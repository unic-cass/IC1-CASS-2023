magic
tech sky130A
magscale 1 2
timestamp 1676037725
<< via4 >>
rect 2269 33811 2505 34047
rect 2589 33811 2825 34047
rect 2909 33811 3145 34047
rect 3229 33811 3465 34047
rect 3549 33811 3785 34047
rect 3869 33811 4105 34047
rect 4189 33811 4425 34047
rect 4509 33811 4745 34047
rect 4829 33811 5065 34047
rect 5149 33811 5385 34047
rect 5469 33811 5705 34047
rect 5789 33811 6025 34047
rect 6109 33811 6345 34047
rect 6429 33811 6665 34047
rect 6749 33811 6985 34047
rect 7069 33811 7305 34047
rect 7389 33811 7625 34047
rect 7709 33811 7945 34047
rect 8029 33811 8265 34047
rect 8349 33811 8585 34047
rect 8669 33811 8905 34047
rect 8989 33811 9225 34047
rect 9309 33811 9545 34047
rect 9629 33811 9865 34047
rect 9949 33811 10185 34047
rect 10269 33811 10505 34047
rect 10589 33811 10825 34047
rect 10909 33811 11145 34047
rect 11229 33811 11465 34047
rect 11549 33811 11785 34047
rect 11869 33811 12105 34047
rect 12189 33811 12425 34047
rect 12509 33811 12745 34047
rect 1947 33503 2183 33739
rect 12871 33449 13107 33685
rect 1627 33183 1863 33419
rect 13191 33129 13427 33365
rect 1307 32863 1543 33099
rect 13511 32809 13747 33045
rect 984 32540 1220 32776
rect 984 32220 1220 32456
rect 13780 32446 14016 32682
rect 984 31900 1220 32136
rect 13780 32126 14016 32362
rect 984 31580 1220 31816
rect 13780 31806 14016 32042
rect 984 31260 1220 31496
rect 13780 31486 14016 31722
rect 984 30940 1220 31176
rect 13780 31166 14016 31402
rect 984 30620 1220 30856
rect 13780 30846 14016 31082
rect 984 30300 1220 30536
rect 13780 30526 14016 30762
rect 984 29980 1220 30216
rect 13780 30206 14016 30442
rect 984 29660 1220 29896
rect 13780 29886 14016 30122
rect 984 29340 1220 29576
rect 13780 29566 14016 29802
rect 984 29020 1220 29256
rect 13780 29246 14016 29482
rect 984 28700 1220 28936
rect 13780 28926 14016 29162
rect 984 28380 1220 28616
rect 13780 28606 14016 28842
rect 984 28060 1220 28296
rect 13780 28286 14016 28522
rect 984 27740 1220 27976
rect 13780 27966 14016 28202
rect 984 27420 1220 27656
rect 13780 27646 14016 27882
rect 984 27100 1220 27336
rect 13780 27326 14016 27562
rect 984 26780 1220 27016
rect 13780 27006 14016 27242
rect 984 26460 1220 26696
rect 13780 26686 14016 26922
rect 984 26140 1220 26376
rect 13780 26366 14016 26602
rect 984 25820 1220 26056
rect 13780 26046 14016 26282
rect 984 25500 1220 25736
rect 13780 25726 14016 25962
rect 984 25180 1220 25416
rect 13780 25406 14016 25642
rect 984 24860 1220 25096
rect 13780 25086 14016 25322
rect 984 24540 1220 24776
rect 13780 24766 14016 25002
rect 984 24220 1220 24456
rect 13780 24446 14016 24682
rect 984 23900 1220 24136
rect 13780 24126 14016 24362
rect 984 23580 1220 23816
rect 13780 23806 14016 24042
rect 984 23260 1220 23496
rect 13780 23486 14016 23722
rect 984 22940 1220 23176
rect 13780 23166 14016 23402
rect 984 22620 1220 22856
rect 13780 22846 14016 23082
rect 984 22300 1220 22536
rect 13780 22526 14016 22762
rect 984 21980 1220 22216
rect 13780 22206 14016 22442
rect 984 21660 1220 21896
rect 13780 21886 14016 22122
rect 984 21340 1220 21576
rect 13780 21566 14016 21802
rect 984 21020 1220 21256
rect 13780 21246 14016 21482
rect 984 20700 1220 20936
rect 13780 20926 14016 21162
rect 984 20380 1220 20616
rect 13780 20606 14016 20842
rect 13780 20286 14016 20522
rect 1253 20017 1489 20253
rect 13457 19963 13693 20199
rect 1573 19697 1809 19933
rect 13137 19643 13373 19879
rect 1893 19377 2129 19613
rect 12817 19323 13053 19559
rect 2255 19015 2491 19251
rect 2575 19015 2811 19251
rect 2895 19015 3131 19251
rect 3215 19015 3451 19251
rect 3535 19015 3771 19251
rect 3855 19015 4091 19251
rect 4175 19015 4411 19251
rect 4495 19015 4731 19251
rect 4815 19015 5051 19251
rect 5135 19015 5371 19251
rect 5455 19015 5691 19251
rect 5775 19015 6011 19251
rect 6095 19015 6331 19251
rect 6415 19015 6651 19251
rect 6735 19015 6971 19251
rect 7055 19015 7291 19251
rect 7375 19015 7611 19251
rect 7695 19015 7931 19251
rect 8015 19015 8251 19251
rect 8335 19015 8571 19251
rect 8655 19015 8891 19251
rect 8975 19015 9211 19251
rect 9295 19015 9531 19251
rect 9615 19015 9851 19251
rect 9935 19015 10171 19251
rect 10255 19015 10491 19251
rect 10575 19015 10811 19251
rect 10895 19015 11131 19251
rect 11215 19015 11451 19251
rect 11535 19015 11771 19251
rect 11855 19015 12091 19251
rect 12175 19015 12411 19251
rect 12495 19015 12731 19251
use sky130_fd_pr__padplhp__example_559591418080  sky130_fd_pr__padplhp__example_559591418080_0
timestamp 1676037725
transform 1 0 1500 0 1 19531
box -540 -540 12540 14540
<< properties >>
string GDS_END 16518
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 16446
<< end >>
