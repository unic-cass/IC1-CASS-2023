magic
tech sky130B
magscale 1 2
timestamp 1676037725
<< metal1 >>
tri 16238 -6692 16244 -6686 se
tri 17056 -6692 17090 -6658 sw
tri 17392 -6692 17426 -6658 se
tri 17472 -6718 17506 -6684 nw
tri 16159 -6772 16193 -6738 nw
rect 21087 -7345 21112 -7317
tri 19541 -7746 19566 -7721 se
rect 19566 -7746 20102 -7721
tri 20102 -7746 20127 -7721 sw
rect 16678 -7749 20715 -7746
rect 16678 -7774 19594 -7749
tri 19594 -7774 19619 -7749 nw
tri 20049 -7774 20074 -7749 ne
rect 20074 -7774 20715 -7749
rect 16678 -7799 16730 -7774
tri 16730 -7808 16764 -7774 nw
tri 19621 -7802 19646 -7777 se
rect 19646 -7802 19993 -7777
tri 19993 -7802 20018 -7777 sw
rect 16791 -7805 20600 -7802
rect 16791 -7830 19674 -7805
tri 19674 -7830 19699 -7805 nw
tri 19940 -7830 19965 -7805 ne
rect 19965 -7830 20600 -7805
tri 16830 -7864 16864 -7830 nw
tri 19694 -7858 19719 -7833 se
tri 16883 -7864 16889 -7858 se
rect 16889 -7864 19827 -7858
tri 16858 -7889 16883 -7864 se
rect 16883 -7886 19827 -7864
rect 16883 -7889 16886 -7886
tri 16505 -8035 16539 -8001 sw
tri 16824 -8035 16858 -8001 se
rect 16858 -8035 16886 -7889
tri 16886 -7912 16912 -7886 nw
tri 17104 -7916 17106 -7914 se
rect 17106 -7916 17574 -7914
rect 16500 -8063 16886 -8035
rect 16500 -8092 16505 -8063
tri 16500 -8097 16505 -8092 ne
tri 16505 -8097 16539 -8063 nw
rect 16922 -8111 17574 -7916
rect 19038 -8681 19039 -8675
tri 19039 -8681 19045 -8675 sw
tri 20148 -9598 20208 -9538 se
rect 20208 -9598 20290 -9538
rect 20036 -9728 20290 -9598
rect 18053 -9806 18125 -9790
tri 18125 -9806 18141 -9790 sw
tri 16159 -9957 16290 -9826 sw
rect 18053 -9836 18141 -9806
tri 18116 -9861 18141 -9836 ne
tri 18141 -9861 18196 -9806 sw
tri 18141 -9916 18196 -9861 ne
tri 18196 -9916 18251 -9861 sw
tri 18827 -9916 18853 -9890 se
rect 18853 -9916 18899 -9888
tri 18899 -9916 18933 -9882 sw
rect 19909 -9916 19955 -9888
tri 18196 -9944 18224 -9916 ne
rect 18224 -9944 19955 -9916
rect 16159 -10159 16389 -9957
tri 18155 -10028 18226 -9957 sw
rect 18155 -10159 18343 -10028
tri 18343 -10159 18344 -10158 nw
tri 16159 -10269 16269 -10159 nw
rect 16668 -10233 18067 -10187
tri 16674 -10262 16703 -10233 nw
tri 16902 -10267 16936 -10233 ne
rect 16936 -10281 18067 -10233
tri 19123 -10267 19189 -10201 se
rect 19189 -10247 19891 -10201
tri 19189 -10267 19209 -10247 nw
rect 16547 -10427 16593 -10397
tri 16547 -10472 16592 -10427 ne
rect 16592 -10444 16593 -10427
tri 16593 -10444 16618 -10419 sw
rect 16592 -10457 16678 -10444
tri 16678 -10457 16691 -10444 sw
rect 16592 -10472 16691 -10457
tri 16662 -10501 16691 -10472 ne
tri 16691 -10501 16735 -10457 sw
rect 16936 -10462 17137 -10281
tri 17137 -10328 17184 -10281 nw
tri 19081 -10309 19123 -10267 se
rect 19123 -10309 19147 -10267
tri 19147 -10309 19189 -10267 nw
rect 17460 -10354 18234 -10309
rect 17460 -10355 18195 -10354
tri 18195 -10355 18196 -10354 nw
tri 18233 -10355 18234 -10354 ne
rect 18364 -10354 19102 -10309
tri 19102 -10354 19147 -10309 nw
tri 18364 -10355 18365 -10354 nw
tri 17323 -10401 17369 -10355 ne
tri 17137 -10462 17171 -10428 sw
tri 16691 -10545 16735 -10501 ne
tri 16735 -10545 16779 -10501 sw
rect 16936 -10508 17210 -10462
tri 17343 -10545 17369 -10519 se
rect 17369 -10545 17397 -10355
tri 17397 -10401 17443 -10355 nw
tri 16735 -10573 16763 -10545 ne
rect 16763 -10553 17397 -10545
rect 16763 -10573 17377 -10553
tri 17377 -10573 17397 -10553 nw
rect 17535 -10542 17581 -10506
tri 17535 -10588 17581 -10542 ne
tri 17581 -10572 17631 -10522 sw
rect 17581 -10588 17907 -10572
tri 17581 -10618 17611 -10588 ne
rect 17611 -10618 17907 -10588
tri 18926 -10743 19098 -10571 se
rect 19098 -10701 19615 -10571
rect 19098 -10738 19236 -10701
rect 19098 -10743 19159 -10738
tri 19236 -10767 19302 -10701 nw
tri 17385 -10825 17419 -10791 ne
tri 17465 -10825 17499 -10791 nw
tri 17925 -10825 17959 -10791 ne
tri 18005 -10825 18039 -10791 nw
tri 18121 -10797 18127 -10791 ne
tri 18257 -10845 18291 -10811 se
tri 18365 -10924 18399 -10890 se
tri 18445 -10934 18479 -10900 sw
tri 18389 -10980 18399 -10970 ne
tri 17797 -11010 17800 -11007 se
rect 17800 -11010 17801 -11007
rect 17927 -11010 17928 -11007
tri 17928 -11010 17931 -11007 sw
tri 17797 -11059 17800 -11056 ne
tri 17928 -11059 17931 -11056 nw
tri 18679 -11104 18713 -11070 se
tri 18759 -11090 18793 -11056 nw
tri 18772 -11178 18806 -11144 se
tri 18834 -11164 18868 -11130 nw
tri 20093 -11335 20096 -11332 se
tri 20315 -11335 20318 -11332 sw
tri 20639 -11335 20673 -11301 se
rect 17333 -11434 17354 -11376
tri 17354 -11434 17412 -11376 nw
tri 20093 -11384 20096 -11381 ne
tri 20315 -11384 20318 -11381 nw
rect 17059 -11489 17060 -11465
tri 17060 -11489 17084 -11465 sw
tri 19593 -11489 19618 -11464 se
tri 19746 -11489 19771 -11464 sw
tri 19989 -11490 19993 -11486 se
rect 19993 -11490 19994 -11486
tri 19972 -11538 19993 -11517 ne
tri 16635 -11564 16636 -11563 sw
rect 16863 -11581 19775 -11553
rect 16863 -11605 16990 -11581
tri 16990 -11605 17014 -11581 nw
rect 16633 -11615 16635 -11610
tri 16635 -11615 16640 -11610 nw
tri 18081 -11624 18095 -11610 se
rect 18095 -11624 18105 -11610
tri 19741 -11615 19775 -11581 ne
tri 18084 -11662 18095 -11651 ne
rect 18095 -11662 18101 -11651
rect 18222 -11662 18223 -11648
tri 18223 -11662 18237 -11648 nw
tri 19518 -11662 19532 -11648 ne
rect 19532 -11662 19534 -11648
tri 17525 -11699 17535 -11689 sw
tri 18345 -11699 18368 -11676 se
tri 17525 -11761 17559 -11727 nw
tri 18366 -11728 18368 -11726 ne
rect 18368 -11728 18369 -11726
tri 18478 -11762 18484 -11756 se
tri 17700 -11814 17724 -11790 nw
tri 18466 -11808 18484 -11790 ne
tri 17795 -11868 17819 -11844 se
rect 20992 -11873 21032 -7425
rect 21072 -11800 21112 -7345
rect 21160 -11744 21188 -7816
rect 21236 -11687 21264 -7832
tri 22737 -8633 22755 -8615 se
rect 22881 -8639 22883 -8615
tri 22883 -8639 22907 -8615 sw
rect 22881 -8640 25670 -8639
rect 22883 -8664 25670 -8640
tri 25670 -8664 25695 -8639 sw
tri 26724 -8664 26773 -8615 se
rect 26773 -8664 26774 -8615
rect 22883 -8667 26906 -8664
tri 25585 -8696 25614 -8667 ne
rect 25614 -8696 26906 -8667
tri 23054 -9427 23088 -9393 sw
tri 22876 -9465 22910 -9431 se
tri 23356 -10151 23361 -10146 sw
tri 23356 -10198 23361 -10193 nw
tri 21264 -11687 21298 -11653 sw
rect 23829 -11687 24082 -11663
rect 21236 -11691 24082 -11687
tri 21188 -11744 21222 -11710 sw
rect 21236 -11715 23857 -11691
tri 21112 -11800 21146 -11766 sw
rect 21160 -11772 23909 -11744
tri 24112 -11800 24138 -11774 se
rect 24138 -11800 24142 -11774
rect 21072 -11824 24142 -11800
tri 21072 -11839 21087 -11824 ne
rect 21087 -11826 24142 -11824
rect 21087 -11839 24129 -11826
tri 24129 -11839 24142 -11826 nw
rect 24471 -11831 24667 -11629
tri 22784 -11873 22790 -11867 se
tri 22918 -11873 22924 -11867 sw
tri 24139 -11873 24158 -11854 se
rect 24158 -11873 24159 -11854
rect 20992 -11906 24189 -11873
rect 20992 -11913 22867 -11906
tri 22784 -11919 22790 -11913 ne
tri 22918 -11919 22931 -11906 nw
tri 19639 -11947 19663 -11923 se
tri 19791 -11947 19815 -11923 sw
tri 16459 -12009 16493 -11975 nw
tri 17047 -12016 17060 -12003 sw
rect 17047 -12046 24298 -12016
tri 17047 -12055 17056 -12046 nw
tri 24438 -12076 24471 -12043 se
rect 24471 -12076 24601 -11831
tri 24601 -11897 24667 -11831 nw
tri 17457 -12126 17481 -12102 nw
tri 16789 -12170 16823 -12136 sw
tri 16696 -12226 16725 -12197 sw
rect 24360 -12206 24601 -12076
rect 16691 -12255 16696 -12251
tri 16696 -12255 16700 -12251 nw
tri 16576 -12293 16610 -12259 sw
tri 23721 -12323 23727 -12317 ne
tri 23855 -12323 23861 -12317 nw
tri 17700 -12404 17722 -12382 nw
tri 24281 -12392 24288 -12385 se
tri 17950 -12549 18089 -12410 se
rect 18089 -12549 18800 -12410
tri 24592 -12507 24693 -12406 se
tri 24760 -12485 24820 -12425 sw
rect 18009 -12569 18800 -12549
tri 18009 -12717 18157 -12569 nw
tri 24617 -12666 24647 -12636 ne
tri 17408 -12785 17414 -12779 se
tri 17524 -13055 17562 -13017 ne
tri 17614 -13051 17648 -13017 nw
tri 16942 -13089 16960 -13071 se
tri 17012 -13090 17041 -13061 sw
tri 16775 -13156 16809 -13122 ne
tri 17865 -13173 17899 -13139 se
tri 16634 -13286 16668 -13252 sw
tri 16223 -13372 16267 -13328 se
tri 16338 -13405 16397 -13346 sw
tri 16634 -13366 16668 -13332 nw
tri 16482 -13405 16502 -13385 se
tri 16548 -13405 16568 -13385 sw
<< metal2 >>
tri 16970 -6686 17004 -6652 se
rect 18357 -7479 18385 -7412
tri 18385 -7479 18392 -7472 sw
rect 18357 -7496 18392 -7479
tri 18357 -7531 18392 -7496 ne
tri 18392 -7531 18444 -7479 sw
tri 18392 -7583 18444 -7531 ne
tri 18444 -7583 18496 -7531 sw
tri 18444 -7607 18468 -7583 ne
tri 16658 -8734 16697 -8695 se
rect 16697 -8725 16725 -7816
tri 17523 -7972 17577 -7918 se
rect 17577 -7934 17615 -7718
tri 17615 -7808 17705 -7718 nw
tri 17577 -7972 17615 -7934 nw
tri 17498 -7997 17523 -7972 se
rect 17523 -7997 17536 -7972
rect 17498 -8681 17536 -7997
tri 17536 -8013 17577 -7972 nw
rect 16697 -8734 16716 -8725
tri 16716 -8734 16725 -8725 nw
rect 16648 -8786 16664 -8734
tri 16664 -8786 16716 -8734 nw
rect 16648 -9557 16673 -9513
tri 16673 -9557 16717 -9513 sw
rect 16648 -9565 16717 -9557
tri 16659 -9595 16689 -9565 ne
tri 16668 -9751 16689 -9730 se
rect 16689 -9751 16717 -9565
tri 16775 -9582 16809 -9548 nw
rect 16668 -9764 16717 -9751
tri 16539 -11002 16573 -10968 ne
tri 16539 -11154 16573 -11120 se
tri 16610 -11154 16640 -11124 sw
tri 16478 -11164 16484 -11158 nw
tri 16539 -11240 16573 -11206 ne
tri 16610 -11236 16640 -11206 nw
tri 16539 -11563 16573 -11529 se
tri 16613 -11563 16635 -11541 sw
tri 16473 -11654 16484 -11643 sw
tri 16340 -11711 16352 -11699 se
tri 16276 -11768 16300 -11744 sw
tri 16407 -12099 16431 -12075 ne
rect 16431 -13054 16459 -12075
tri 16644 -12127 16668 -12103 se
tri 16644 -12279 16668 -12255 ne
tri 16625 -13046 16668 -13003 se
rect 16668 -13018 16696 -9764
tri 16696 -9785 16717 -9764 nw
rect 17779 -10890 17831 -8811
rect 18127 -10554 18330 -8141
rect 18127 -10792 18258 -10554
tri 18258 -10626 18330 -10554 nw
tri 17779 -10942 17831 -10890 ne
tri 17831 -10895 17858 -10868 sw
rect 17831 -10942 17961 -10895
tri 17831 -10947 17836 -10942 ne
rect 17836 -10947 17961 -10942
tri 17939 -10969 17961 -10947 ne
tri 17961 -10948 18014 -10895 sw
rect 17961 -10969 18014 -10948
tri 17961 -10990 17982 -10969 ne
tri 17473 -11841 17497 -11817 ne
tri 17340 -12074 17374 -12040 se
tri 17426 -12074 17457 -12043 sw
tri 17464 -12779 17497 -12746 se
rect 17497 -12779 17525 -11817
tri 17600 -11848 17634 -11814 nw
tri 17841 -11844 17875 -11810 se
tri 17903 -11844 17937 -11810 sw
tri 17600 -12352 17634 -12318 sw
tri 17600 -12438 17634 -12404 nw
tri 17525 -12779 17542 -12762 sw
tri 17936 -12887 17982 -12841 se
rect 17982 -12855 18014 -10969
rect 18468 -11688 18496 -7583
tri 18903 -7755 18940 -7718 ne
tri 18910 -8675 18940 -8645 se
rect 18940 -8675 18984 -7718
tri 18984 -7765 19031 -7718 nw
tri 18984 -8675 19039 -8620 sw
rect 19454 -9144 20370 -9116
rect 19454 -9393 19506 -9144
tri 19506 -9178 19540 -9144 nw
tri 20290 -9178 20324 -9144 ne
rect 19355 -10032 19407 -9887
tri 19355 -10082 19405 -10032 ne
rect 19405 -10060 19407 -10032
tri 19407 -10060 19457 -10010 sw
tri 19371 -11409 19405 -11375 se
rect 19405 -11409 19457 -10060
tri 19457 -11409 19471 -11395 sw
tri 19684 -11464 19718 -11430 se
tri 19684 -11550 19718 -11516 ne
tri 19532 -11610 19535 -11607 se
tri 19572 -11610 19606 -11576 sw
tri 18512 -11756 18546 -11722 se
tri 18574 -11756 18608 -11722 sw
tri 18014 -11836 18048 -11802 sw
tri 18014 -11922 18048 -11888 nw
tri 19663 -11923 19718 -11868 se
rect 19718 -11975 19746 -9216
tri 19746 -9302 19780 -9268 nw
tri 19982 -9456 20048 -9390 se
rect 20048 -9410 20094 -9312
tri 20048 -9456 20094 -9410 nw
tri 19916 -9522 19982 -9456 se
tri 19982 -9522 20048 -9456 nw
tri 19890 -9548 19916 -9522 se
rect 19916 -9548 19936 -9522
rect 19890 -10195 19936 -9548
tri 19936 -9568 19982 -9522 nw
rect 20324 -9665 20370 -9144
rect 22787 -9694 22839 -8667
rect 22776 -9746 22839 -9694
rect 22776 -10046 22821 -9746
tri 22821 -10046 22839 -10028 sw
rect 22776 -10098 22839 -10046
tri 22776 -10109 22787 -10098 ne
tri 19936 -10195 19970 -10161 sw
rect 22787 -10518 22839 -10098
tri 23269 -10232 23303 -10198 ne
rect 23303 -10200 23356 -10198
rect 22787 -10570 23094 -10518
tri 19993 -11486 20023 -11456 se
tri 20051 -11486 20085 -11452 sw
rect 23042 -11760 23094 -10570
rect 23303 -11599 23355 -10200
tri 23355 -10201 23356 -10200 nw
rect 23042 -11797 23809 -11760
tri 23042 -11812 23057 -11797 ne
rect 23057 -11812 23809 -11797
tri 19746 -11923 19791 -11878 sw
tri 20912 -11926 20946 -11892 ne
tri 22822 -12002 22918 -11906 ne
tri 22918 -11941 22931 -11928 sw
rect 22918 -12002 22931 -11941
tri 22918 -12015 22931 -12002 ne
tri 22931 -12015 23005 -11941 sw
tri 22931 -12089 23005 -12015 ne
tri 23005 -12089 23079 -12015 sw
tri 23005 -12163 23079 -12089 ne
tri 23079 -12163 23153 -12089 sw
tri 23079 -12237 23153 -12163 ne
tri 23153 -12237 23227 -12163 sw
tri 23153 -12259 23175 -12237 ne
rect 23175 -12346 23227 -12237
rect 23757 -12271 23809 -11812
rect 23980 -12143 24008 -11772
rect 24082 -12071 24110 -11715
rect 24267 -11826 25445 -11774
tri 25445 -11826 25497 -11774 sw
tri 25439 -11884 25497 -11826 ne
tri 25497 -11865 25536 -11826 sw
rect 25497 -11884 25603 -11865
tri 25497 -11917 25530 -11884 ne
rect 25530 -11917 25603 -11884
tri 26070 -11890 26126 -11834 se
rect 26126 -11862 27734 -11834
tri 27734 -11862 27762 -11834 sw
rect 26126 -11890 26128 -11862
tri 26128 -11890 26156 -11862 nw
rect 24152 -11949 24581 -11934
tri 24581 -11949 24596 -11934 sw
tri 26012 -11948 26070 -11890 se
tri 26070 -11948 26128 -11890 nw
tri 27710 -11914 27762 -11862 ne
tri 27762 -11914 27814 -11862 sw
rect 24152 -11962 24596 -11949
rect 24426 -12001 24529 -11996
tri 24529 -12001 24534 -11996 sw
tri 24557 -12001 24596 -11962 ne
tri 24596 -12001 24648 -11949 sw
tri 25982 -11978 26012 -11948 se
rect 24426 -12035 24534 -12001
tri 24534 -12035 24568 -12001 sw
rect 24426 -12048 24568 -12035
tri 24082 -12099 24110 -12071 ne
tri 24110 -12089 24146 -12053 sw
tri 24531 -12085 24568 -12048 ne
tri 24568 -12053 24586 -12035 sw
tri 24596 -12053 24648 -12001 ne
tri 24648 -12053 24700 -12001 sw
tri 25429 -12006 25457 -11978 se
rect 25457 -12006 26012 -11978
tri 26012 -12006 26070 -11948 nw
tri 27762 -11966 27814 -11914 ne
tri 27814 -11966 27866 -11914 sw
tri 26118 -11973 26125 -11966 se
rect 26125 -11973 27119 -11966
tri 27119 -11973 27126 -11966 sw
rect 24568 -12085 24586 -12053
tri 24586 -12085 24618 -12053 sw
rect 24110 -12099 24488 -12089
tri 24110 -12117 24128 -12099 ne
rect 24128 -12117 24488 -12099
tri 24008 -12143 24021 -12130 sw
tri 24462 -12143 24488 -12117 ne
tri 24488 -12135 24534 -12089 sw
tri 24568 -12135 24618 -12085 ne
tri 24618 -12105 24638 -12085 sw
tri 24648 -12105 24700 -12053 ne
tri 24700 -12105 24752 -12053 sw
tri 25380 -12055 25429 -12006 se
rect 25429 -12055 25431 -12006
tri 25431 -12055 25480 -12006 nw
tri 26073 -12018 26118 -11973 se
rect 26118 -11994 27126 -11973
rect 26118 -12018 26125 -11994
tri 26065 -12026 26073 -12018 se
rect 26073 -12026 26125 -12018
tri 26125 -12026 26157 -11994 nw
tri 27098 -12022 27126 -11994 ne
tri 27126 -12022 27175 -11973 sw
tri 27814 -12018 27866 -11966 ne
tri 27866 -12018 27918 -11966 sw
rect 24618 -12135 24638 -12105
tri 24638 -12135 24668 -12105 sw
rect 24488 -12143 24534 -12135
rect 23980 -12153 24021 -12143
tri 23980 -12192 24019 -12153 ne
rect 24019 -12192 24021 -12153
tri 24021 -12192 24070 -12143 sw
tri 24488 -12187 24532 -12143 ne
rect 24532 -12187 24534 -12143
tri 24534 -12187 24586 -12135 sw
tri 24618 -12185 24668 -12135 ne
tri 24668 -12156 24689 -12135 sw
tri 24700 -12156 24751 -12105 ne
rect 24751 -12129 24810 -12105
tri 25329 -12106 25380 -12055 se
tri 25380 -12106 25431 -12055 nw
tri 26005 -12086 26065 -12026 se
tri 26065 -12086 26125 -12026 nw
tri 27126 -12043 27147 -12022 ne
tri 25306 -12129 25329 -12106 se
rect 24668 -12185 24689 -12156
tri 24689 -12185 24718 -12156 sw
rect 24751 -12157 25329 -12129
tri 25329 -12157 25380 -12106 nw
tri 25945 -12146 26005 -12086 se
tri 26005 -12146 26065 -12086 nw
tri 26469 -12103 26521 -12051 se
rect 26521 -12103 26678 -12051
tri 25922 -12169 25945 -12146 se
rect 25945 -12169 25948 -12146
tri 25460 -12185 25466 -12179 se
rect 25466 -12185 25717 -12179
tri 24019 -12220 24047 -12192 ne
rect 24047 -12220 24446 -12192
tri 24424 -12242 24446 -12220 ne
tri 24446 -12241 24495 -12192 sw
tri 24532 -12241 24586 -12187 ne
tri 24586 -12241 24640 -12187 sw
tri 24668 -12213 24696 -12185 ne
rect 24696 -12207 25717 -12185
rect 25791 -12203 25948 -12169
tri 25948 -12203 26005 -12146 nw
tri 26419 -12153 26469 -12103 se
tri 26469 -12153 26519 -12103 nw
tri 26369 -12203 26419 -12153 se
tri 26419 -12203 26469 -12153 nw
rect 27147 -12179 27175 -12022
tri 27866 -12070 27918 -12018 ne
tri 27918 -12070 27970 -12018 sw
tri 27918 -12106 27954 -12070 ne
rect 27954 -12082 27970 -12070
tri 27970 -12082 27982 -12070 sw
rect 27954 -12148 27982 -12082
rect 24696 -12213 25484 -12207
tri 25484 -12213 25490 -12207 nw
rect 25791 -12221 25930 -12203
tri 25930 -12221 25948 -12203 nw
rect 24446 -12242 24495 -12241
tri 24446 -12281 24485 -12242 ne
rect 24485 -12281 24495 -12242
tri 24495 -12281 24535 -12241 sw
tri 24586 -12269 24614 -12241 ne
rect 24614 -12269 24796 -12241
tri 25017 -12281 25049 -12249 se
rect 25049 -12281 25064 -12249
tri 26319 -12253 26369 -12203 se
tri 26369 -12253 26419 -12203 nw
tri 24485 -12331 24535 -12281 ne
tri 24535 -12331 24585 -12281 sw
tri 25003 -12295 25017 -12281 se
rect 25017 -12293 25064 -12281
rect 25017 -12295 25041 -12293
tri 24967 -12331 25003 -12295 se
rect 25003 -12303 25041 -12295
tri 25041 -12303 25051 -12293 nw
tri 26269 -12303 26319 -12253 se
tri 26319 -12303 26369 -12253 nw
rect 25003 -12331 25013 -12303
tri 25013 -12331 25041 -12303 nw
tri 24535 -12359 24563 -12331 ne
rect 24563 -12359 24985 -12331
tri 24985 -12359 25013 -12331 nw
tri 26219 -12353 26269 -12303 se
tri 26269 -12353 26319 -12303 nw
rect 24416 -12392 24523 -12385
tri 24523 -12392 24530 -12385 sw
tri 26180 -12392 26219 -12353 se
rect 24416 -12403 26219 -12392
tri 26219 -12403 26269 -12353 nw
rect 24416 -12420 26202 -12403
tri 26202 -12420 26219 -12403 nw
tri 24416 -12437 24433 -12420 nw
tri 17982 -12887 18014 -12855 nw
tri 16668 -13046 16696 -13018 nw
tri 17899 -12924 17936 -12887 se
rect 17936 -12924 17951 -12887
tri 17951 -12918 17982 -12887 nw
tri 16582 -13089 16625 -13046 se
tri 16625 -13089 16668 -13046 nw
tri 16539 -13132 16582 -13089 se
tri 16582 -13132 16625 -13089 nw
tri 16529 -13142 16539 -13132 se
rect 16539 -13142 16572 -13132
tri 16572 -13142 16582 -13132 nw
rect 16502 -13194 16520 -13142
tri 16520 -13194 16572 -13142 nw
tri 16719 -13162 16747 -13134 se
rect 17899 -13207 17951 -12924
<< metal3 >>
tri 17694 -8710 17844 -8560 se
rect 17844 -8677 18073 -7911
rect 17844 -8710 17962 -8677
rect 17694 -9077 17962 -8710
tri 17962 -8788 18073 -8677 nw
tri 17962 -9077 18038 -9001 sw
rect 17694 -9079 18038 -9077
tri 17694 -9179 17794 -9079 ne
rect 17794 -9253 18038 -9079
tri 17448 -13661 17794 -13315 se
rect 17794 -13417 18038 -13207
tri 17794 -13661 18038 -13417 nw
tri 26847 -13573 27137 -13283 se
rect 27137 -13403 27423 -11215
rect 27137 -13573 27299 -13403
tri 27299 -13527 27423 -13403 nw
tri 17220 -13889 17448 -13661 se
rect 17448 -13889 17464 -13661
rect 17220 -15244 17464 -13889
tri 17464 -13991 17794 -13661 nw
use sky130_fd_io__amx_inv1  sky130_fd_io__amx_inv1_0
timestamp 1676037725
transform -1 0 16742 0 -1 -10035
box 118 36 220 682
use sky130_fd_io__amx_inv1  sky130_fd_io__amx_inv1_1
timestamp 1676037725
transform 1 0 20176 0 -1 -9456
box 118 36 220 682
use sky130_fd_io__amx_inv1  sky130_fd_io__amx_inv1_2
timestamp 1676037725
transform 1 0 16560 0 -1 -10035
box 118 36 220 682
use sky130_fd_io__gpiov2_amux_drvr_ls  sky130_fd_io__gpiov2_amux_drvr_ls_0
timestamp 1676037725
transform 1 0 16331 0 1 -9217
box 38 39 1829 964
use sky130_fd_io__gpiov2_amux_drvr_ls  sky130_fd_io__gpiov2_amux_drvr_ls_1
timestamp 1676037725
transform 1 0 24609 0 1 -12705
box 38 39 1829 964
use sky130_fd_io__gpiov2_amux_drvr_ls  sky130_fd_io__gpiov2_amux_drvr_ls_2
timestamp 1676037725
transform -1 0 20092 0 1 -9217
box 38 39 1829 964
use sky130_fd_io__gpiov2_amux_drvr_ls  sky130_fd_io__gpiov2_amux_drvr_ls_3
timestamp 1676037725
transform 1 0 16331 0 -1 -9083
box 38 39 1829 964
use sky130_fd_io__gpiov2_amux_drvr_ls  sky130_fd_io__gpiov2_amux_drvr_ls_4
timestamp 1676037725
transform 1 0 16185 0 1 -13625
box 38 39 1829 964
use sky130_fd_io__gpiov2_amux_drvr_ls  sky130_fd_io__gpiov2_amux_drvr_ls_5
timestamp 1676037725
transform -1 0 28283 0 1 -12705
box 38 39 1829 964
use sky130_fd_io__gpiov2_amux_drvr_lshv2hv2  sky130_fd_io__gpiov2_amux_drvr_lshv2hv2_0
timestamp 1676037725
transform -1 0 21030 0 1 -8115
box 371 123 4711 3822
use sky130_fd_io__gpiov2_amux_drvr_lshv2hv  sky130_fd_io__gpiov2_amux_drvr_lshv2hv_0
timestamp 1676037725
transform 1 0 17744 0 1 -8115
box -1425 123 1533 3328
use sky130_fd_io__gpiov2_amx_inv4  sky130_fd_io__gpiov2_amx_inv4_0
timestamp 1676037725
transform 1 0 19218 0 -1 -9588
box 118 36 416 351
use sky130_fd_io__gpiov2_amx_inv4  sky130_fd_io__gpiov2_amx_inv4_1
timestamp 1676037725
transform -1 0 19400 0 -1 -9588
box 118 36 416 351
use sky130_fd_io__gpiov2_amx_inv4  sky130_fd_io__gpiov2_amx_inv4_2
timestamp 1676037725
transform -1 0 23372 0 1 -12646
box 118 36 416 351
use sky130_fd_io__gpiov2_amx_inv4  sky130_fd_io__gpiov2_amx_inv4_3
timestamp 1676037725
transform -1 0 20104 0 -1 -9588
box 118 36 416 351
use sky130_fd_io__gpiov2_amx_inv4  sky130_fd_io__gpiov2_amx_inv4_4
timestamp 1676037725
transform 1 0 22486 0 1 -12646
box 118 36 416 351
use sky130_fd_io__gpiov2_amx_inv4  sky130_fd_io__gpiov2_amx_inv4_5
timestamp 1676037725
transform -1 0 19048 0 -1 -9588
box 118 36 416 351
use sky130_fd_io__gpiov2_amx_pucsd_inv  sky130_fd_io__gpiov2_amx_pucsd_inv_0
timestamp 1676037725
transform 1 0 23189 0 1 -12655
box 119 45 1297 360
use sky130_fd_io__hvsbt_inv_x1  sky130_fd_io__hvsbt_inv_x1_0
timestamp 1676037725
transform 1 0 23264 0 1 -11502
box 107 226 240 873
use sky130_fd_io__hvsbt_inv_x1  sky130_fd_io__hvsbt_inv_x1_1
timestamp 1676037725
transform -1 0 22742 0 1 -11502
box 107 226 240 873
use sky130_fd_io__hvsbt_inv_x2  sky130_fd_io__hvsbt_inv_x2_0
timestamp 1676037725
transform 1 0 22912 0 1 -11502
box 107 226 460 873
use sky130_fd_io__hvsbt_inv_x2  sky130_fd_io__hvsbt_inv_x2_1
timestamp 1676037725
transform 1 0 22560 0 1 -11502
box 107 226 460 873
use sky130_fd_pr__nfet_01v8__example_55959141808576  sky130_fd_pr__nfet_01v8__example_55959141808576_0
timestamp 1676037725
transform 1 0 19943 0 1 -9509
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808577  sky130_fd_pr__nfet_01v8__example_55959141808577_0
timestamp 1676037725
transform 0 -1 17492 1 0 -10306
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808578  sky130_fd_pr__nfet_01v8__example_55959141808578_0
timestamp 1676037725
transform 0 -1 17492 1 0 -10462
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808579  sky130_fd_pr__nfet_01v8__example_55959141808579_0
timestamp 1676037725
transform 1 0 19676 0 1 -9509
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808579  sky130_fd_pr__nfet_01v8__example_55959141808579_1
timestamp 1676037725
transform -1 0 18914 0 -1 -9309
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808579  sky130_fd_pr__nfet_01v8__example_55959141808579_2
timestamp 1676037725
transform -1 0 19620 0 1 -9509
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808579  sky130_fd_pr__nfet_01v8__example_55959141808579_3
timestamp 1676037725
transform 1 0 18970 0 -1 -9309
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808572  sky130_fd_pr__pfet_01v8__example_55959141808572_0
timestamp 1676037725
transform 1 0 18313 0 1 -10530
box -1 0 401 1
use sky130_fd_pr__pfet_01v8__example_55959141808573  sky130_fd_pr__pfet_01v8__example_55959141808573_0
timestamp 1676037725
transform 1 0 17857 0 1 -10530
box -1 0 401 1
<< properties >>
string GDS_END 43750940
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 43608254
<< end >>
