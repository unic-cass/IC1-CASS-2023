magic
tech sky130A
magscale 1 2
timestamp 1676037725
<< metal2 >>
rect -6231 23152 -1085 23500
rect -6231 22896 -6130 23152
rect -5874 22896 -5606 23152
rect -5350 22896 -5052 23152
rect -4796 22896 -4498 23152
rect -4242 22896 -3944 23152
rect -3688 22896 -3390 23152
rect -3134 22896 -2836 23152
rect -2580 22896 -2312 23152
rect -2056 22896 -1085 23152
rect -6231 22628 -1085 22896
rect -6231 22372 -6130 22628
rect -5874 22372 -5606 22628
rect -5350 22372 -5052 22628
rect -4796 22372 -4498 22628
rect -4242 22372 -3944 22628
rect -3688 22372 -3390 22628
rect -3134 22372 -2836 22628
rect -2580 22372 -2312 22628
rect -2056 22372 -1085 22628
rect -6231 22104 -1085 22372
rect -6231 21848 -6130 22104
rect -5874 21848 -5606 22104
rect -5350 21848 -5052 22104
rect -4796 21848 -4498 22104
rect -4242 21848 -3944 22104
rect -3688 21848 -3390 22104
rect -3134 21848 -2836 22104
rect -2580 21848 -2312 22104
rect -2056 21848 -1085 22104
rect -6231 21500 -1085 21848
tri -1915 21330 -1745 21500 ne
rect -1745 21330 -1085 21500
tri -1085 21330 1085 23500 sw
tri -1745 18500 1085 21330 ne
tri 1085 20500 1915 21330 sw
rect 1085 20151 6008 20500
rect 1085 19895 1833 20151
rect 2089 19895 2357 20151
rect 2613 19895 2911 20151
rect 3167 19895 3465 20151
rect 3721 19895 4019 20151
rect 4275 19895 4573 20151
rect 4829 19895 5127 20151
rect 5383 19895 5651 20151
rect 5907 19895 6008 20151
rect 1085 19627 6008 19895
rect 1085 19371 1833 19627
rect 2089 19371 2357 19627
rect 2613 19371 2911 19627
rect 3167 19371 3465 19627
rect 3721 19371 4019 19627
rect 4275 19371 4573 19627
rect 4829 19371 5127 19627
rect 5383 19371 5651 19627
rect 5907 19371 6008 19627
rect 1085 19103 6008 19371
rect 1085 18847 1833 19103
rect 2089 18847 2357 19103
rect 2613 18847 2911 19103
rect 3167 18847 3465 19103
rect 3721 18847 4019 19103
rect 4275 18847 4573 19103
rect 4829 18847 5127 19103
rect 5383 18847 5651 19103
rect 5907 18847 6008 19103
rect 1085 18500 6008 18847
rect -6231 17153 -1085 17500
rect -6231 16897 -6131 17153
rect -5875 16897 -5607 17153
rect -5351 16897 -5053 17153
rect -4797 16897 -4499 17153
rect -4243 16897 -3945 17153
rect -3689 16897 -3391 17153
rect -3135 16897 -2837 17153
rect -2581 16897 -2313 17153
rect -2057 16897 -1085 17153
rect -6231 16629 -1085 16897
rect -6231 16373 -6131 16629
rect -5875 16373 -5607 16629
rect -5351 16373 -5053 16629
rect -4797 16373 -4499 16629
rect -4243 16373 -3945 16629
rect -3689 16373 -3391 16629
rect -3135 16373 -2837 16629
rect -2581 16373 -2313 16629
rect -2057 16373 -1085 16629
rect -6231 16105 -1085 16373
rect -6231 15849 -6131 16105
rect -5875 15849 -5607 16105
rect -5351 15849 -5053 16105
rect -4797 15849 -4499 16105
rect -4243 15849 -3945 16105
rect -3689 15849 -3391 16105
rect -3135 15849 -2837 16105
rect -2581 15849 -2313 16105
rect -2057 15849 -1085 16105
rect -6231 15500 -1085 15849
tri -1915 15330 -1745 15500 ne
rect -1745 15330 -1085 15500
tri -1085 15330 1085 17500 sw
tri -1745 12500 1085 15330 ne
tri 1085 14500 1915 15330 sw
rect 1085 14153 6008 14500
rect 1085 13897 1833 14153
rect 2089 13897 2357 14153
rect 2613 13897 2911 14153
rect 3167 13897 3465 14153
rect 3721 13897 4019 14153
rect 4275 13897 4573 14153
rect 4829 13897 5127 14153
rect 5383 13897 5651 14153
rect 5907 13897 6008 14153
rect 1085 13629 6008 13897
rect 1085 13373 1833 13629
rect 2089 13373 2357 13629
rect 2613 13373 2911 13629
rect 3167 13373 3465 13629
rect 3721 13373 4019 13629
rect 4275 13373 4573 13629
rect 4829 13373 5127 13629
rect 5383 13373 5651 13629
rect 5907 13373 6008 13629
rect 1085 13105 6008 13373
rect 1085 12849 1833 13105
rect 2089 12849 2357 13105
rect 2613 12849 2911 13105
rect 3167 12849 3465 13105
rect 3721 12849 4019 13105
rect 4275 12849 4573 13105
rect 4829 12849 5127 13105
rect 5383 12849 5651 13105
rect 5907 12849 6008 13105
rect 1085 12500 6008 12849
rect 9908 652 27500 1000
rect 9908 396 10052 652
rect 10308 396 10576 652
rect 10832 396 11130 652
rect 11386 396 27500 652
rect 9908 128 27500 396
rect 9908 -128 10052 128
rect 10308 -128 10576 128
rect 10832 -128 11130 128
rect 11386 -128 27500 128
rect 9908 -396 27500 -128
rect 9908 -652 10052 -396
rect 10308 -652 10576 -396
rect 10832 -652 11130 -396
rect 11386 -652 27500 -396
rect 9908 -1000 27500 -652
tri -1745 -18330 1085 -15500 se
rect 1085 -15849 6008 -15500
rect 1085 -16105 1832 -15849
rect 2088 -16105 2356 -15849
rect 2612 -16105 2910 -15849
rect 3166 -16105 3464 -15849
rect 3720 -16105 4018 -15849
rect 4274 -16105 4572 -15849
rect 4828 -16105 5126 -15849
rect 5382 -16105 5650 -15849
rect 5906 -16105 6008 -15849
rect 1085 -16373 6008 -16105
rect 1085 -16629 1832 -16373
rect 2088 -16629 2356 -16373
rect 2612 -16629 2910 -16373
rect 3166 -16629 3464 -16373
rect 3720 -16629 4018 -16373
rect 4274 -16629 4572 -16373
rect 4828 -16629 5126 -16373
rect 5382 -16629 5650 -16373
rect 5906 -16629 6008 -16373
rect 1085 -16897 6008 -16629
rect 1085 -17153 1832 -16897
rect 2088 -17153 2356 -16897
rect 2612 -17153 2910 -16897
rect 3166 -17153 3464 -16897
rect 3720 -17153 4018 -16897
rect 4274 -17153 4572 -16897
rect 4828 -17153 5126 -16897
rect 5382 -17153 5650 -16897
rect 5906 -17153 6008 -16897
rect 1085 -17500 6008 -17153
tri 1085 -18330 1915 -17500 nw
tri -1915 -18500 -1745 -18330 se
rect -1745 -18500 -1085 -18330
rect -6231 -18848 -1085 -18500
rect -6231 -19104 -6130 -18848
rect -5874 -19104 -5606 -18848
rect -5350 -19104 -5052 -18848
rect -4796 -19104 -4498 -18848
rect -4242 -19104 -3944 -18848
rect -3688 -19104 -3390 -18848
rect -3134 -19104 -2836 -18848
rect -2580 -19104 -2312 -18848
rect -2056 -19104 -1085 -18848
rect -6231 -19372 -1085 -19104
rect -6231 -19628 -6130 -19372
rect -5874 -19628 -5606 -19372
rect -5350 -19628 -5052 -19372
rect -4796 -19628 -4498 -19372
rect -4242 -19628 -3944 -19372
rect -3688 -19628 -3390 -19372
rect -3134 -19628 -2836 -19372
rect -2580 -19628 -2312 -19372
rect -2056 -19628 -1085 -19372
rect -6231 -19896 -1085 -19628
rect -6231 -20152 -6130 -19896
rect -5874 -20152 -5606 -19896
rect -5350 -20152 -5052 -19896
rect -4796 -20152 -4498 -19896
rect -4242 -20152 -3944 -19896
rect -3688 -20152 -3390 -19896
rect -3134 -20152 -2836 -19896
rect -2580 -20152 -2312 -19896
rect -2056 -20152 -1085 -19896
rect -6231 -20500 -1085 -20152
tri -1085 -20500 1085 -18330 nw
tri -1745 -24330 1085 -21500 se
rect 1085 -21848 6008 -21500
rect 1085 -22104 1833 -21848
rect 2089 -22104 2357 -21848
rect 2613 -22104 2911 -21848
rect 3167 -22104 3465 -21848
rect 3721 -22104 4019 -21848
rect 4275 -22104 4573 -21848
rect 4829 -22104 5127 -21848
rect 5383 -22104 5651 -21848
rect 5907 -22104 6008 -21848
rect 1085 -22372 6008 -22104
rect 1085 -22628 1833 -22372
rect 2089 -22628 2357 -22372
rect 2613 -22628 2911 -22372
rect 3167 -22628 3465 -22372
rect 3721 -22628 4019 -22372
rect 4275 -22628 4573 -22372
rect 4829 -22628 5127 -22372
rect 5383 -22628 5651 -22372
rect 5907 -22628 6008 -22372
rect 1085 -22896 6008 -22628
rect 1085 -23152 1833 -22896
rect 2089 -23152 2357 -22896
rect 2613 -23152 2911 -22896
rect 3167 -23152 3465 -22896
rect 3721 -23152 4019 -22896
rect 4275 -23152 4573 -22896
rect 4829 -23152 5127 -22896
rect 5383 -23152 5651 -22896
rect 5907 -23152 6008 -22896
rect 1085 -23500 6008 -23152
tri 1085 -24330 1915 -23500 nw
tri -1915 -24500 -1745 -24330 se
rect -1745 -24500 -1085 -24330
rect -6231 -24848 -1085 -24500
rect -6231 -25104 -6130 -24848
rect -5874 -25104 -5606 -24848
rect -5350 -25104 -5052 -24848
rect -4796 -25104 -4498 -24848
rect -4242 -25104 -3944 -24848
rect -3688 -25104 -3390 -24848
rect -3134 -25104 -2836 -24848
rect -2580 -25104 -2312 -24848
rect -2056 -25104 -1085 -24848
rect -6231 -25372 -1085 -25104
rect -6231 -25628 -6130 -25372
rect -5874 -25628 -5606 -25372
rect -5350 -25628 -5052 -25372
rect -4796 -25628 -4498 -25372
rect -4242 -25628 -3944 -25372
rect -3688 -25628 -3390 -25372
rect -3134 -25628 -2836 -25372
rect -2580 -25628 -2312 -25372
rect -2056 -25628 -1085 -25372
rect -6231 -25896 -1085 -25628
rect -6231 -26152 -6130 -25896
rect -5874 -26152 -5606 -25896
rect -5350 -26152 -5052 -25896
rect -4796 -26152 -4498 -25896
rect -4242 -26152 -3944 -25896
rect -3688 -26152 -3390 -25896
rect -3134 -26152 -2836 -25896
rect -2580 -26152 -2312 -25896
rect -2056 -26152 -1085 -25896
rect -6231 -26500 -1085 -26152
tri -1085 -26500 1085 -24330 nw
<< via2 >>
rect -6130 22896 -5874 23152
rect -5606 22896 -5350 23152
rect -5052 22896 -4796 23152
rect -4498 22896 -4242 23152
rect -3944 22896 -3688 23152
rect -3390 22896 -3134 23152
rect -2836 22896 -2580 23152
rect -2312 22896 -2056 23152
rect -6130 22372 -5874 22628
rect -5606 22372 -5350 22628
rect -5052 22372 -4796 22628
rect -4498 22372 -4242 22628
rect -3944 22372 -3688 22628
rect -3390 22372 -3134 22628
rect -2836 22372 -2580 22628
rect -2312 22372 -2056 22628
rect -6130 21848 -5874 22104
rect -5606 21848 -5350 22104
rect -5052 21848 -4796 22104
rect -4498 21848 -4242 22104
rect -3944 21848 -3688 22104
rect -3390 21848 -3134 22104
rect -2836 21848 -2580 22104
rect -2312 21848 -2056 22104
rect 1833 19895 2089 20151
rect 2357 19895 2613 20151
rect 2911 19895 3167 20151
rect 3465 19895 3721 20151
rect 4019 19895 4275 20151
rect 4573 19895 4829 20151
rect 5127 19895 5383 20151
rect 5651 19895 5907 20151
rect 1833 19371 2089 19627
rect 2357 19371 2613 19627
rect 2911 19371 3167 19627
rect 3465 19371 3721 19627
rect 4019 19371 4275 19627
rect 4573 19371 4829 19627
rect 5127 19371 5383 19627
rect 5651 19371 5907 19627
rect 1833 18847 2089 19103
rect 2357 18847 2613 19103
rect 2911 18847 3167 19103
rect 3465 18847 3721 19103
rect 4019 18847 4275 19103
rect 4573 18847 4829 19103
rect 5127 18847 5383 19103
rect 5651 18847 5907 19103
rect -6131 16897 -5875 17153
rect -5607 16897 -5351 17153
rect -5053 16897 -4797 17153
rect -4499 16897 -4243 17153
rect -3945 16897 -3689 17153
rect -3391 16897 -3135 17153
rect -2837 16897 -2581 17153
rect -2313 16897 -2057 17153
rect -6131 16373 -5875 16629
rect -5607 16373 -5351 16629
rect -5053 16373 -4797 16629
rect -4499 16373 -4243 16629
rect -3945 16373 -3689 16629
rect -3391 16373 -3135 16629
rect -2837 16373 -2581 16629
rect -2313 16373 -2057 16629
rect -6131 15849 -5875 16105
rect -5607 15849 -5351 16105
rect -5053 15849 -4797 16105
rect -4499 15849 -4243 16105
rect -3945 15849 -3689 16105
rect -3391 15849 -3135 16105
rect -2837 15849 -2581 16105
rect -2313 15849 -2057 16105
rect 1833 13897 2089 14153
rect 2357 13897 2613 14153
rect 2911 13897 3167 14153
rect 3465 13897 3721 14153
rect 4019 13897 4275 14153
rect 4573 13897 4829 14153
rect 5127 13897 5383 14153
rect 5651 13897 5907 14153
rect 1833 13373 2089 13629
rect 2357 13373 2613 13629
rect 2911 13373 3167 13629
rect 3465 13373 3721 13629
rect 4019 13373 4275 13629
rect 4573 13373 4829 13629
rect 5127 13373 5383 13629
rect 5651 13373 5907 13629
rect 1833 12849 2089 13105
rect 2357 12849 2613 13105
rect 2911 12849 3167 13105
rect 3465 12849 3721 13105
rect 4019 12849 4275 13105
rect 4573 12849 4829 13105
rect 5127 12849 5383 13105
rect 5651 12849 5907 13105
rect 10052 396 10308 652
rect 10576 396 10832 652
rect 11130 396 11386 652
rect 10052 -128 10308 128
rect 10576 -128 10832 128
rect 11130 -128 11386 128
rect 10052 -652 10308 -396
rect 10576 -652 10832 -396
rect 11130 -652 11386 -396
rect 1832 -16105 2088 -15849
rect 2356 -16105 2612 -15849
rect 2910 -16105 3166 -15849
rect 3464 -16105 3720 -15849
rect 4018 -16105 4274 -15849
rect 4572 -16105 4828 -15849
rect 5126 -16105 5382 -15849
rect 5650 -16105 5906 -15849
rect 1832 -16629 2088 -16373
rect 2356 -16629 2612 -16373
rect 2910 -16629 3166 -16373
rect 3464 -16629 3720 -16373
rect 4018 -16629 4274 -16373
rect 4572 -16629 4828 -16373
rect 5126 -16629 5382 -16373
rect 5650 -16629 5906 -16373
rect 1832 -17153 2088 -16897
rect 2356 -17153 2612 -16897
rect 2910 -17153 3166 -16897
rect 3464 -17153 3720 -16897
rect 4018 -17153 4274 -16897
rect 4572 -17153 4828 -16897
rect 5126 -17153 5382 -16897
rect 5650 -17153 5906 -16897
rect -6130 -19104 -5874 -18848
rect -5606 -19104 -5350 -18848
rect -5052 -19104 -4796 -18848
rect -4498 -19104 -4242 -18848
rect -3944 -19104 -3688 -18848
rect -3390 -19104 -3134 -18848
rect -2836 -19104 -2580 -18848
rect -2312 -19104 -2056 -18848
rect -6130 -19628 -5874 -19372
rect -5606 -19628 -5350 -19372
rect -5052 -19628 -4796 -19372
rect -4498 -19628 -4242 -19372
rect -3944 -19628 -3688 -19372
rect -3390 -19628 -3134 -19372
rect -2836 -19628 -2580 -19372
rect -2312 -19628 -2056 -19372
rect -6130 -20152 -5874 -19896
rect -5606 -20152 -5350 -19896
rect -5052 -20152 -4796 -19896
rect -4498 -20152 -4242 -19896
rect -3944 -20152 -3688 -19896
rect -3390 -20152 -3134 -19896
rect -2836 -20152 -2580 -19896
rect -2312 -20152 -2056 -19896
rect 1833 -22104 2089 -21848
rect 2357 -22104 2613 -21848
rect 2911 -22104 3167 -21848
rect 3465 -22104 3721 -21848
rect 4019 -22104 4275 -21848
rect 4573 -22104 4829 -21848
rect 5127 -22104 5383 -21848
rect 5651 -22104 5907 -21848
rect 1833 -22628 2089 -22372
rect 2357 -22628 2613 -22372
rect 2911 -22628 3167 -22372
rect 3465 -22628 3721 -22372
rect 4019 -22628 4275 -22372
rect 4573 -22628 4829 -22372
rect 5127 -22628 5383 -22372
rect 5651 -22628 5907 -22372
rect 1833 -23152 2089 -22896
rect 2357 -23152 2613 -22896
rect 2911 -23152 3167 -22896
rect 3465 -23152 3721 -22896
rect 4019 -23152 4275 -22896
rect 4573 -23152 4829 -22896
rect 5127 -23152 5383 -22896
rect 5651 -23152 5907 -22896
rect -6130 -25104 -5874 -24848
rect -5606 -25104 -5350 -24848
rect -5052 -25104 -4796 -24848
rect -4498 -25104 -4242 -24848
rect -3944 -25104 -3688 -24848
rect -3390 -25104 -3134 -24848
rect -2836 -25104 -2580 -24848
rect -2312 -25104 -2056 -24848
rect -6130 -25628 -5874 -25372
rect -5606 -25628 -5350 -25372
rect -5052 -25628 -4796 -25372
rect -4498 -25628 -4242 -25372
rect -3944 -25628 -3688 -25372
rect -3390 -25628 -3134 -25372
rect -2836 -25628 -2580 -25372
rect -2312 -25628 -2056 -25372
rect -6130 -26152 -5874 -25896
rect -5606 -26152 -5350 -25896
rect -5052 -26152 -4796 -25896
rect -4498 -26152 -4242 -25896
rect -3944 -26152 -3688 -25896
rect -3390 -26152 -3134 -25896
rect -2836 -26152 -2580 -25896
rect -2312 -26152 -2056 -25896
<< metal3 >>
tri -13806 23672 -10978 26500 se
rect -10978 25118 10978 26500
tri 10978 25118 12360 26500 sw
rect -10978 24500 12360 25118
tri -10978 23672 -10150 24500 nw
tri -16634 20844 -13806 23672 se
rect -13806 22258 -12392 23672
tri -12392 22258 -10978 23672 nw
tri 10150 23500 11150 24500 ne
rect 11150 23500 12360 24500
tri -10978 22258 -9736 23500 se
rect -9736 23253 -2202 23500
tri -2202 23253 -1955 23500 sw
rect -9736 23152 -1955 23253
rect -9736 22896 -6130 23152
rect -5874 22896 -5606 23152
rect -5350 22896 -5052 23152
rect -4796 22896 -4498 23152
rect -4242 22896 -3944 23152
rect -3688 22896 -3390 23152
rect -3134 22896 -2836 23152
rect -2580 22896 -2312 23152
rect -2056 22896 -1955 23152
rect -9736 22628 -1955 22896
rect -9736 22372 -6130 22628
rect -5874 22372 -5606 22628
rect -5350 22372 -5052 22628
rect -4796 22372 -4498 22628
rect -4242 22372 -3944 22628
rect -3688 22372 -3390 22628
rect -3134 22372 -2836 22628
rect -2580 22372 -2312 22628
rect -2056 22372 -1955 22628
rect -9736 22258 -1955 22372
tri -13806 20844 -12392 22258 nw
tri -12392 20844 -10978 22258 se
rect -10978 22104 -1955 22258
rect -10978 21848 -6130 22104
rect -5874 21848 -5606 22104
rect -5350 21848 -5052 22104
rect -4796 21848 -4498 22104
rect -4242 21848 -3944 22104
rect -3688 21848 -3390 22104
rect -3134 21848 -2836 22104
rect -2580 21848 -2312 22104
rect -2056 21848 -1955 22104
rect -10978 21747 -1955 21848
rect -10978 21500 -2202 21747
tri -2202 21500 -1955 21747 nw
rect -10978 20844 -9736 21500
tri -19462 18016 -16634 20844 se
rect -16634 19430 -15220 20844
tri -15220 19430 -13806 20844 nw
tri -12564 20672 -12392 20844 se
rect -12392 20672 -9736 20844
tri -9736 20672 -8908 21500 nw
tri -13806 19430 -12564 20672 se
rect -12564 19430 -11151 20672
tri -16634 18016 -15220 19430 nw
tri -15220 18016 -13806 19430 se
rect -13806 19257 -11151 19430
tri -11151 19257 -9736 20672 nw
tri -1745 20670 1085 23500 se
rect 1085 22290 9736 23500
tri 9736 22290 10946 23500 sw
tri 11150 22290 12360 23500 ne
tri 12360 22290 15188 25118 sw
rect 1085 21500 10946 22290
tri 1085 20670 1915 21500 nw
tri 8908 20672 9736 21500 ne
rect 9736 21048 10946 21500
tri 10946 21048 12188 22290 sw
rect 9736 20876 12188 21048
tri 12188 20876 12360 21048 sw
tri 12360 20876 13774 22290 ne
rect 13774 20876 15188 22290
rect 9736 20672 12360 20876
tri -1915 20500 -1745 20670 se
rect -1745 20500 -1085 20670
tri -9736 19257 -8493 20500 se
rect -8493 19257 -1085 20500
rect -13806 18016 -12564 19257
tri -22290 15188 -19462 18016 se
rect -19462 16602 -18048 18016
tri -18048 16602 -16634 18016 nw
tri -15392 17844 -15220 18016 se
rect -15220 17844 -12564 18016
tri -12564 17844 -11151 19257 nw
tri -11149 17844 -9736 19257 se
rect -9736 18500 -1085 19257
tri -1085 18500 1085 20670 nw
tri 1732 20253 1979 20500 se
rect 1979 20253 8493 20500
rect 1732 20151 8493 20253
rect 1732 19895 1833 20151
rect 2089 19895 2357 20151
rect 2613 19895 2911 20151
rect 3167 19895 3465 20151
rect 3721 19895 4019 20151
rect 4275 19895 4573 20151
rect 4829 19895 5127 20151
rect 5383 19895 5651 20151
rect 5907 19895 8493 20151
rect 1732 19805 8493 19895
tri 8493 19805 9188 20500 sw
rect 1732 19627 9188 19805
rect 1732 19371 1833 19627
rect 2089 19371 2357 19627
rect 2613 19371 2911 19627
rect 3167 19371 3465 19627
rect 3721 19371 4019 19627
rect 4275 19371 4573 19627
rect 4829 19371 5127 19627
rect 5383 19371 5651 19627
rect 5907 19371 9188 19627
rect 1732 19257 9188 19371
tri 9188 19257 9736 19805 sw
tri 9736 19257 11151 20672 ne
rect 11151 19462 12360 20672
tri 12360 19462 13774 20876 sw
tri 13774 19462 15188 20876 ne
tri 15188 19462 18016 22290 sw
rect 11151 19257 13774 19462
rect 1732 19103 9736 19257
rect 1732 18847 1833 19103
rect 2089 18847 2357 19103
rect 2613 18847 2911 19103
rect 3167 18847 3465 19103
rect 3721 18847 4019 19103
rect 4275 18847 4573 19103
rect 4829 18847 5127 19103
rect 5383 18847 5651 19103
rect 5907 18847 9736 19103
rect 1732 18747 9736 18847
tri 1732 18500 1979 18747 ne
rect 1979 18500 9736 18747
rect -9736 17844 -8493 18500
tri -16634 16602 -15392 17844 se
rect -15392 16602 -13979 17844
tri -19462 15188 -18048 16602 nw
tri -18048 15188 -16634 16602 se
rect -16634 16429 -13979 16602
tri -13979 16429 -12564 17844 nw
tri -11321 17672 -11149 17844 se
rect -11149 17672 -8493 17844
tri -8493 17672 -7665 18500 nw
tri -12564 16429 -11321 17672 se
rect -11321 16429 -9907 17672
rect -16634 15188 -15392 16429
tri -25118 12360 -22290 15188 se
rect -22290 13774 -20876 15188
tri -20876 13774 -19462 15188 nw
tri -18220 15016 -18048 15188 se
rect -18048 15016 -15392 15188
tri -15392 15016 -13979 16429 nw
tri -13977 15016 -12564 16429 se
rect -12564 16258 -9907 16429
tri -9907 16258 -8493 17672 nw
tri 7665 17500 8665 18500 ne
rect 8665 18220 9736 18500
tri 9736 18220 10773 19257 sw
tri 11151 18220 12188 19257 ne
rect 12188 18220 13774 19257
tri 13774 18220 15016 19462 sw
rect 8665 17500 10773 18220
tri -8493 16258 -7251 17500 se
rect -7251 17253 -2202 17500
tri -2202 17253 -1955 17500 sw
rect -7251 17153 -1955 17253
rect -7251 16897 -6131 17153
rect -5875 16897 -5607 17153
rect -5351 16897 -5053 17153
rect -4797 16897 -4499 17153
rect -4243 16897 -3945 17153
rect -3689 16897 -3391 17153
rect -3135 16897 -2837 17153
rect -2581 16897 -2313 17153
rect -2057 16897 -1955 17153
rect -7251 16629 -1955 16897
rect -7251 16373 -6131 16629
rect -5875 16373 -5607 16629
rect -5351 16373 -5053 16629
rect -4797 16373 -4499 16629
rect -4243 16373 -3945 16629
rect -3689 16373 -3391 16629
rect -3135 16373 -2837 16629
rect -2581 16373 -2313 16629
rect -2057 16373 -1955 16629
rect -7251 16258 -1955 16373
rect -12564 15016 -11321 16258
tri -19462 13774 -18220 15016 se
rect -18220 13774 -16807 15016
tri -22290 12360 -20876 13774 nw
tri -20876 12360 -19462 13774 se
rect -19462 13601 -16807 13774
tri -16807 13601 -15392 15016 nw
tri -14149 14844 -13977 15016 se
rect -13977 14844 -11321 15016
tri -11321 14844 -9907 16258 nw
tri -9907 14844 -8493 16258 se
rect -8493 16105 -1955 16258
rect -8493 15849 -6131 16105
rect -5875 15849 -5607 16105
rect -5351 15849 -5053 16105
rect -4797 15849 -4499 16105
rect -4243 15849 -3945 16105
rect -3689 15849 -3391 16105
rect -3135 15849 -2837 16105
rect -2581 15849 -2313 16105
rect -2057 15849 -1955 16105
rect -8493 15747 -1955 15849
rect -8493 15500 -2202 15747
tri -2202 15500 -1955 15747 nw
rect -8493 14844 -7251 15500
tri -15392 13601 -14149 14844 se
rect -14149 13601 -12735 14844
rect -19462 12360 -18220 13601
tri -26500 10978 -25118 12360 se
rect -25118 10978 -23672 12360
tri -23672 10978 -22290 12360 nw
tri -22258 10978 -20876 12360 se
rect -20876 12188 -18220 12360
tri -18220 12188 -16807 13601 nw
tri -16805 12188 -15392 13601 se
rect -15392 13430 -12735 13601
tri -12735 13430 -11321 14844 nw
tri -10079 14672 -9907 14844 se
rect -9907 14672 -7251 14844
tri -7251 14672 -6423 15500 nw
tri -11321 13430 -10079 14672 se
rect -10079 13430 -8666 14672
rect -15392 12188 -14149 13430
rect -20876 10978 -19635 12188
rect -26500 -10978 -24500 10978
tri -24500 10150 -23672 10978 nw
tri -23500 9736 -22258 10978 se
rect -22258 10773 -19635 10978
tri -19635 10773 -18220 12188 nw
tri -16977 12016 -16805 12188 se
rect -16805 12016 -14149 12188
tri -14149 12016 -12735 13430 nw
tri -12735 12016 -11321 13430 se
rect -11321 13257 -8666 13430
tri -8666 13257 -7251 14672 nw
tri -1745 14670 1085 17500 se
rect 1085 16977 7251 17500
tri 7251 16977 7774 17500 sw
tri 8665 16977 9188 17500 ne
rect 9188 16977 10773 17500
tri 10773 16977 12016 18220 sw
rect 1085 15735 7774 16977
tri 7774 15735 9016 16977 sw
rect 1085 15563 9016 15735
tri 9016 15563 9188 15735 sw
tri 9188 15563 10602 16977 ne
rect 10602 16805 12016 16977
tri 12016 16805 12188 16977 sw
tri 12188 16805 13603 18220 ne
rect 13603 18048 15016 18220
tri 15016 18048 15188 18220 sw
tri 15188 18048 16602 19462 ne
rect 16602 18048 18016 19462
rect 13603 16805 15188 18048
rect 10602 15563 12188 16805
rect 1085 15500 9188 15563
tri 1085 14670 1915 15500 nw
tri -1915 14500 -1745 14670 se
rect -1745 14500 -1085 14670
tri -7251 13257 -6008 14500 se
rect -6008 13257 -1085 14500
rect -11321 12016 -10079 13257
tri -18220 10773 -16977 12016 se
rect -16977 10773 -15563 12016
rect -22258 9736 -20672 10773
tri -20672 9736 -19635 10773 nw
tri -19257 9736 -18220 10773 se
rect -18220 10602 -15563 10773
tri -15563 10602 -14149 12016 nw
tri -12907 11844 -12735 12016 se
rect -12735 11844 -10079 12016
tri -10079 11844 -8666 13257 nw
tri -8664 11844 -7251 13257 se
rect -7251 12500 -1085 13257
tri -1085 12500 1085 14670 nw
tri 1732 14253 1979 14500 se
rect 1979 14492 6008 14500
tri 6008 14492 6016 14500 sw
tri 6423 14492 7431 15500 ne
rect 7431 14492 9188 15500
rect 1979 14253 6016 14492
rect 1732 14153 6016 14253
rect 1732 13897 1833 14153
rect 2089 13897 2357 14153
rect 2613 13897 2911 14153
rect 3167 13897 3465 14153
rect 3721 13897 4019 14153
rect 4275 13897 4573 14153
rect 4829 13897 5127 14153
rect 5383 13897 5651 14153
rect 5907 13897 6016 14153
rect 1732 13629 6016 13897
rect 1732 13373 1833 13629
rect 2089 13373 2357 13629
rect 2613 13373 2911 13629
rect 3167 13373 3465 13629
rect 3721 13373 4019 13629
rect 4275 13373 4573 13629
rect 4829 13373 5127 13629
rect 5383 13373 5651 13629
rect 5907 13373 6016 13629
rect 1732 13257 6016 13373
tri 6016 13257 7251 14492 sw
tri 7431 13257 8666 14492 ne
rect 8666 14149 9188 14492
tri 9188 14149 10602 15563 sw
tri 10602 14149 12016 15563 ne
rect 12016 15392 12188 15563
tri 12188 15392 13601 16805 sw
tri 13603 15392 15016 16805 ne
rect 15016 16634 15188 16805
tri 15188 16634 16602 18048 sw
tri 16602 16634 18016 18048 ne
tri 18016 16634 20844 19462 sw
rect 15016 15392 16602 16634
tri 16602 15392 17844 16634 sw
rect 12016 14149 13601 15392
tri 13601 14149 14844 15392 sw
rect 8666 13257 10602 14149
rect 1732 13105 7251 13257
rect 1732 12849 1833 13105
rect 2089 12849 2357 13105
rect 2613 12849 2911 13105
rect 3167 12849 3465 13105
rect 3721 12849 4019 13105
rect 4275 12849 4573 13105
rect 4829 12849 5127 13105
rect 5383 12849 5651 13105
rect 5907 12907 7251 13105
tri 7251 12907 7601 13257 sw
tri 8666 12907 9016 13257 ne
rect 9016 12907 10602 13257
tri 10602 12907 11844 14149 sw
rect 5907 12849 7601 12907
rect 1732 12747 7601 12849
tri 1732 12500 1979 12747 ne
rect 1979 12500 7601 12747
rect -7251 11844 -6008 12500
tri -14149 10602 -12907 11844 se
rect -12907 10602 -11494 11844
rect -18220 9736 -16977 10602
rect -23500 -9736 -21500 9736
tri -21500 8908 -20672 9736 nw
tri -20500 8493 -19257 9736 se
rect -19257 9188 -16977 9736
tri -16977 9188 -15563 10602 nw
tri -15563 9188 -14149 10602 se
rect -14149 10429 -11494 10602
tri -11494 10429 -10079 11844 nw
tri -8836 11672 -8664 11844 se
rect -8664 11672 -6008 11844
tri -6008 11672 -5180 12500 nw
tri -10079 10429 -8836 11672 se
rect -14149 9188 -12907 10429
rect -19257 8493 -17672 9188
tri -17672 8493 -16977 9188 nw
tri -16258 8493 -15563 9188 se
rect -15563 9016 -12907 9188
tri -12907 9016 -11494 10429 nw
tri -11492 9016 -10079 10429 se
rect -10079 9016 -8836 10429
rect -15563 8493 -14322 9016
rect -20500 -8493 -18500 8493
tri -18500 7665 -17672 8493 nw
tri -17500 7251 -16258 8493 se
rect -16258 7601 -14322 8493
tri -14322 7601 -12907 9016 nw
tri -11664 8844 -11492 9016 se
rect -11492 8844 -8836 9016
tri -8836 8844 -6008 11672 nw
tri 5180 11664 6016 12500 ne
rect 6016 11664 7601 12500
tri 7601 11664 8844 12907 sw
tri -12907 7601 -11664 8844 se
rect -16258 7251 -14672 7601
tri -14672 7251 -14322 7601 nw
tri -13257 7251 -12907 7601 se
rect -12907 7251 -11664 7601
rect -17500 -7251 -15500 7251
tri -15500 6423 -14672 7251 nw
tri -14500 6008 -13257 7251 se
rect -13257 6016 -11664 7251
tri -11664 6016 -8836 8844 nw
tri 6016 8836 8844 11664 ne
tri 8844 11492 9016 11664 sw
tri 9016 11492 10431 12907 ne
rect 10431 12735 11844 12907
tri 11844 12735 12016 12907 sw
tri 12016 12735 13430 14149 ne
rect 13430 13977 14844 14149
tri 14844 13977 15016 14149 sw
tri 15016 13977 16431 15392 ne
rect 16431 15220 17844 15392
tri 17844 15220 18016 15392 sw
tri 18016 15220 19430 16634 ne
rect 19430 15220 20844 16634
rect 16431 13977 18016 15220
rect 13430 12735 15016 13977
rect 10431 11492 12016 12735
rect 8844 10079 9016 11492
tri 9016 10079 10429 11492 sw
tri 10431 10079 11844 11492 ne
rect 11844 11321 12016 11492
tri 12016 11321 13430 12735 sw
tri 13430 11321 14844 12735 ne
rect 14844 12564 15016 12735
tri 15016 12564 16429 13977 sw
tri 16431 12564 17844 13977 ne
rect 17844 13806 18016 13977
tri 18016 13806 19430 15220 sw
tri 19430 13806 20844 15220 ne
tri 20844 13806 23672 16634 sw
rect 17844 12564 19430 13806
tri 19430 12564 20672 13806 sw
rect 14844 11321 16429 12564
tri 16429 11321 17672 12564 sw
rect 11844 10079 13430 11321
tri 13430 10079 14672 11321 sw
rect 8844 8836 10429 10079
tri 10429 8836 11672 10079 sw
rect -13257 6008 -12500 6016
rect -14500 1000 -12500 6008
tri -12500 5180 -11664 6016 nw
tri 8844 6008 11672 8836 ne
tri 11672 8664 11844 8836 sw
tri 11844 8664 13259 10079 ne
rect 13259 9907 14672 10079
tri 14672 9907 14844 10079 sw
tri 14844 9907 16258 11321 ne
rect 16258 11149 17672 11321
tri 17672 11149 17844 11321 sw
tri 17844 11149 19259 12564 ne
rect 19259 12392 20672 12564
tri 20672 12392 20844 12564 sw
tri 20844 12392 22258 13806 ne
rect 22258 12392 23672 13806
rect 19259 11149 20844 12392
rect 16258 9907 17844 11149
rect 13259 8664 14844 9907
rect 11672 7251 11844 8664
tri 11844 7251 13257 8664 sw
tri 13259 7251 14672 8664 ne
rect 14672 8493 14844 8664
tri 14844 8493 16258 9907 sw
tri 16258 8493 17672 9907 ne
rect 17672 9736 17844 9907
tri 17844 9736 19257 11149 sw
tri 19259 9736 20672 11149 ne
rect 20672 10978 20844 11149
tri 20844 10978 22258 12392 sw
tri 22258 10978 23672 12392 ne
tri 23672 10978 26500 13806 sw
rect 20672 9736 22258 10978
tri 22258 9736 23500 10978 sw
tri 23672 10150 24500 10978 ne
rect 17672 8493 19257 9736
tri 19257 8493 20500 9736 sw
tri 20672 8908 21500 9736 ne
rect 14672 7251 16258 8493
tri 16258 7251 17500 8493 sw
tri 17672 7665 18500 8493 ne
rect 11672 6008 13257 7251
tri 13257 6008 14500 7251 sw
tri 14672 6423 15500 7251 ne
tri 11672 5180 12500 6008 ne
rect -14500 652 11500 1000
rect -14500 396 10052 652
rect 10308 396 10576 652
rect 10832 396 11130 652
rect 11386 396 11500 652
rect -14500 128 11500 396
rect -14500 -128 10052 128
rect 10308 -128 10576 128
rect 10832 -128 11130 128
rect 11386 -128 11500 128
rect -14500 -396 11500 -128
rect -14500 -652 10052 -396
rect 10308 -652 10576 -396
rect 10832 -652 11130 -396
rect 11386 -652 11500 -396
rect -14500 -1000 11500 -652
rect -14500 -6008 -12500 -1000
tri -12500 -6008 -11672 -5180 sw
tri -15500 -7251 -14672 -6423 sw
tri -14500 -7251 -13257 -6008 ne
rect -13257 -7251 -11672 -6008
tri -18500 -8493 -17672 -7665 sw
tri -17500 -8493 -16258 -7251 ne
rect -16258 -8493 -14672 -7251
tri -21500 -9736 -20672 -8908 sw
tri -20500 -9736 -19257 -8493 ne
rect -19257 -9736 -17672 -8493
tri -24500 -10978 -23672 -10150 sw
tri -23500 -10978 -22258 -9736 ne
rect -22258 -10978 -20672 -9736
tri -26500 -13806 -23672 -10978 ne
tri -23672 -12392 -22258 -10978 sw
tri -22258 -12392 -20844 -10978 ne
rect -20844 -11149 -20672 -10978
tri -20672 -11149 -19259 -9736 sw
tri -19257 -11149 -17844 -9736 ne
rect -17844 -9907 -17672 -9736
tri -17672 -9907 -16258 -8493 sw
tri -16258 -9907 -14844 -8493 ne
rect -14844 -8664 -14672 -8493
tri -14672 -8664 -13259 -7251 sw
tri -13257 -8664 -11844 -7251 ne
rect -11844 -8664 -11672 -7251
rect -14844 -9907 -13259 -8664
rect -17844 -11149 -16258 -9907
rect -20844 -12392 -19259 -11149
rect -23672 -13806 -22258 -12392
tri -22258 -13806 -20844 -12392 sw
tri -20844 -12564 -20672 -12392 ne
rect -20672 -12564 -19259 -12392
tri -19259 -12564 -17844 -11149 sw
tri -17844 -11321 -17672 -11149 ne
rect -17672 -11321 -16258 -11149
tri -16258 -11321 -14844 -9907 sw
tri -14844 -10079 -14672 -9907 ne
rect -14672 -10079 -13259 -9907
tri -13259 -10079 -11844 -8664 sw
tri -11844 -8836 -11672 -8664 ne
tri -11672 -8836 -8844 -6008 sw
tri 11664 -6016 12500 -5180 se
rect 12500 -6008 14500 6008
rect 12500 -6016 13257 -6008
tri -11672 -10079 -10429 -8836 ne
rect -10429 -10079 -8844 -8836
tri -14672 -11321 -13430 -10079 ne
rect -13430 -11321 -11844 -10079
tri -17672 -12564 -16429 -11321 ne
rect -16429 -12564 -14844 -11321
tri -20672 -13806 -19430 -12564 ne
rect -19430 -13806 -17844 -12564
tri -23672 -16634 -20844 -13806 ne
tri -20844 -15220 -19430 -13806 sw
tri -19430 -15220 -18016 -13806 ne
rect -18016 -13977 -17844 -13806
tri -17844 -13977 -16431 -12564 sw
tri -16429 -13977 -15016 -12564 ne
rect -15016 -12735 -14844 -12564
tri -14844 -12735 -13430 -11321 sw
tri -13430 -12735 -12016 -11321 ne
rect -12016 -11492 -11844 -11321
tri -11844 -11492 -10431 -10079 sw
tri -10429 -11492 -9016 -10079 ne
rect -9016 -11492 -8844 -10079
rect -12016 -12735 -10431 -11492
rect -15016 -13977 -13430 -12735
rect -18016 -15220 -16431 -13977
rect -20844 -16634 -19430 -15220
tri -19430 -16634 -18016 -15220 sw
tri -18016 -15392 -17844 -15220 ne
rect -17844 -15392 -16431 -15220
tri -16431 -15392 -15016 -13977 sw
tri -15016 -14149 -14844 -13977 ne
rect -14844 -14149 -13430 -13977
tri -13430 -14149 -12016 -12735 sw
tri -12016 -12907 -11844 -12735 ne
rect -11844 -12907 -10431 -12735
tri -10431 -12907 -9016 -11492 sw
tri -9016 -11664 -8844 -11492 ne
tri -8844 -11664 -6016 -8836 sw
tri 8836 -8844 11664 -6016 se
rect 11664 -7251 13257 -6016
tri 13257 -7251 14500 -6008 nw
tri 14672 -7251 15500 -6423 se
rect 15500 -7251 17500 7251
rect 11664 -7601 12907 -7251
tri 12907 -7601 13257 -7251 nw
tri 11664 -8844 12907 -7601 nw
tri 13430 -8493 14672 -7251 se
rect 14672 -8493 16258 -7251
tri 16258 -8493 17500 -7251 nw
tri 17672 -8493 18500 -7665 se
rect 18500 -8493 20500 8493
tri -8844 -12907 -7601 -11664 ne
rect -7601 -12500 -6016 -11664
tri -6016 -12500 -5180 -11664 sw
tri 6008 -11672 8836 -8844 se
rect 8836 -9016 11492 -8844
tri 11492 -9016 11664 -8844 nw
tri 12907 -9016 13430 -8493 se
rect 13430 -9016 15015 -8493
rect 8836 -10429 10079 -9016
tri 10079 -10429 11492 -9016 nw
tri 11494 -10429 12907 -9016 se
rect 12907 -9736 15015 -9016
tri 15015 -9736 16258 -8493 nw
tri 16429 -9736 17672 -8493 se
rect 17672 -9736 19257 -8493
tri 19257 -9736 20500 -8493 nw
tri 20672 -9736 21500 -8908 se
rect 21500 -9736 23500 9736
rect 24500 5000 26500 10978
rect 24500 3000 27500 5000
rect 12907 -10429 14149 -9736
tri 8836 -11672 10079 -10429 nw
tri 5180 -12500 6008 -11672 se
rect 6008 -11844 8664 -11672
tri 8664 -11844 8836 -11672 nw
tri 10079 -11844 11494 -10429 se
rect 11494 -10602 14149 -10429
tri 14149 -10602 15015 -9736 nw
rect 11494 -11844 12907 -10602
tri 12907 -11844 14149 -10602 nw
tri 15187 -10978 16429 -9736 se
rect 16429 -10978 18015 -9736
tri 18015 -10978 19257 -9736 nw
tri 19430 -10978 20672 -9736 se
rect 20672 -10978 22258 -9736
tri 22258 -10978 23500 -9736 nw
rect 24500 -5000 27500 -3000
tri 23672 -10978 24500 -10150 se
rect 24500 -10978 26500 -5000
rect 6008 -12500 7251 -11844
rect -7601 -12907 7251 -12500
tri -11844 -14149 -10602 -12907 ne
rect -10602 -13257 -9016 -12907
tri -9016 -13257 -8666 -12907 sw
tri -7601 -13257 -7251 -12907 ne
rect -7251 -13257 7251 -12907
tri 7251 -13257 8664 -11844 nw
tri 8666 -13257 10079 -11844 se
rect 10079 -12016 12735 -11844
tri 12735 -12016 12907 -11844 nw
tri 14149 -12016 15187 -10978 se
rect 15187 -12016 16977 -10978
tri 16977 -12016 18015 -10978 nw
rect 10079 -13257 11321 -12016
rect -10602 -14149 -8666 -13257
tri -14844 -15392 -13601 -14149 ne
rect -13601 -15392 -12016 -14149
tri -17844 -16634 -16602 -15392 ne
rect -16602 -16634 -15016 -15392
tri -20844 -19462 -18016 -16634 ne
tri -18016 -18048 -16602 -16634 sw
tri -16602 -18048 -15188 -16634 ne
rect -15188 -16805 -15016 -16634
tri -15016 -16805 -13603 -15392 sw
tri -13601 -16805 -12188 -15392 ne
rect -12188 -15563 -12016 -15392
tri -12016 -15563 -10602 -14149 sw
tri -10602 -15563 -9188 -14149 ne
rect -9188 -14672 -8666 -14149
tri -8666 -14672 -7251 -13257 sw
tri -7251 -14500 -6008 -13257 ne
rect -6008 -14500 6008 -13257
tri 6008 -14500 7251 -13257 nw
tri 7251 -14672 8666 -13257 se
rect 8666 -13430 11321 -13257
tri 11321 -13430 12735 -12016 nw
tri 12735 -13430 14149 -12016 se
rect 14149 -12188 16805 -12016
tri 16805 -12188 16977 -12016 nw
tri 18220 -12188 19430 -10978 se
rect 19430 -12188 21048 -10978
tri 21048 -12188 22258 -10978 nw
rect 14149 -13430 15392 -12188
rect 8666 -14672 10079 -13430
tri 10079 -14672 11321 -13430 nw
rect -9188 -15500 -7251 -14672
tri -7251 -15500 -6423 -14672 sw
tri 6423 -15500 7251 -14672 se
rect 7251 -14844 9907 -14672
tri 9907 -14844 10079 -14672 nw
tri 11321 -14844 12735 -13430 se
rect 12735 -13601 15392 -13430
tri 15392 -13601 16805 -12188 nw
tri 16807 -13601 18220 -12188 se
rect 18220 -12360 20876 -12188
tri 20876 -12360 21048 -12188 nw
tri 22290 -12360 23672 -10978 se
rect 23672 -12360 25118 -10978
tri 25118 -12360 26500 -10978 nw
rect 18220 -13601 19462 -12360
rect 12735 -14844 14149 -13601
tri 14149 -14844 15392 -13601 nw
rect 7251 -15500 8493 -14844
rect -9188 -15563 -1085 -15500
rect -12188 -16805 -10602 -15563
rect -15188 -18048 -13603 -16805
rect -18016 -19462 -16602 -18048
tri -16602 -19462 -15188 -18048 sw
tri -15188 -18220 -15016 -18048 ne
rect -15016 -18220 -13603 -18048
tri -13603 -18220 -12188 -16805 sw
tri -12188 -16977 -12016 -16805 ne
rect -12016 -16977 -10602 -16805
tri -10602 -16977 -9188 -15563 sw
tri -9188 -16977 -7774 -15563 ne
rect -7774 -16977 -1085 -15563
tri -12016 -18220 -10773 -16977 ne
rect -10773 -17500 -9188 -16977
tri -9188 -17500 -8665 -16977 sw
tri -7774 -17500 -7251 -16977 ne
rect -7251 -17500 -1085 -16977
rect -10773 -18220 -8665 -17500
tri -15016 -19462 -13774 -18220 ne
rect -13774 -19257 -12188 -18220
tri -12188 -19257 -11151 -18220 sw
tri -10773 -19257 -9736 -18220 ne
rect -9736 -18500 -8665 -18220
tri -8665 -18500 -7665 -17500 sw
tri -1915 -17672 -1743 -17500 ne
rect -1743 -17672 -1085 -17500
tri -1085 -17672 1087 -15500 sw
tri 1732 -15747 1979 -15500 se
rect 1979 -15747 8493 -15500
rect 1732 -15849 8493 -15747
rect 1732 -16105 1832 -15849
rect 2088 -16105 2356 -15849
rect 2612 -16105 2910 -15849
rect 3166 -16105 3464 -15849
rect 3720 -16105 4018 -15849
rect 4274 -16105 4572 -15849
rect 4828 -16105 5126 -15849
rect 5382 -16105 5650 -15849
rect 5906 -16105 8493 -15849
rect 1732 -16258 8493 -16105
tri 8493 -16258 9907 -14844 nw
tri 9907 -16258 11321 -14844 se
rect 11321 -15016 13977 -14844
tri 13977 -15016 14149 -14844 nw
tri 15392 -15016 16807 -13601 se
rect 16807 -13774 19462 -13601
tri 19462 -13774 20876 -12360 nw
tri 20876 -13774 22290 -12360 se
rect 16807 -15016 18220 -13774
tri 18220 -15016 19462 -13774 nw
rect 11321 -16258 12564 -15016
rect 1732 -16373 7251 -16258
rect 1732 -16629 1832 -16373
rect 2088 -16629 2356 -16373
rect 2612 -16629 2910 -16373
rect 3166 -16629 3464 -16373
rect 3720 -16629 4018 -16373
rect 4274 -16629 4572 -16373
rect 4828 -16629 5126 -16373
rect 5382 -16629 5650 -16373
rect 5906 -16629 7251 -16373
rect 1732 -16897 7251 -16629
rect 1732 -17153 1832 -16897
rect 2088 -17153 2356 -16897
rect 2612 -17153 2910 -16897
rect 3166 -17153 3464 -16897
rect 3720 -17153 4018 -16897
rect 4274 -17153 4572 -16897
rect 4828 -17153 5126 -16897
rect 5382 -17153 5650 -16897
rect 5906 -17153 7251 -16897
rect 1732 -17253 7251 -17153
tri 1732 -17500 1979 -17253 ne
rect 1979 -17500 7251 -17253
tri 7251 -17500 8493 -16258 nw
tri 8493 -17672 9907 -16258 se
rect 9907 -16429 12564 -16258
tri 12564 -16429 13977 -15016 nw
tri 13979 -16429 15392 -15016 se
rect 15392 -15188 18048 -15016
tri 18048 -15188 18220 -15016 nw
tri 19462 -15188 20876 -13774 se
rect 20876 -15188 22290 -13774
tri 22290 -15188 25118 -12360 nw
rect 15392 -16429 16634 -15188
rect 9907 -17672 11321 -16429
tri 11321 -17672 12564 -16429 nw
rect -9736 -18747 -2202 -18500
tri -2202 -18747 -1955 -18500 sw
rect -9736 -18848 -1955 -18747
rect -9736 -19104 -6130 -18848
rect -5874 -19104 -5606 -18848
rect -5350 -19104 -5052 -18848
rect -4796 -19104 -4498 -18848
rect -4242 -19104 -3944 -18848
rect -3688 -19104 -3390 -18848
rect -3134 -19104 -2836 -18848
rect -2580 -19104 -2312 -18848
rect -2056 -19104 -1955 -18848
rect -9736 -19257 -1955 -19104
rect -13774 -19462 -11151 -19257
tri -18016 -22290 -15188 -19462 ne
tri -15188 -20876 -13774 -19462 sw
tri -13774 -20876 -12360 -19462 ne
rect -12360 -20672 -11151 -19462
tri -11151 -20672 -9736 -19257 sw
tri -9736 -20500 -8493 -19257 ne
rect -8493 -19372 -1955 -19257
rect -8493 -19628 -6130 -19372
rect -5874 -19628 -5606 -19372
rect -5350 -19628 -5052 -19372
rect -4796 -19628 -4498 -19372
rect -4242 -19628 -3944 -19372
rect -3688 -19628 -3390 -19372
rect -3134 -19628 -2836 -19372
rect -2580 -19628 -2312 -19372
rect -2056 -19628 -1955 -19372
rect -8493 -19896 -1955 -19628
rect -8493 -20152 -6130 -19896
rect -5874 -20152 -5606 -19896
rect -5350 -20152 -5052 -19896
rect -4796 -20152 -4498 -19896
rect -4242 -20152 -3944 -19896
rect -3688 -20152 -3390 -19896
rect -3134 -20152 -2836 -19896
rect -2580 -20152 -2312 -19896
rect -2056 -20152 -1955 -19896
rect -8493 -20253 -1955 -20152
rect -8493 -20500 -2202 -20253
tri -2202 -20500 -1955 -20253 nw
tri -1743 -20500 1085 -17672 ne
rect 1085 -18500 1087 -17672
tri 1087 -18500 1915 -17672 sw
tri 7665 -18500 8493 -17672 se
rect 8493 -17844 11149 -17672
tri 11149 -17844 11321 -17672 nw
tri 12564 -17844 13979 -16429 se
rect 13979 -16602 16634 -16429
tri 16634 -16602 18048 -15188 nw
tri 18048 -16602 19462 -15188 se
rect 13979 -17844 15392 -16602
tri 15392 -17844 16634 -16602 nw
rect 8493 -18500 9736 -17844
rect 1085 -19257 9736 -18500
tri 9736 -19257 11149 -17844 nw
tri 11151 -19257 12564 -17844 se
rect 12564 -18016 15220 -17844
tri 15220 -18016 15392 -17844 nw
tri 16634 -18016 18048 -16602 se
rect 18048 -18016 19462 -16602
tri 19462 -18016 22290 -15188 nw
rect 12564 -19257 13806 -18016
rect 1085 -20500 8493 -19257
tri 8493 -20500 9736 -19257 nw
tri 9736 -20672 11151 -19257 se
rect 11151 -19430 13806 -19257
tri 13806 -19430 15220 -18016 nw
tri 15220 -19430 16634 -18016 se
rect 11151 -20672 12564 -19430
tri 12564 -20672 13806 -19430 nw
rect -12360 -20876 -9736 -20672
rect -15188 -22290 -13774 -20876
tri -13774 -22290 -12360 -20876 sw
tri -12360 -22290 -10946 -20876 ne
rect -10946 -21500 -9736 -20876
tri -9736 -21500 -8908 -20672 sw
tri 8908 -21500 9736 -20672 se
rect 9736 -20844 12392 -20672
tri 12392 -20844 12564 -20672 nw
tri 13806 -20844 15220 -19430 se
rect 15220 -20844 16634 -19430
tri 16634 -20844 19462 -18016 nw
rect 9736 -21500 10978 -20844
rect -10946 -22290 -1085 -21500
tri -15188 -25118 -12360 -22290 ne
tri -12360 -23670 -10980 -22290 sw
tri -10946 -23500 -9736 -22290 ne
rect -9736 -23500 -1085 -22290
tri -1915 -23670 -1745 -23500 ne
rect -1745 -23670 -1085 -23500
tri -1085 -23670 1085 -21500 sw
tri 1732 -21747 1979 -21500 se
rect 1979 -21747 10978 -21500
rect 1732 -21848 10978 -21747
rect 1732 -22104 1833 -21848
rect 2089 -22104 2357 -21848
rect 2613 -22104 2911 -21848
rect 3167 -22104 3465 -21848
rect 3721 -22104 4019 -21848
rect 4275 -22104 4573 -21848
rect 4829 -22104 5127 -21848
rect 5383 -22104 5651 -21848
rect 5907 -22104 10978 -21848
rect 1732 -22258 10978 -22104
tri 10978 -22258 12392 -20844 nw
tri 12392 -22258 13806 -20844 se
rect 1732 -22372 9736 -22258
rect 1732 -22628 1833 -22372
rect 2089 -22628 2357 -22372
rect 2613 -22628 2911 -22372
rect 3167 -22628 3465 -22372
rect 3721 -22628 4019 -22372
rect 4275 -22628 4573 -22372
rect 4829 -22628 5127 -22372
rect 5383 -22628 5651 -22372
rect 5907 -22628 9736 -22372
rect 1732 -22896 9736 -22628
rect 1732 -23152 1833 -22896
rect 2089 -23152 2357 -22896
rect 2613 -23152 2911 -22896
rect 3167 -23152 3465 -22896
rect 3721 -23152 4019 -22896
rect 4275 -23152 4573 -22896
rect 4829 -23152 5127 -22896
rect 5383 -23152 5651 -22896
rect 5907 -23152 9736 -22896
rect 1732 -23253 9736 -23152
tri 1732 -23500 1979 -23253 ne
rect 1979 -23500 9736 -23253
tri 9736 -23500 10978 -22258 nw
rect -12360 -24500 -10980 -23670
tri -10980 -24500 -10150 -23670 sw
rect -12360 -24747 -2202 -24500
tri -2202 -24747 -1955 -24500 sw
rect -12360 -24848 -1955 -24747
rect -12360 -25104 -6130 -24848
rect -5874 -25104 -5606 -24848
rect -5350 -25104 -5052 -24848
rect -4796 -25104 -4498 -24848
rect -4242 -25104 -3944 -24848
rect -3688 -25104 -3390 -24848
rect -3134 -25104 -2836 -24848
rect -2580 -25104 -2312 -24848
rect -2056 -25104 -1955 -24848
rect -12360 -25118 -1955 -25104
tri -12360 -26500 -10978 -25118 ne
rect -10978 -25372 -1955 -25118
rect -10978 -25628 -6130 -25372
rect -5874 -25628 -5606 -25372
rect -5350 -25628 -5052 -25372
rect -4796 -25628 -4498 -25372
rect -4242 -25628 -3944 -25372
rect -3688 -25628 -3390 -25372
rect -3134 -25628 -2836 -25372
rect -2580 -25628 -2312 -25372
rect -2056 -25628 -1955 -25372
rect -10978 -25896 -1955 -25628
rect -10978 -26152 -6130 -25896
rect -5874 -26152 -5606 -25896
rect -5350 -26152 -5052 -25896
rect -4796 -26152 -4498 -25896
rect -4242 -26152 -3944 -25896
rect -3688 -26152 -3390 -25896
rect -3134 -26152 -2836 -25896
rect -2580 -26152 -2312 -25896
rect -2056 -26152 -1955 -25896
rect -10978 -26253 -1955 -26152
rect -10978 -26500 -2202 -26253
tri -2202 -26500 -1955 -26253 nw
tri -1745 -26500 1085 -23670 ne
tri 1085 -24500 1915 -23670 sw
tri 10978 -23672 12392 -22258 se
rect 12392 -23672 13806 -22258
tri 13806 -23672 16634 -20844 nw
tri 10150 -24500 10978 -23672 se
rect 1085 -26500 10978 -24500
tri 10978 -26500 13806 -23672 nw
<< comment >>
tri -10979 10979 -4549 26500 ne
rect -4549 10979 4549 26500
tri 4549 10980 10979 26500 nw
tri -26500 4549 -10979 10979 sw
tri -4549 4549 -1885 10979 ne
rect -1885 4549 1885 10979
tri 1885 4550 4549 10979 nw
tri 10979 4549 26500 10979 se
rect -26500 781 -10979 4549
tri -10979 781 -1885 4549 sw
tri -1885 781 -324 4549 ne
rect -324 781 324 4549
tri 324 782 1885 4549 nw
tri 1885 781 10979 4549 se
rect 10979 781 26500 4549
rect -26500 134 -1885 781
tri -1885 134 -324 781 sw
tri -324 134 -56 781 ne
rect -56 134 56 781
tri 56 135 324 781 nw
tri 324 134 1885 781 se
rect 1885 134 26500 781
rect -26500 23 -324 134
tri -324 23 -56 134 sw
tri -56 23 -10 134 ne
rect -10 23 10 134
tri 10 24 56 134 nw
tri 56 23 324 134 se
rect 324 23 26500 134
rect -26500 4 -56 23
tri -56 4 -10 23 sw
tri -10 4 -2 23 ne
rect -2 4 2 23
tri 2 5 10 23 nw
tri 10 4 56 23 se
rect 56 4 26500 23
rect -26500 1 -10 4
tri -10 1 -2 4 sw
tri -2 2 -1 4 ne
rect -1 1 1 4
tri 1 2 2 4 nw
tri 2 1 10 4 se
rect 10 1 26500 4
rect -26500 0 -2 1
tri -2 0 -1 1 sw
tri -1 0 0 1 ne
rect 0 0 26500 1
rect -26500 -1 -2 0
tri -2 -1 0 0 nw
tri 0 -1 1 0 ne
rect 1 -1 26500 0
rect -26500 -4 -10 -1
tri -10 -4 -2 -1 nw
tri -2 -4 0 -1 se
tri 0 -2 1 -1 sw
tri 2 -2 4 -1 ne
rect 4 -2 26500 -1
rect 0 -4 1 -2
rect -26500 -23 -56 -4
tri -56 -23 -10 -4 nw
tri -10 -23 -2 -5 se
rect -2 -10 1 -4
tri 1 -10 4 -2 sw
tri 4 -10 23 -2 ne
rect 23 -10 26500 -2
rect -2 -23 4 -10
rect -26500 -134 -324 -23
tri -324 -134 -56 -23 nw
tri -56 -134 -10 -24 se
rect -10 -56 4 -23
tri 4 -56 23 -10 sw
tri 23 -56 134 -10 ne
rect 134 -56 26500 -10
rect -10 -134 23 -56
rect -26500 -781 -1885 -134
tri -1885 -781 -324 -134 nw
tri -324 -781 -56 -135 se
rect -56 -324 23 -134
tri 23 -324 134 -56 sw
tri 134 -324 781 -56 ne
rect 781 -324 26500 -56
rect -56 -781 134 -324
rect -26500 -4549 -10979 -781
tri -10979 -4549 -1885 -781 nw
tri -1885 -4549 -324 -782 se
rect -324 -1885 134 -781
tri 134 -1885 781 -324 sw
tri 781 -1885 4549 -324 ne
rect 4549 -1885 26500 -324
rect -324 -4549 781 -1885
tri -26500 -10979 -10979 -4549 nw
tri -4549 -10979 -1885 -4550 se
rect -1885 -10979 781 -4549
tri 781 -10979 4549 -1885 sw
tri 4549 -10979 26500 -1885 ne
tri -10979 -26500 -4549 -10980 se
rect -4549 -26500 4549 -10979
tri 4549 -26500 10979 -10979 sw
<< properties >>
string GDS_END 10411040
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 10392572
string gencell sky130_fd_pr__rf_test_coil2
string library sky130
string parameter m=1
string path 637.500 -274.450 637.500 -75.000 
<< end >>
