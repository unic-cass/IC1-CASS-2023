magic
tech sky130A
magscale 1 2
timestamp 1676037725
<< locali >>
rect 165 1160 177 1194
rect 211 1160 249 1194
rect 283 1160 321 1194
rect 355 1160 393 1194
rect 427 1160 439 1194
rect 48 1020 82 1058
rect 48 948 82 986
rect 48 876 82 914
rect 48 804 82 842
rect 48 732 82 770
rect 48 660 82 698
rect 48 588 82 626
rect 48 516 82 554
rect 48 444 82 482
rect 48 372 82 410
rect 48 300 82 338
rect 48 228 82 266
rect 48 122 82 194
rect 522 1020 556 1058
rect 522 948 556 986
rect 522 876 556 914
rect 522 804 556 842
rect 522 732 556 770
rect 522 660 556 698
rect 522 588 556 626
rect 522 516 556 554
rect 522 444 556 482
rect 522 372 556 410
rect 522 300 556 338
rect 522 228 556 266
rect 522 122 556 194
rect 165 20 177 54
rect 211 20 249 54
rect 283 20 321 54
rect 355 20 393 54
rect 427 20 439 54
<< viali >>
rect 177 1160 211 1194
rect 249 1160 283 1194
rect 321 1160 355 1194
rect 393 1160 427 1194
rect 48 1058 82 1092
rect 48 986 82 1020
rect 48 914 82 948
rect 48 842 82 876
rect 48 770 82 804
rect 48 698 82 732
rect 48 626 82 660
rect 48 554 82 588
rect 48 482 82 516
rect 48 410 82 444
rect 48 338 82 372
rect 48 266 82 300
rect 48 194 82 228
rect 522 1058 556 1092
rect 522 986 556 1020
rect 522 914 556 948
rect 522 842 556 876
rect 522 770 556 804
rect 522 698 556 732
rect 522 626 556 660
rect 522 554 556 588
rect 522 482 556 516
rect 522 410 556 444
rect 522 338 556 372
rect 522 266 556 300
rect 522 194 556 228
rect 177 20 211 54
rect 249 20 283 54
rect 321 20 355 54
rect 393 20 427 54
<< obsli1 >>
rect 159 98 193 1116
rect 285 98 319 1116
rect 411 98 445 1116
<< metal1 >>
rect 165 1194 439 1214
rect 165 1160 177 1194
rect 211 1160 249 1194
rect 283 1160 321 1194
rect 355 1160 393 1194
rect 427 1160 439 1194
rect 165 1148 439 1160
rect 36 1092 94 1104
rect 36 1058 48 1092
rect 82 1058 94 1092
rect 36 1020 94 1058
rect 36 986 48 1020
rect 82 986 94 1020
rect 36 948 94 986
rect 36 914 48 948
rect 82 914 94 948
rect 36 876 94 914
rect 36 842 48 876
rect 82 842 94 876
rect 36 804 94 842
rect 36 770 48 804
rect 82 770 94 804
rect 36 732 94 770
rect 36 698 48 732
rect 82 698 94 732
rect 36 660 94 698
rect 36 626 48 660
rect 82 626 94 660
rect 36 588 94 626
rect 36 554 48 588
rect 82 554 94 588
rect 36 516 94 554
rect 36 482 48 516
rect 82 482 94 516
rect 36 444 94 482
rect 36 410 48 444
rect 82 410 94 444
rect 36 372 94 410
rect 36 338 48 372
rect 82 338 94 372
rect 36 300 94 338
rect 36 266 48 300
rect 82 266 94 300
rect 36 228 94 266
rect 36 194 48 228
rect 82 194 94 228
rect 36 110 94 194
rect 510 1092 568 1104
rect 510 1058 522 1092
rect 556 1058 568 1092
rect 510 1020 568 1058
rect 510 986 522 1020
rect 556 986 568 1020
rect 510 948 568 986
rect 510 914 522 948
rect 556 914 568 948
rect 510 876 568 914
rect 510 842 522 876
rect 556 842 568 876
rect 510 804 568 842
rect 510 770 522 804
rect 556 770 568 804
rect 510 732 568 770
rect 510 698 522 732
rect 556 698 568 732
rect 510 660 568 698
rect 510 626 522 660
rect 556 626 568 660
rect 510 588 568 626
rect 510 554 522 588
rect 556 554 568 588
rect 510 516 568 554
rect 510 482 522 516
rect 556 482 568 516
rect 510 444 568 482
rect 510 410 522 444
rect 556 410 568 444
rect 510 372 568 410
rect 510 338 522 372
rect 556 338 568 372
rect 510 300 568 338
rect 510 266 522 300
rect 556 266 568 300
rect 510 228 568 266
rect 510 194 522 228
rect 556 194 568 228
rect 510 110 568 194
rect 165 54 439 66
rect 165 20 177 54
rect 211 20 249 54
rect 283 20 321 54
rect 355 20 393 54
rect 427 20 439 54
rect 165 0 439 20
<< obsm1 >>
rect 150 110 202 1104
rect 276 110 328 1104
rect 402 110 454 1104
<< metal2 >>
rect 10 632 594 1104
rect 10 110 594 582
<< labels >>
rlabel viali s 522 1058 556 1092 6 BULK
port 1 nsew
rlabel viali s 522 986 556 1020 6 BULK
port 1 nsew
rlabel viali s 522 914 556 948 6 BULK
port 1 nsew
rlabel viali s 522 842 556 876 6 BULK
port 1 nsew
rlabel viali s 522 770 556 804 6 BULK
port 1 nsew
rlabel viali s 522 698 556 732 6 BULK
port 1 nsew
rlabel viali s 522 626 556 660 6 BULK
port 1 nsew
rlabel viali s 522 554 556 588 6 BULK
port 1 nsew
rlabel viali s 522 482 556 516 6 BULK
port 1 nsew
rlabel viali s 522 410 556 444 6 BULK
port 1 nsew
rlabel viali s 522 338 556 372 6 BULK
port 1 nsew
rlabel viali s 522 266 556 300 6 BULK
port 1 nsew
rlabel viali s 522 194 556 228 6 BULK
port 1 nsew
rlabel viali s 48 1058 82 1092 6 BULK
port 1 nsew
rlabel viali s 48 986 82 1020 6 BULK
port 1 nsew
rlabel viali s 48 914 82 948 6 BULK
port 1 nsew
rlabel viali s 48 842 82 876 6 BULK
port 1 nsew
rlabel viali s 48 770 82 804 6 BULK
port 1 nsew
rlabel viali s 48 698 82 732 6 BULK
port 1 nsew
rlabel viali s 48 626 82 660 6 BULK
port 1 nsew
rlabel viali s 48 554 82 588 6 BULK
port 1 nsew
rlabel viali s 48 482 82 516 6 BULK
port 1 nsew
rlabel viali s 48 410 82 444 6 BULK
port 1 nsew
rlabel viali s 48 338 82 372 6 BULK
port 1 nsew
rlabel viali s 48 266 82 300 6 BULK
port 1 nsew
rlabel viali s 48 194 82 228 6 BULK
port 1 nsew
rlabel locali s 522 122 556 1092 6 BULK
port 1 nsew
rlabel locali s 48 122 82 1092 6 BULK
port 1 nsew
rlabel metal1 s 510 110 568 1104 6 BULK
port 1 nsew
rlabel metal1 s 36 110 94 1104 6 BULK
port 1 nsew
rlabel metal2 s 10 632 594 1104 6 DRAIN
port 2 nsew
rlabel viali s 393 1160 427 1194 6 GATE
port 3 nsew
rlabel viali s 393 20 427 54 6 GATE
port 3 nsew
rlabel viali s 321 1160 355 1194 6 GATE
port 3 nsew
rlabel viali s 321 20 355 54 6 GATE
port 3 nsew
rlabel viali s 249 1160 283 1194 6 GATE
port 3 nsew
rlabel viali s 249 20 283 54 6 GATE
port 3 nsew
rlabel viali s 177 1160 211 1194 6 GATE
port 3 nsew
rlabel viali s 177 20 211 54 6 GATE
port 3 nsew
rlabel locali s 165 1160 439 1194 6 GATE
port 3 nsew
rlabel locali s 165 20 439 54 6 GATE
port 3 nsew
rlabel metal1 s 165 1148 439 1214 6 GATE
port 3 nsew
rlabel metal1 s 165 0 439 66 6 GATE
port 3 nsew
rlabel metal2 s 10 110 594 582 6 SOURCE
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 604 1214
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 9967686
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 9952034
<< end >>
