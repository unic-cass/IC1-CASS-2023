magic
tech sky130A
magscale 1 2
timestamp 1698801689
<< obsli1 >>
rect 1104 2159 51980 52785
<< obsm1 >>
rect 566 76 53070 52816
<< metal2 >>
rect 754 0 810 800
rect 2318 0 2374 800
rect 3882 0 3938 800
rect 5446 0 5502 800
rect 7010 0 7066 800
rect 8574 0 8630 800
rect 10138 0 10194 800
rect 11702 0 11758 800
rect 13266 0 13322 800
rect 14830 0 14886 800
rect 16394 0 16450 800
rect 17958 0 18014 800
rect 19522 0 19578 800
rect 21086 0 21142 800
rect 22650 0 22706 800
rect 24214 0 24270 800
rect 25778 0 25834 800
rect 27342 0 27398 800
rect 28906 0 28962 800
rect 30470 0 30526 800
rect 32034 0 32090 800
rect 33598 0 33654 800
rect 35162 0 35218 800
rect 36726 0 36782 800
rect 38290 0 38346 800
rect 39854 0 39910 800
rect 41418 0 41474 800
rect 42982 0 43038 800
rect 44546 0 44602 800
rect 46110 0 46166 800
rect 47674 0 47730 800
rect 49238 0 49294 800
rect 50802 0 50858 800
rect 52366 0 52422 800
<< obsm2 >>
rect 572 856 53144 52805
rect 572 70 698 856
rect 866 70 2262 856
rect 2430 70 3826 856
rect 3994 70 5390 856
rect 5558 70 6954 856
rect 7122 70 8518 856
rect 8686 70 10082 856
rect 10250 70 11646 856
rect 11814 70 13210 856
rect 13378 70 14774 856
rect 14942 70 16338 856
rect 16506 70 17902 856
rect 18070 70 19466 856
rect 19634 70 21030 856
rect 21198 70 22594 856
rect 22762 70 24158 856
rect 24326 70 25722 856
rect 25890 70 27286 856
rect 27454 70 28850 856
rect 29018 70 30414 856
rect 30582 70 31978 856
rect 32146 70 33542 856
rect 33710 70 35106 856
rect 35274 70 36670 856
rect 36838 70 38234 856
rect 38402 70 39798 856
rect 39966 70 41362 856
rect 41530 70 42926 856
rect 43094 70 44490 856
rect 44658 70 46054 856
rect 46222 70 47618 856
rect 47786 70 49182 856
rect 49350 70 50746 856
rect 50914 70 52310 856
rect 52478 70 53144 856
<< metal3 >>
rect 0 27480 800 27600
<< obsm3 >>
rect 749 27680 53071 52801
rect 880 27400 53071 27680
rect 749 851 53071 27400
<< metal4 >>
rect 4208 2128 4528 52816
rect 19568 2128 19888 52816
rect 34928 2128 35248 52816
rect 50288 2128 50608 52816
<< obsm4 >>
rect 979 2048 4128 47565
rect 4608 2048 19488 47565
rect 19968 2048 34848 47565
rect 35328 2048 50208 47565
rect 50688 2048 52381 47565
rect 979 851 52381 2048
<< labels >>
rlabel metal2 s 24214 0 24270 800 6 la_data_in_58_43[0]
port 1 nsew signal input
rlabel metal2 s 39854 0 39910 800 6 la_data_in_58_43[10]
port 2 nsew signal input
rlabel metal2 s 41418 0 41474 800 6 la_data_in_58_43[11]
port 3 nsew signal input
rlabel metal2 s 42982 0 43038 800 6 la_data_in_58_43[12]
port 4 nsew signal input
rlabel metal2 s 44546 0 44602 800 6 la_data_in_58_43[13]
port 5 nsew signal input
rlabel metal2 s 46110 0 46166 800 6 la_data_in_58_43[14]
port 6 nsew signal input
rlabel metal2 s 47674 0 47730 800 6 la_data_in_58_43[15]
port 7 nsew signal input
rlabel metal2 s 25778 0 25834 800 6 la_data_in_58_43[1]
port 8 nsew signal input
rlabel metal2 s 27342 0 27398 800 6 la_data_in_58_43[2]
port 9 nsew signal input
rlabel metal2 s 28906 0 28962 800 6 la_data_in_58_43[3]
port 10 nsew signal input
rlabel metal2 s 30470 0 30526 800 6 la_data_in_58_43[4]
port 11 nsew signal input
rlabel metal2 s 32034 0 32090 800 6 la_data_in_58_43[5]
port 12 nsew signal input
rlabel metal2 s 33598 0 33654 800 6 la_data_in_58_43[6]
port 13 nsew signal input
rlabel metal2 s 35162 0 35218 800 6 la_data_in_58_43[7]
port 14 nsew signal input
rlabel metal2 s 36726 0 36782 800 6 la_data_in_58_43[8]
port 15 nsew signal input
rlabel metal2 s 38290 0 38346 800 6 la_data_in_58_43[9]
port 16 nsew signal input
rlabel metal2 s 49238 0 49294 800 6 la_data_in_60_59[0]
port 17 nsew signal input
rlabel metal2 s 50802 0 50858 800 6 la_data_in_60_59[1]
port 18 nsew signal input
rlabel metal2 s 52366 0 52422 800 6 la_data_in_65
port 19 nsew signal input
rlabel metal2 s 754 0 810 800 6 la_data_out_23_16[0]
port 20 nsew signal output
rlabel metal2 s 2318 0 2374 800 6 la_data_out_23_16[1]
port 21 nsew signal output
rlabel metal2 s 3882 0 3938 800 6 la_data_out_23_16[2]
port 22 nsew signal output
rlabel metal2 s 5446 0 5502 800 6 la_data_out_23_16[3]
port 23 nsew signal output
rlabel metal2 s 7010 0 7066 800 6 la_data_out_23_16[4]
port 24 nsew signal output
rlabel metal2 s 8574 0 8630 800 6 la_data_out_23_16[5]
port 25 nsew signal output
rlabel metal2 s 10138 0 10194 800 6 la_data_out_23_16[6]
port 26 nsew signal output
rlabel metal2 s 11702 0 11758 800 6 la_data_out_23_16[7]
port 27 nsew signal output
rlabel metal2 s 13266 0 13322 800 6 la_data_out_26_24[0]
port 28 nsew signal output
rlabel metal2 s 14830 0 14886 800 6 la_data_out_26_24[1]
port 29 nsew signal output
rlabel metal2 s 16394 0 16450 800 6 la_data_out_26_24[2]
port 30 nsew signal output
rlabel metal2 s 17958 0 18014 800 6 la_data_out_30_27[0]
port 31 nsew signal output
rlabel metal2 s 19522 0 19578 800 6 la_data_out_30_27[1]
port 32 nsew signal output
rlabel metal2 s 21086 0 21142 800 6 la_data_out_30_27[2]
port 33 nsew signal output
rlabel metal2 s 22650 0 22706 800 6 la_data_out_30_27[3]
port 34 nsew signal output
rlabel metal4 s 4208 2128 4528 52816 6 vccd1
port 35 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 52816 6 vccd1
port 35 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 52816 6 vssd1
port 36 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 52816 6 vssd1
port 36 nsew ground bidirectional
rlabel metal3 s 0 27480 800 27600 6 wb_clk_i
port 37 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 53159 55303
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 11255716
string GDS_FILE /home/rodrigowue/IC1-V2/openlane/egd_top_wrapper/runs/23_10_31_22_11/results/signoff/egd_top_wrapper.magic.gds
string GDS_START 562642
<< end >>

