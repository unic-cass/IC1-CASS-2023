magic
tech sky130A
magscale 1 2
timestamp 1698545845
<< obsli1 >>
rect 1104 2159 558808 349809
<< obsm1 >>
rect 934 892 559070 349840
<< metal2 >>
rect 139950 351200 140006 352000
rect 419906 351200 419962 352000
rect 11702 0 11758 800
rect 34058 0 34114 800
rect 56414 0 56470 800
rect 78770 0 78826 800
rect 101126 0 101182 800
rect 123482 0 123538 800
rect 145838 0 145894 800
rect 168194 0 168250 800
rect 190550 0 190606 800
rect 212906 0 212962 800
rect 235262 0 235318 800
rect 257618 0 257674 800
rect 279974 0 280030 800
rect 302330 0 302386 800
rect 324686 0 324742 800
rect 347042 0 347098 800
rect 369398 0 369454 800
rect 391754 0 391810 800
rect 414110 0 414166 800
rect 436466 0 436522 800
rect 458822 0 458878 800
rect 481178 0 481234 800
rect 503534 0 503590 800
rect 525890 0 525946 800
rect 548246 0 548302 800
<< obsm2 >>
rect 938 351144 139894 351200
rect 140062 351144 419850 351200
rect 420018 351144 559066 351200
rect 938 856 559066 351144
rect 938 800 11646 856
rect 11814 800 34002 856
rect 34170 800 56358 856
rect 56526 800 78714 856
rect 78882 800 101070 856
rect 101238 800 123426 856
rect 123594 800 145782 856
rect 145950 800 168138 856
rect 168306 800 190494 856
rect 190662 800 212850 856
rect 213018 800 235206 856
rect 235374 800 257562 856
rect 257730 800 279918 856
rect 280086 800 302274 856
rect 302442 800 324630 856
rect 324798 800 346986 856
rect 347154 800 369342 856
rect 369510 800 391698 856
rect 391866 800 414054 856
rect 414222 800 436410 856
rect 436578 800 458766 856
rect 458934 800 481122 856
rect 481290 800 503478 856
rect 503646 800 525834 856
rect 526002 800 548190 856
rect 548358 800 559066 856
<< metal3 >>
rect 0 343816 800 343936
rect 0 340280 800 340400
rect 0 336744 800 336864
rect 0 333208 800 333328
rect 0 329672 800 329792
rect 0 326136 800 326256
rect 0 322600 800 322720
rect 0 319064 800 319184
rect 559200 316480 560000 316600
rect 0 315528 800 315648
rect 0 311992 800 312112
rect 0 308456 800 308576
rect 0 304920 800 305040
rect 0 301384 800 301504
rect 0 297848 800 297968
rect 0 294312 800 294432
rect 0 290776 800 290896
rect 0 287240 800 287360
rect 0 283704 800 283824
rect 0 280168 800 280288
rect 0 276632 800 276752
rect 0 273096 800 273216
rect 0 269560 800 269680
rect 0 266024 800 266144
rect 0 262488 800 262608
rect 0 258952 800 259072
rect 0 255416 800 255536
rect 0 251880 800 252000
rect 0 248344 800 248464
rect 559200 246168 560000 246288
rect 0 244808 800 244928
rect 0 241272 800 241392
rect 0 237736 800 237856
rect 0 234200 800 234320
rect 0 230664 800 230784
rect 0 227128 800 227248
rect 0 223592 800 223712
rect 0 220056 800 220176
rect 0 216520 800 216640
rect 0 212984 800 213104
rect 0 209448 800 209568
rect 0 205912 800 206032
rect 0 202376 800 202496
rect 0 198840 800 198960
rect 0 195304 800 195424
rect 0 191768 800 191888
rect 0 188232 800 188352
rect 0 184696 800 184816
rect 0 181160 800 181280
rect 0 177624 800 177744
rect 559200 175856 560000 175976
rect 0 174088 800 174208
rect 0 170552 800 170672
rect 0 167016 800 167136
rect 0 163480 800 163600
rect 0 159944 800 160064
rect 0 156408 800 156528
rect 0 152872 800 152992
rect 0 149336 800 149456
rect 0 145800 800 145920
rect 0 142264 800 142384
rect 0 138728 800 138848
rect 0 135192 800 135312
rect 0 131656 800 131776
rect 0 128120 800 128240
rect 0 124584 800 124704
rect 0 121048 800 121168
rect 0 117512 800 117632
rect 0 113976 800 114096
rect 0 110440 800 110560
rect 0 106904 800 107024
rect 559200 105544 560000 105664
rect 0 103368 800 103488
rect 0 99832 800 99952
rect 0 96296 800 96416
rect 0 92760 800 92880
rect 0 89224 800 89344
rect 0 85688 800 85808
rect 0 82152 800 82272
rect 0 78616 800 78736
rect 0 75080 800 75200
rect 0 71544 800 71664
rect 0 68008 800 68128
rect 0 64472 800 64592
rect 0 60936 800 61056
rect 0 57400 800 57520
rect 0 53864 800 53984
rect 0 50328 800 50448
rect 0 46792 800 46912
rect 0 43256 800 43376
rect 0 39720 800 39840
rect 0 36184 800 36304
rect 559200 35232 560000 35352
rect 0 32648 800 32768
rect 0 29112 800 29232
rect 0 25576 800 25696
rect 0 22040 800 22160
rect 0 18504 800 18624
rect 0 14968 800 15088
rect 0 11432 800 11552
rect 0 7896 800 8016
<< obsm3 >>
rect 800 344016 559200 349825
rect 880 343736 559200 344016
rect 800 340480 559200 343736
rect 880 340200 559200 340480
rect 800 336944 559200 340200
rect 880 336664 559200 336944
rect 800 333408 559200 336664
rect 880 333128 559200 333408
rect 800 329872 559200 333128
rect 880 329592 559200 329872
rect 800 326336 559200 329592
rect 880 326056 559200 326336
rect 800 322800 559200 326056
rect 880 322520 559200 322800
rect 800 319264 559200 322520
rect 880 318984 559200 319264
rect 800 316680 559200 318984
rect 800 316400 559120 316680
rect 800 315728 559200 316400
rect 880 315448 559200 315728
rect 800 312192 559200 315448
rect 880 311912 559200 312192
rect 800 308656 559200 311912
rect 880 308376 559200 308656
rect 800 305120 559200 308376
rect 880 304840 559200 305120
rect 800 301584 559200 304840
rect 880 301304 559200 301584
rect 800 298048 559200 301304
rect 880 297768 559200 298048
rect 800 294512 559200 297768
rect 880 294232 559200 294512
rect 800 290976 559200 294232
rect 880 290696 559200 290976
rect 800 287440 559200 290696
rect 880 287160 559200 287440
rect 800 283904 559200 287160
rect 880 283624 559200 283904
rect 800 280368 559200 283624
rect 880 280088 559200 280368
rect 800 276832 559200 280088
rect 880 276552 559200 276832
rect 800 273296 559200 276552
rect 880 273016 559200 273296
rect 800 269760 559200 273016
rect 880 269480 559200 269760
rect 800 266224 559200 269480
rect 880 265944 559200 266224
rect 800 262688 559200 265944
rect 880 262408 559200 262688
rect 800 259152 559200 262408
rect 880 258872 559200 259152
rect 800 255616 559200 258872
rect 880 255336 559200 255616
rect 800 252080 559200 255336
rect 880 251800 559200 252080
rect 800 248544 559200 251800
rect 880 248264 559200 248544
rect 800 246368 559200 248264
rect 800 246088 559120 246368
rect 800 245008 559200 246088
rect 880 244728 559200 245008
rect 800 241472 559200 244728
rect 880 241192 559200 241472
rect 800 237936 559200 241192
rect 880 237656 559200 237936
rect 800 234400 559200 237656
rect 880 234120 559200 234400
rect 800 230864 559200 234120
rect 880 230584 559200 230864
rect 800 227328 559200 230584
rect 880 227048 559200 227328
rect 800 223792 559200 227048
rect 880 223512 559200 223792
rect 800 220256 559200 223512
rect 880 219976 559200 220256
rect 800 216720 559200 219976
rect 880 216440 559200 216720
rect 800 213184 559200 216440
rect 880 212904 559200 213184
rect 800 209648 559200 212904
rect 880 209368 559200 209648
rect 800 206112 559200 209368
rect 880 205832 559200 206112
rect 800 202576 559200 205832
rect 880 202296 559200 202576
rect 800 199040 559200 202296
rect 880 198760 559200 199040
rect 800 195504 559200 198760
rect 880 195224 559200 195504
rect 800 191968 559200 195224
rect 880 191688 559200 191968
rect 800 188432 559200 191688
rect 880 188152 559200 188432
rect 800 184896 559200 188152
rect 880 184616 559200 184896
rect 800 181360 559200 184616
rect 880 181080 559200 181360
rect 800 177824 559200 181080
rect 880 177544 559200 177824
rect 800 176056 559200 177544
rect 800 175776 559120 176056
rect 800 174288 559200 175776
rect 880 174008 559200 174288
rect 800 170752 559200 174008
rect 880 170472 559200 170752
rect 800 167216 559200 170472
rect 880 166936 559200 167216
rect 800 163680 559200 166936
rect 880 163400 559200 163680
rect 800 160144 559200 163400
rect 880 159864 559200 160144
rect 800 156608 559200 159864
rect 880 156328 559200 156608
rect 800 153072 559200 156328
rect 880 152792 559200 153072
rect 800 149536 559200 152792
rect 880 149256 559200 149536
rect 800 146000 559200 149256
rect 880 145720 559200 146000
rect 800 142464 559200 145720
rect 880 142184 559200 142464
rect 800 138928 559200 142184
rect 880 138648 559200 138928
rect 800 135392 559200 138648
rect 880 135112 559200 135392
rect 800 131856 559200 135112
rect 880 131576 559200 131856
rect 800 128320 559200 131576
rect 880 128040 559200 128320
rect 800 124784 559200 128040
rect 880 124504 559200 124784
rect 800 121248 559200 124504
rect 880 120968 559200 121248
rect 800 117712 559200 120968
rect 880 117432 559200 117712
rect 800 114176 559200 117432
rect 880 113896 559200 114176
rect 800 110640 559200 113896
rect 880 110360 559200 110640
rect 800 107104 559200 110360
rect 880 106824 559200 107104
rect 800 105744 559200 106824
rect 800 105464 559120 105744
rect 800 103568 559200 105464
rect 880 103288 559200 103568
rect 800 100032 559200 103288
rect 880 99752 559200 100032
rect 800 96496 559200 99752
rect 880 96216 559200 96496
rect 800 92960 559200 96216
rect 880 92680 559200 92960
rect 800 89424 559200 92680
rect 880 89144 559200 89424
rect 800 85888 559200 89144
rect 880 85608 559200 85888
rect 800 82352 559200 85608
rect 880 82072 559200 82352
rect 800 78816 559200 82072
rect 880 78536 559200 78816
rect 800 75280 559200 78536
rect 880 75000 559200 75280
rect 800 71744 559200 75000
rect 880 71464 559200 71744
rect 800 68208 559200 71464
rect 880 67928 559200 68208
rect 800 64672 559200 67928
rect 880 64392 559200 64672
rect 800 61136 559200 64392
rect 880 60856 559200 61136
rect 800 57600 559200 60856
rect 880 57320 559200 57600
rect 800 54064 559200 57320
rect 880 53784 559200 54064
rect 800 50528 559200 53784
rect 880 50248 559200 50528
rect 800 46992 559200 50248
rect 880 46712 559200 46992
rect 800 43456 559200 46712
rect 880 43176 559200 43456
rect 800 39920 559200 43176
rect 880 39640 559200 39920
rect 800 36384 559200 39640
rect 880 36104 559200 36384
rect 800 35432 559200 36104
rect 800 35152 559120 35432
rect 800 32848 559200 35152
rect 880 32568 559200 32848
rect 800 29312 559200 32568
rect 880 29032 559200 29312
rect 800 25776 559200 29032
rect 880 25496 559200 25776
rect 800 22240 559200 25496
rect 880 21960 559200 22240
rect 800 18704 559200 21960
rect 880 18424 559200 18704
rect 800 15168 559200 18424
rect 880 14888 559200 15168
rect 800 11632 559200 14888
rect 880 11352 559200 11632
rect 800 8096 559200 11352
rect 880 7816 559200 8096
rect 800 2143 559200 7816
<< metal4 >>
rect 4208 2128 4528 349840
rect 19568 2128 19888 349840
rect 34928 2128 35248 349840
rect 50288 2128 50608 349840
rect 65648 2128 65968 349840
rect 81008 2128 81328 349840
rect 96368 2128 96688 349840
rect 111728 2128 112048 349840
rect 127088 2128 127408 349840
rect 142448 2128 142768 349840
rect 157808 2128 158128 349840
rect 173168 2128 173488 349840
rect 188528 2128 188848 349840
rect 203888 2128 204208 349840
rect 219248 2128 219568 349840
rect 234608 2128 234928 349840
rect 249968 2128 250288 349840
rect 265328 2128 265648 349840
rect 280688 2128 281008 349840
rect 296048 2128 296368 349840
rect 311408 2128 311728 349840
rect 326768 2128 327088 349840
rect 342128 2128 342448 349840
rect 357488 2128 357808 349840
rect 372848 2128 373168 349840
rect 388208 2128 388528 349840
rect 403568 2128 403888 349840
rect 418928 2128 419248 349840
rect 434288 2128 434608 349840
rect 449648 2128 449968 349840
rect 465008 2128 465328 349840
rect 480368 2128 480688 349840
rect 495728 2128 496048 349840
rect 511088 2128 511408 349840
rect 526448 2128 526768 349840
rect 541808 2128 542128 349840
rect 557168 2128 557488 349840
<< obsm4 >>
rect 1899 174523 4128 262989
rect 4608 174523 19488 262989
rect 19968 174523 34848 262989
rect 35328 174523 50208 262989
rect 50688 174523 65568 262989
rect 66048 174523 80928 262989
rect 81408 174523 96288 262989
rect 96768 174523 111648 262989
rect 112128 174523 127008 262989
rect 127488 174523 142368 262989
rect 142848 174523 157728 262989
rect 158208 174523 168485 262989
<< labels >>
rlabel metal2 s 11702 0 11758 800 6 buttons
port 1 nsew signal input
rlabel metal2 s 419906 351200 419962 352000 6 clk
port 2 nsew signal input
rlabel metal3 s 0 7896 800 8016 6 i_wb_addr[0]
port 3 nsew signal input
rlabel metal3 s 0 43256 800 43376 6 i_wb_addr[10]
port 4 nsew signal input
rlabel metal3 s 0 46792 800 46912 6 i_wb_addr[11]
port 5 nsew signal input
rlabel metal3 s 0 50328 800 50448 6 i_wb_addr[12]
port 6 nsew signal input
rlabel metal3 s 0 53864 800 53984 6 i_wb_addr[13]
port 7 nsew signal input
rlabel metal3 s 0 57400 800 57520 6 i_wb_addr[14]
port 8 nsew signal input
rlabel metal3 s 0 60936 800 61056 6 i_wb_addr[15]
port 9 nsew signal input
rlabel metal3 s 0 64472 800 64592 6 i_wb_addr[16]
port 10 nsew signal input
rlabel metal3 s 0 68008 800 68128 6 i_wb_addr[17]
port 11 nsew signal input
rlabel metal3 s 0 71544 800 71664 6 i_wb_addr[18]
port 12 nsew signal input
rlabel metal3 s 0 75080 800 75200 6 i_wb_addr[19]
port 13 nsew signal input
rlabel metal3 s 0 11432 800 11552 6 i_wb_addr[1]
port 14 nsew signal input
rlabel metal3 s 0 78616 800 78736 6 i_wb_addr[20]
port 15 nsew signal input
rlabel metal3 s 0 82152 800 82272 6 i_wb_addr[21]
port 16 nsew signal input
rlabel metal3 s 0 85688 800 85808 6 i_wb_addr[22]
port 17 nsew signal input
rlabel metal3 s 0 89224 800 89344 6 i_wb_addr[23]
port 18 nsew signal input
rlabel metal3 s 0 92760 800 92880 6 i_wb_addr[24]
port 19 nsew signal input
rlabel metal3 s 0 96296 800 96416 6 i_wb_addr[25]
port 20 nsew signal input
rlabel metal3 s 0 99832 800 99952 6 i_wb_addr[26]
port 21 nsew signal input
rlabel metal3 s 0 103368 800 103488 6 i_wb_addr[27]
port 22 nsew signal input
rlabel metal3 s 0 106904 800 107024 6 i_wb_addr[28]
port 23 nsew signal input
rlabel metal3 s 0 110440 800 110560 6 i_wb_addr[29]
port 24 nsew signal input
rlabel metal3 s 0 14968 800 15088 6 i_wb_addr[2]
port 25 nsew signal input
rlabel metal3 s 0 113976 800 114096 6 i_wb_addr[30]
port 26 nsew signal input
rlabel metal3 s 0 117512 800 117632 6 i_wb_addr[31]
port 27 nsew signal input
rlabel metal3 s 0 18504 800 18624 6 i_wb_addr[3]
port 28 nsew signal input
rlabel metal3 s 0 22040 800 22160 6 i_wb_addr[4]
port 29 nsew signal input
rlabel metal3 s 0 25576 800 25696 6 i_wb_addr[5]
port 30 nsew signal input
rlabel metal3 s 0 29112 800 29232 6 i_wb_addr[6]
port 31 nsew signal input
rlabel metal3 s 0 32648 800 32768 6 i_wb_addr[7]
port 32 nsew signal input
rlabel metal3 s 0 36184 800 36304 6 i_wb_addr[8]
port 33 nsew signal input
rlabel metal3 s 0 39720 800 39840 6 i_wb_addr[9]
port 34 nsew signal input
rlabel metal3 s 559200 35232 560000 35352 6 i_wb_cyc
port 35 nsew signal input
rlabel metal3 s 0 121048 800 121168 6 i_wb_data[0]
port 36 nsew signal input
rlabel metal3 s 0 156408 800 156528 6 i_wb_data[10]
port 37 nsew signal input
rlabel metal3 s 0 159944 800 160064 6 i_wb_data[11]
port 38 nsew signal input
rlabel metal3 s 0 163480 800 163600 6 i_wb_data[12]
port 39 nsew signal input
rlabel metal3 s 0 167016 800 167136 6 i_wb_data[13]
port 40 nsew signal input
rlabel metal3 s 0 170552 800 170672 6 i_wb_data[14]
port 41 nsew signal input
rlabel metal3 s 0 174088 800 174208 6 i_wb_data[15]
port 42 nsew signal input
rlabel metal3 s 0 177624 800 177744 6 i_wb_data[16]
port 43 nsew signal input
rlabel metal3 s 0 181160 800 181280 6 i_wb_data[17]
port 44 nsew signal input
rlabel metal3 s 0 184696 800 184816 6 i_wb_data[18]
port 45 nsew signal input
rlabel metal3 s 0 188232 800 188352 6 i_wb_data[19]
port 46 nsew signal input
rlabel metal3 s 0 124584 800 124704 6 i_wb_data[1]
port 47 nsew signal input
rlabel metal3 s 0 191768 800 191888 6 i_wb_data[20]
port 48 nsew signal input
rlabel metal3 s 0 195304 800 195424 6 i_wb_data[21]
port 49 nsew signal input
rlabel metal3 s 0 198840 800 198960 6 i_wb_data[22]
port 50 nsew signal input
rlabel metal3 s 0 202376 800 202496 6 i_wb_data[23]
port 51 nsew signal input
rlabel metal3 s 0 205912 800 206032 6 i_wb_data[24]
port 52 nsew signal input
rlabel metal3 s 0 209448 800 209568 6 i_wb_data[25]
port 53 nsew signal input
rlabel metal3 s 0 212984 800 213104 6 i_wb_data[26]
port 54 nsew signal input
rlabel metal3 s 0 216520 800 216640 6 i_wb_data[27]
port 55 nsew signal input
rlabel metal3 s 0 220056 800 220176 6 i_wb_data[28]
port 56 nsew signal input
rlabel metal3 s 0 223592 800 223712 6 i_wb_data[29]
port 57 nsew signal input
rlabel metal3 s 0 128120 800 128240 6 i_wb_data[2]
port 58 nsew signal input
rlabel metal3 s 0 227128 800 227248 6 i_wb_data[30]
port 59 nsew signal input
rlabel metal3 s 0 230664 800 230784 6 i_wb_data[31]
port 60 nsew signal input
rlabel metal3 s 0 131656 800 131776 6 i_wb_data[3]
port 61 nsew signal input
rlabel metal3 s 0 135192 800 135312 6 i_wb_data[4]
port 62 nsew signal input
rlabel metal3 s 0 138728 800 138848 6 i_wb_data[5]
port 63 nsew signal input
rlabel metal3 s 0 142264 800 142384 6 i_wb_data[6]
port 64 nsew signal input
rlabel metal3 s 0 145800 800 145920 6 i_wb_data[7]
port 65 nsew signal input
rlabel metal3 s 0 149336 800 149456 6 i_wb_data[8]
port 66 nsew signal input
rlabel metal3 s 0 152872 800 152992 6 i_wb_data[9]
port 67 nsew signal input
rlabel metal3 s 559200 105544 560000 105664 6 i_wb_stb
port 68 nsew signal input
rlabel metal3 s 559200 175856 560000 175976 6 i_wb_we
port 69 nsew signal input
rlabel metal2 s 34058 0 34114 800 6 led_enb[0]
port 70 nsew signal output
rlabel metal2 s 257618 0 257674 800 6 led_enb[10]
port 71 nsew signal output
rlabel metal2 s 279974 0 280030 800 6 led_enb[11]
port 72 nsew signal output
rlabel metal2 s 56414 0 56470 800 6 led_enb[1]
port 73 nsew signal output
rlabel metal2 s 78770 0 78826 800 6 led_enb[2]
port 74 nsew signal output
rlabel metal2 s 101126 0 101182 800 6 led_enb[3]
port 75 nsew signal output
rlabel metal2 s 123482 0 123538 800 6 led_enb[4]
port 76 nsew signal output
rlabel metal2 s 145838 0 145894 800 6 led_enb[5]
port 77 nsew signal output
rlabel metal2 s 168194 0 168250 800 6 led_enb[6]
port 78 nsew signal output
rlabel metal2 s 190550 0 190606 800 6 led_enb[7]
port 79 nsew signal output
rlabel metal2 s 212906 0 212962 800 6 led_enb[8]
port 80 nsew signal output
rlabel metal2 s 235262 0 235318 800 6 led_enb[9]
port 81 nsew signal output
rlabel metal2 s 302330 0 302386 800 6 leds[0]
port 82 nsew signal output
rlabel metal2 s 525890 0 525946 800 6 leds[10]
port 83 nsew signal output
rlabel metal2 s 548246 0 548302 800 6 leds[11]
port 84 nsew signal output
rlabel metal2 s 324686 0 324742 800 6 leds[1]
port 85 nsew signal output
rlabel metal2 s 347042 0 347098 800 6 leds[2]
port 86 nsew signal output
rlabel metal2 s 369398 0 369454 800 6 leds[3]
port 87 nsew signal output
rlabel metal2 s 391754 0 391810 800 6 leds[4]
port 88 nsew signal output
rlabel metal2 s 414110 0 414166 800 6 leds[5]
port 89 nsew signal output
rlabel metal2 s 436466 0 436522 800 6 leds[6]
port 90 nsew signal output
rlabel metal2 s 458822 0 458878 800 6 leds[7]
port 91 nsew signal output
rlabel metal2 s 481178 0 481234 800 6 leds[8]
port 92 nsew signal output
rlabel metal2 s 503534 0 503590 800 6 leds[9]
port 93 nsew signal output
rlabel metal3 s 559200 246168 560000 246288 6 o_wb_ack
port 94 nsew signal output
rlabel metal3 s 0 234200 800 234320 6 o_wb_data[0]
port 95 nsew signal output
rlabel metal3 s 0 269560 800 269680 6 o_wb_data[10]
port 96 nsew signal output
rlabel metal3 s 0 273096 800 273216 6 o_wb_data[11]
port 97 nsew signal output
rlabel metal3 s 0 276632 800 276752 6 o_wb_data[12]
port 98 nsew signal output
rlabel metal3 s 0 280168 800 280288 6 o_wb_data[13]
port 99 nsew signal output
rlabel metal3 s 0 283704 800 283824 6 o_wb_data[14]
port 100 nsew signal output
rlabel metal3 s 0 287240 800 287360 6 o_wb_data[15]
port 101 nsew signal output
rlabel metal3 s 0 290776 800 290896 6 o_wb_data[16]
port 102 nsew signal output
rlabel metal3 s 0 294312 800 294432 6 o_wb_data[17]
port 103 nsew signal output
rlabel metal3 s 0 297848 800 297968 6 o_wb_data[18]
port 104 nsew signal output
rlabel metal3 s 0 301384 800 301504 6 o_wb_data[19]
port 105 nsew signal output
rlabel metal3 s 0 237736 800 237856 6 o_wb_data[1]
port 106 nsew signal output
rlabel metal3 s 0 304920 800 305040 6 o_wb_data[20]
port 107 nsew signal output
rlabel metal3 s 0 308456 800 308576 6 o_wb_data[21]
port 108 nsew signal output
rlabel metal3 s 0 311992 800 312112 6 o_wb_data[22]
port 109 nsew signal output
rlabel metal3 s 0 315528 800 315648 6 o_wb_data[23]
port 110 nsew signal output
rlabel metal3 s 0 319064 800 319184 6 o_wb_data[24]
port 111 nsew signal output
rlabel metal3 s 0 322600 800 322720 6 o_wb_data[25]
port 112 nsew signal output
rlabel metal3 s 0 326136 800 326256 6 o_wb_data[26]
port 113 nsew signal output
rlabel metal3 s 0 329672 800 329792 6 o_wb_data[27]
port 114 nsew signal output
rlabel metal3 s 0 333208 800 333328 6 o_wb_data[28]
port 115 nsew signal output
rlabel metal3 s 0 336744 800 336864 6 o_wb_data[29]
port 116 nsew signal output
rlabel metal3 s 0 241272 800 241392 6 o_wb_data[2]
port 117 nsew signal output
rlabel metal3 s 0 340280 800 340400 6 o_wb_data[30]
port 118 nsew signal output
rlabel metal3 s 0 343816 800 343936 6 o_wb_data[31]
port 119 nsew signal output
rlabel metal3 s 0 244808 800 244928 6 o_wb_data[3]
port 120 nsew signal output
rlabel metal3 s 0 248344 800 248464 6 o_wb_data[4]
port 121 nsew signal output
rlabel metal3 s 0 251880 800 252000 6 o_wb_data[5]
port 122 nsew signal output
rlabel metal3 s 0 255416 800 255536 6 o_wb_data[6]
port 123 nsew signal output
rlabel metal3 s 0 258952 800 259072 6 o_wb_data[7]
port 124 nsew signal output
rlabel metal3 s 0 262488 800 262608 6 o_wb_data[8]
port 125 nsew signal output
rlabel metal3 s 0 266024 800 266144 6 o_wb_data[9]
port 126 nsew signal output
rlabel metal3 s 559200 316480 560000 316600 6 o_wb_stall
port 127 nsew signal output
rlabel metal2 s 139950 351200 140006 352000 6 reset
port 128 nsew signal input
rlabel metal4 s 4208 2128 4528 349840 6 vccd1
port 129 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 349840 6 vccd1
port 129 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 349840 6 vccd1
port 129 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 349840 6 vccd1
port 129 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 349840 6 vccd1
port 129 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 349840 6 vccd1
port 129 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 349840 6 vccd1
port 129 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 349840 6 vccd1
port 129 nsew power bidirectional
rlabel metal4 s 249968 2128 250288 349840 6 vccd1
port 129 nsew power bidirectional
rlabel metal4 s 280688 2128 281008 349840 6 vccd1
port 129 nsew power bidirectional
rlabel metal4 s 311408 2128 311728 349840 6 vccd1
port 129 nsew power bidirectional
rlabel metal4 s 342128 2128 342448 349840 6 vccd1
port 129 nsew power bidirectional
rlabel metal4 s 372848 2128 373168 349840 6 vccd1
port 129 nsew power bidirectional
rlabel metal4 s 403568 2128 403888 349840 6 vccd1
port 129 nsew power bidirectional
rlabel metal4 s 434288 2128 434608 349840 6 vccd1
port 129 nsew power bidirectional
rlabel metal4 s 465008 2128 465328 349840 6 vccd1
port 129 nsew power bidirectional
rlabel metal4 s 495728 2128 496048 349840 6 vccd1
port 129 nsew power bidirectional
rlabel metal4 s 526448 2128 526768 349840 6 vccd1
port 129 nsew power bidirectional
rlabel metal4 s 557168 2128 557488 349840 6 vccd1
port 129 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 349840 6 vssd1
port 130 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 349840 6 vssd1
port 130 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 349840 6 vssd1
port 130 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 349840 6 vssd1
port 130 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 349840 6 vssd1
port 130 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 349840 6 vssd1
port 130 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 349840 6 vssd1
port 130 nsew ground bidirectional
rlabel metal4 s 234608 2128 234928 349840 6 vssd1
port 130 nsew ground bidirectional
rlabel metal4 s 265328 2128 265648 349840 6 vssd1
port 130 nsew ground bidirectional
rlabel metal4 s 296048 2128 296368 349840 6 vssd1
port 130 nsew ground bidirectional
rlabel metal4 s 326768 2128 327088 349840 6 vssd1
port 130 nsew ground bidirectional
rlabel metal4 s 357488 2128 357808 349840 6 vssd1
port 130 nsew ground bidirectional
rlabel metal4 s 388208 2128 388528 349840 6 vssd1
port 130 nsew ground bidirectional
rlabel metal4 s 418928 2128 419248 349840 6 vssd1
port 130 nsew ground bidirectional
rlabel metal4 s 449648 2128 449968 349840 6 vssd1
port 130 nsew ground bidirectional
rlabel metal4 s 480368 2128 480688 349840 6 vssd1
port 130 nsew ground bidirectional
rlabel metal4 s 511088 2128 511408 349840 6 vssd1
port 130 nsew ground bidirectional
rlabel metal4 s 541808 2128 542128 349840 6 vssd1
port 130 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 560000 352000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 75313290
string GDS_FILE /home/bignixon/unic-cass/caravel_tutorial/caravel_user_project/openlane/wb_buttons_leds/runs/23_10_28_22_43/results/signoff/wb_buttons_leds.magic.gds
string GDS_START 1519226
<< end >>

