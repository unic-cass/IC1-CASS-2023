magic
tech sky130A
magscale 1 2
timestamp 1676037725
<< nwell >>
rect 2735 1206 3201 1878
rect -91 798 247 925
rect -91 166 817 798
rect 195 66 817 166
<< pwell >>
rect 1232 2195 2455 2228
rect 1232 2050 2563 2195
rect 4 1056 464 1308
rect 747 1056 2563 2050
rect 1225 1050 2563 1056
rect 1225 880 3126 1050
rect 917 798 3126 880
rect 917 102 2563 798
rect 917 66 1187 102
rect 2477 82 2563 102
<< nmos >>
rect 2679 824 2729 1024
rect 2785 824 2835 1024
rect 2891 824 2941 1024
rect 2997 824 3047 1024
<< mvnmos >>
rect 826 1424 946 2024
rect 1002 1424 1122 2024
rect 86 1082 206 1282
rect 262 1082 382 1282
rect 826 1082 946 1222
rect 1002 1082 1122 1222
rect 1311 1202 1411 2202
rect 1620 1202 1720 2202
<< mvpmos >>
rect 28 659 128 859
rect 28 232 128 432
rect 314 132 414 732
rect 470 132 570 732
<< mvnnmos >>
rect 1900 2002 2080 2202
rect 1900 1742 2080 1942
rect 1900 1482 2080 1682
rect 1900 1222 2080 1422
rect 1304 908 1484 1108
rect 1540 908 1720 1108
rect 1900 908 2080 1108
rect 1304 648 1484 848
rect 1540 648 1720 848
rect 1900 648 2080 848
rect 1304 388 1484 588
rect 1540 388 1720 588
rect 1900 388 2080 588
rect 1304 128 1484 328
rect 1540 128 1720 328
rect 1900 128 2080 328
<< pmoshvt >>
rect 2824 1242 2874 1842
rect 2930 1242 2980 1842
<< nmoslvt >>
rect 2260 2002 2290 2202
rect 2346 2002 2376 2202
rect 2260 1742 2290 1942
rect 2346 1742 2376 1942
rect 2260 1482 2290 1682
rect 2346 1482 2376 1682
rect 2260 1222 2290 1422
rect 2346 1222 2376 1422
rect 2260 908 2290 1108
rect 2346 908 2376 1108
rect 2260 648 2290 848
rect 2346 648 2376 848
rect 2260 388 2290 588
rect 2346 388 2376 588
rect 2260 128 2290 328
rect 2346 128 2376 328
<< ndiff >>
rect 2207 2184 2260 2202
rect 2207 2150 2215 2184
rect 2249 2150 2260 2184
rect 2207 2116 2260 2150
rect 2207 2082 2215 2116
rect 2249 2082 2260 2116
rect 2207 2048 2260 2082
rect 2207 2014 2215 2048
rect 2249 2014 2260 2048
rect 2207 2002 2260 2014
rect 2290 2184 2346 2202
rect 2290 2150 2301 2184
rect 2335 2150 2346 2184
rect 2290 2116 2346 2150
rect 2290 2082 2301 2116
rect 2335 2082 2346 2116
rect 2290 2048 2346 2082
rect 2290 2014 2301 2048
rect 2335 2014 2346 2048
rect 2290 2002 2346 2014
rect 2376 2184 2429 2202
rect 2376 2150 2387 2184
rect 2421 2150 2429 2184
rect 2376 2116 2429 2150
rect 2376 2082 2387 2116
rect 2421 2082 2429 2116
rect 2376 2048 2429 2082
rect 2376 2014 2387 2048
rect 2421 2014 2429 2048
rect 2376 2002 2429 2014
rect 2207 1924 2260 1942
rect 2207 1890 2215 1924
rect 2249 1890 2260 1924
rect 2207 1856 2260 1890
rect 2207 1822 2215 1856
rect 2249 1822 2260 1856
rect 2207 1788 2260 1822
rect 2207 1754 2215 1788
rect 2249 1754 2260 1788
rect 2207 1742 2260 1754
rect 2290 1924 2346 1942
rect 2290 1890 2301 1924
rect 2335 1890 2346 1924
rect 2290 1856 2346 1890
rect 2290 1822 2301 1856
rect 2335 1822 2346 1856
rect 2290 1788 2346 1822
rect 2290 1754 2301 1788
rect 2335 1754 2346 1788
rect 2290 1742 2346 1754
rect 2376 1924 2429 1942
rect 2376 1890 2387 1924
rect 2421 1890 2429 1924
rect 2376 1856 2429 1890
rect 2376 1822 2387 1856
rect 2421 1822 2429 1856
rect 2376 1788 2429 1822
rect 2376 1754 2387 1788
rect 2421 1754 2429 1788
rect 2376 1742 2429 1754
rect 2207 1664 2260 1682
rect 2207 1630 2215 1664
rect 2249 1630 2260 1664
rect 2207 1596 2260 1630
rect 2207 1562 2215 1596
rect 2249 1562 2260 1596
rect 2207 1528 2260 1562
rect 2207 1494 2215 1528
rect 2249 1494 2260 1528
rect 2207 1482 2260 1494
rect 2290 1664 2346 1682
rect 2290 1630 2301 1664
rect 2335 1630 2346 1664
rect 2290 1596 2346 1630
rect 2290 1562 2301 1596
rect 2335 1562 2346 1596
rect 2290 1528 2346 1562
rect 2290 1494 2301 1528
rect 2335 1494 2346 1528
rect 2290 1482 2346 1494
rect 2376 1664 2429 1682
rect 2376 1630 2387 1664
rect 2421 1630 2429 1664
rect 2376 1596 2429 1630
rect 2376 1562 2387 1596
rect 2421 1562 2429 1596
rect 2376 1528 2429 1562
rect 2376 1494 2387 1528
rect 2421 1494 2429 1528
rect 2376 1482 2429 1494
rect 2207 1404 2260 1422
rect 2207 1370 2215 1404
rect 2249 1370 2260 1404
rect 2207 1336 2260 1370
rect 2207 1302 2215 1336
rect 2249 1302 2260 1336
rect 2207 1268 2260 1302
rect 2207 1234 2215 1268
rect 2249 1234 2260 1268
rect 2207 1222 2260 1234
rect 2290 1404 2346 1422
rect 2290 1370 2301 1404
rect 2335 1370 2346 1404
rect 2290 1336 2346 1370
rect 2290 1302 2301 1336
rect 2335 1302 2346 1336
rect 2290 1268 2346 1302
rect 2290 1234 2301 1268
rect 2335 1234 2346 1268
rect 2290 1222 2346 1234
rect 2376 1404 2429 1422
rect 2376 1370 2387 1404
rect 2421 1370 2429 1404
rect 2376 1336 2429 1370
rect 2376 1302 2387 1336
rect 2421 1302 2429 1336
rect 2376 1268 2429 1302
rect 2376 1234 2387 1268
rect 2421 1234 2429 1268
rect 2376 1222 2429 1234
rect 2207 1090 2260 1108
rect 2207 1056 2215 1090
rect 2249 1056 2260 1090
rect 2207 1022 2260 1056
rect 2207 988 2215 1022
rect 2249 988 2260 1022
rect 2207 954 2260 988
rect 2207 920 2215 954
rect 2249 920 2260 954
rect 2207 908 2260 920
rect 2290 1090 2346 1108
rect 2290 1056 2301 1090
rect 2335 1056 2346 1090
rect 2290 1022 2346 1056
rect 2290 988 2301 1022
rect 2335 988 2346 1022
rect 2290 954 2346 988
rect 2290 920 2301 954
rect 2335 920 2346 954
rect 2290 908 2346 920
rect 2376 1090 2429 1108
rect 2376 1056 2387 1090
rect 2421 1056 2429 1090
rect 2376 1022 2429 1056
rect 2376 988 2387 1022
rect 2421 988 2429 1022
rect 2376 954 2429 988
rect 2376 920 2387 954
rect 2421 920 2429 954
rect 2376 908 2429 920
rect 2207 830 2260 848
rect 2207 796 2215 830
rect 2249 796 2260 830
rect 2207 762 2260 796
rect 2207 728 2215 762
rect 2249 728 2260 762
rect 2207 694 2260 728
rect 2207 660 2215 694
rect 2249 660 2260 694
rect 2207 648 2260 660
rect 2290 830 2346 848
rect 2290 796 2301 830
rect 2335 796 2346 830
rect 2290 762 2346 796
rect 2290 728 2301 762
rect 2335 728 2346 762
rect 2290 694 2346 728
rect 2290 660 2301 694
rect 2335 660 2346 694
rect 2290 648 2346 660
rect 2376 830 2429 848
rect 2376 796 2387 830
rect 2421 796 2429 830
rect 2376 762 2429 796
rect 2376 728 2387 762
rect 2421 728 2429 762
rect 2376 694 2429 728
rect 2376 660 2387 694
rect 2421 660 2429 694
rect 2376 648 2429 660
rect 2626 1006 2679 1024
rect 2626 972 2634 1006
rect 2668 972 2679 1006
rect 2626 938 2679 972
rect 2626 904 2634 938
rect 2668 904 2679 938
rect 2626 870 2679 904
rect 2626 836 2634 870
rect 2668 836 2679 870
rect 2626 824 2679 836
rect 2729 1006 2785 1024
rect 2729 972 2740 1006
rect 2774 972 2785 1006
rect 2729 938 2785 972
rect 2729 904 2740 938
rect 2774 904 2785 938
rect 2729 870 2785 904
rect 2729 836 2740 870
rect 2774 836 2785 870
rect 2729 824 2785 836
rect 2835 1006 2891 1024
rect 2835 972 2846 1006
rect 2880 972 2891 1006
rect 2835 938 2891 972
rect 2835 904 2846 938
rect 2880 904 2891 938
rect 2835 870 2891 904
rect 2835 836 2846 870
rect 2880 836 2891 870
rect 2835 824 2891 836
rect 2941 1006 2997 1024
rect 2941 972 2952 1006
rect 2986 972 2997 1006
rect 2941 938 2997 972
rect 2941 904 2952 938
rect 2986 904 2997 938
rect 2941 870 2997 904
rect 2941 836 2952 870
rect 2986 836 2997 870
rect 2941 824 2997 836
rect 3047 1006 3100 1024
rect 3047 972 3058 1006
rect 3092 972 3100 1006
rect 3047 938 3100 972
rect 3047 904 3058 938
rect 3092 904 3100 938
rect 3047 870 3100 904
rect 3047 836 3058 870
rect 3092 836 3100 870
rect 3047 824 3100 836
rect 2207 570 2260 588
rect 2207 536 2215 570
rect 2249 536 2260 570
rect 2207 502 2260 536
rect 2207 468 2215 502
rect 2249 468 2260 502
rect 2207 434 2260 468
rect 2207 400 2215 434
rect 2249 400 2260 434
rect 2207 388 2260 400
rect 2290 570 2346 588
rect 2290 536 2301 570
rect 2335 536 2346 570
rect 2290 502 2346 536
rect 2290 468 2301 502
rect 2335 468 2346 502
rect 2290 434 2346 468
rect 2290 400 2301 434
rect 2335 400 2346 434
rect 2290 388 2346 400
rect 2376 570 2429 588
rect 2376 536 2387 570
rect 2421 536 2429 570
rect 2376 502 2429 536
rect 2376 468 2387 502
rect 2421 468 2429 502
rect 2376 434 2429 468
rect 2376 400 2387 434
rect 2421 400 2429 434
rect 2376 388 2429 400
rect 2207 310 2260 328
rect 2207 276 2215 310
rect 2249 276 2260 310
rect 2207 242 2260 276
rect 2207 208 2215 242
rect 2249 208 2260 242
rect 2207 174 2260 208
rect 2207 140 2215 174
rect 2249 140 2260 174
rect 2207 128 2260 140
rect 2290 310 2346 328
rect 2290 276 2301 310
rect 2335 276 2346 310
rect 2290 242 2346 276
rect 2290 208 2301 242
rect 2335 208 2346 242
rect 2290 174 2346 208
rect 2290 140 2301 174
rect 2335 140 2346 174
rect 2290 128 2346 140
rect 2376 310 2429 328
rect 2376 276 2387 310
rect 2421 276 2429 310
rect 2376 242 2429 276
rect 2376 208 2387 242
rect 2421 208 2429 242
rect 2376 174 2429 208
rect 2376 140 2387 174
rect 2421 140 2429 174
rect 2376 128 2429 140
<< pdiff >>
rect 2771 1830 2824 1842
rect 2771 1796 2779 1830
rect 2813 1796 2824 1830
rect 2771 1762 2824 1796
rect 2771 1728 2779 1762
rect 2813 1728 2824 1762
rect 2771 1694 2824 1728
rect 2771 1660 2779 1694
rect 2813 1660 2824 1694
rect 2771 1626 2824 1660
rect 2771 1592 2779 1626
rect 2813 1592 2824 1626
rect 2771 1558 2824 1592
rect 2771 1524 2779 1558
rect 2813 1524 2824 1558
rect 2771 1490 2824 1524
rect 2771 1456 2779 1490
rect 2813 1456 2824 1490
rect 2771 1422 2824 1456
rect 2771 1388 2779 1422
rect 2813 1388 2824 1422
rect 2771 1354 2824 1388
rect 2771 1320 2779 1354
rect 2813 1320 2824 1354
rect 2771 1242 2824 1320
rect 2874 1830 2930 1842
rect 2874 1796 2885 1830
rect 2919 1796 2930 1830
rect 2874 1762 2930 1796
rect 2874 1728 2885 1762
rect 2919 1728 2930 1762
rect 2874 1694 2930 1728
rect 2874 1660 2885 1694
rect 2919 1660 2930 1694
rect 2874 1626 2930 1660
rect 2874 1592 2885 1626
rect 2919 1592 2930 1626
rect 2874 1558 2930 1592
rect 2874 1524 2885 1558
rect 2919 1524 2930 1558
rect 2874 1490 2930 1524
rect 2874 1456 2885 1490
rect 2919 1456 2930 1490
rect 2874 1422 2930 1456
rect 2874 1388 2885 1422
rect 2919 1388 2930 1422
rect 2874 1354 2930 1388
rect 2874 1320 2885 1354
rect 2919 1320 2930 1354
rect 2874 1242 2930 1320
rect 2980 1830 3033 1842
rect 2980 1796 2991 1830
rect 3025 1796 3033 1830
rect 2980 1762 3033 1796
rect 2980 1728 2991 1762
rect 3025 1728 3033 1762
rect 2980 1694 3033 1728
rect 2980 1660 2991 1694
rect 3025 1660 3033 1694
rect 2980 1626 3033 1660
rect 2980 1592 2991 1626
rect 3025 1592 3033 1626
rect 2980 1558 3033 1592
rect 2980 1524 2991 1558
rect 3025 1524 3033 1558
rect 2980 1490 3033 1524
rect 2980 1456 2991 1490
rect 3025 1456 3033 1490
rect 2980 1422 3033 1456
rect 2980 1388 2991 1422
rect 3025 1388 3033 1422
rect 2980 1354 3033 1388
rect 2980 1320 2991 1354
rect 3025 1320 3033 1354
rect 2980 1242 3033 1320
<< mvndiff >>
rect 1258 2190 1311 2202
rect 1258 2156 1266 2190
rect 1300 2156 1311 2190
rect 1258 2122 1311 2156
rect 1258 2088 1266 2122
rect 1300 2088 1311 2122
rect 1258 2054 1311 2088
rect 773 2012 826 2024
rect 773 1978 781 2012
rect 815 1978 826 2012
rect 773 1944 826 1978
rect 773 1910 781 1944
rect 815 1910 826 1944
rect 773 1876 826 1910
rect 773 1842 781 1876
rect 815 1842 826 1876
rect 773 1808 826 1842
rect 773 1774 781 1808
rect 815 1774 826 1808
rect 773 1740 826 1774
rect 773 1706 781 1740
rect 815 1706 826 1740
rect 773 1672 826 1706
rect 773 1638 781 1672
rect 815 1638 826 1672
rect 773 1604 826 1638
rect 773 1570 781 1604
rect 815 1570 826 1604
rect 773 1536 826 1570
rect 773 1502 781 1536
rect 815 1502 826 1536
rect 773 1424 826 1502
rect 946 2012 1002 2024
rect 946 1978 957 2012
rect 991 1978 1002 2012
rect 946 1944 1002 1978
rect 946 1910 957 1944
rect 991 1910 1002 1944
rect 946 1876 1002 1910
rect 946 1842 957 1876
rect 991 1842 1002 1876
rect 946 1808 1002 1842
rect 946 1774 957 1808
rect 991 1774 1002 1808
rect 946 1740 1002 1774
rect 946 1706 957 1740
rect 991 1706 1002 1740
rect 946 1672 1002 1706
rect 946 1638 957 1672
rect 991 1638 1002 1672
rect 946 1604 1002 1638
rect 946 1570 957 1604
rect 991 1570 1002 1604
rect 946 1536 1002 1570
rect 946 1502 957 1536
rect 991 1502 1002 1536
rect 946 1424 1002 1502
rect 1122 2012 1175 2024
rect 1122 1978 1133 2012
rect 1167 1978 1175 2012
rect 1122 1944 1175 1978
rect 1122 1910 1133 1944
rect 1167 1910 1175 1944
rect 1122 1876 1175 1910
rect 1122 1842 1133 1876
rect 1167 1842 1175 1876
rect 1122 1808 1175 1842
rect 1122 1774 1133 1808
rect 1167 1774 1175 1808
rect 1122 1740 1175 1774
rect 1122 1706 1133 1740
rect 1167 1706 1175 1740
rect 1122 1672 1175 1706
rect 1122 1638 1133 1672
rect 1167 1638 1175 1672
rect 1122 1604 1175 1638
rect 1122 1570 1133 1604
rect 1167 1570 1175 1604
rect 1122 1536 1175 1570
rect 1122 1502 1133 1536
rect 1167 1502 1175 1536
rect 1122 1424 1175 1502
rect 1258 2020 1266 2054
rect 1300 2020 1311 2054
rect 1258 1986 1311 2020
rect 1258 1952 1266 1986
rect 1300 1952 1311 1986
rect 1258 1918 1311 1952
rect 1258 1884 1266 1918
rect 1300 1884 1311 1918
rect 1258 1850 1311 1884
rect 1258 1816 1266 1850
rect 1300 1816 1311 1850
rect 1258 1782 1311 1816
rect 1258 1748 1266 1782
rect 1300 1748 1311 1782
rect 1258 1714 1311 1748
rect 1258 1680 1266 1714
rect 1300 1680 1311 1714
rect 1258 1646 1311 1680
rect 1258 1612 1266 1646
rect 1300 1612 1311 1646
rect 1258 1578 1311 1612
rect 1258 1544 1266 1578
rect 1300 1544 1311 1578
rect 1258 1510 1311 1544
rect 1258 1476 1266 1510
rect 1300 1476 1311 1510
rect 1258 1442 1311 1476
rect 1258 1408 1266 1442
rect 1300 1408 1311 1442
rect 1258 1374 1311 1408
rect 1258 1340 1266 1374
rect 1300 1340 1311 1374
rect 1258 1306 1311 1340
rect 30 1270 86 1282
rect 30 1236 41 1270
rect 75 1236 86 1270
rect 30 1202 86 1236
rect 30 1168 41 1202
rect 75 1168 86 1202
rect 30 1134 86 1168
rect 30 1100 41 1134
rect 75 1100 86 1134
rect 30 1082 86 1100
rect 206 1270 262 1282
rect 206 1236 217 1270
rect 251 1236 262 1270
rect 206 1202 262 1236
rect 206 1168 217 1202
rect 251 1168 262 1202
rect 206 1134 262 1168
rect 206 1100 217 1134
rect 251 1100 262 1134
rect 206 1082 262 1100
rect 382 1270 438 1282
rect 382 1236 393 1270
rect 427 1236 438 1270
rect 1258 1272 1266 1306
rect 1300 1272 1311 1306
rect 382 1202 438 1236
rect 382 1168 393 1202
rect 427 1168 438 1202
rect 382 1134 438 1168
rect 382 1100 393 1134
rect 427 1100 438 1134
rect 382 1082 438 1100
rect 773 1210 826 1222
rect 773 1176 781 1210
rect 815 1176 826 1210
rect 773 1142 826 1176
rect 773 1108 781 1142
rect 815 1108 826 1142
rect 773 1082 826 1108
rect 946 1210 1002 1222
rect 946 1176 957 1210
rect 991 1176 1002 1210
rect 946 1142 1002 1176
rect 946 1108 957 1142
rect 991 1108 1002 1142
rect 946 1082 1002 1108
rect 1122 1210 1175 1222
rect 1122 1176 1133 1210
rect 1167 1176 1175 1210
rect 1258 1202 1311 1272
rect 1411 2190 1467 2202
rect 1411 2156 1422 2190
rect 1456 2156 1467 2190
rect 1411 2122 1467 2156
rect 1411 2088 1422 2122
rect 1456 2088 1467 2122
rect 1411 2054 1467 2088
rect 1411 2020 1422 2054
rect 1456 2020 1467 2054
rect 1411 1986 1467 2020
rect 1411 1952 1422 1986
rect 1456 1952 1467 1986
rect 1411 1918 1467 1952
rect 1411 1884 1422 1918
rect 1456 1884 1467 1918
rect 1411 1850 1467 1884
rect 1411 1816 1422 1850
rect 1456 1816 1467 1850
rect 1411 1782 1467 1816
rect 1411 1748 1422 1782
rect 1456 1748 1467 1782
rect 1411 1714 1467 1748
rect 1411 1680 1422 1714
rect 1456 1680 1467 1714
rect 1411 1646 1467 1680
rect 1411 1612 1422 1646
rect 1456 1612 1467 1646
rect 1411 1578 1467 1612
rect 1411 1544 1422 1578
rect 1456 1544 1467 1578
rect 1411 1510 1467 1544
rect 1411 1476 1422 1510
rect 1456 1476 1467 1510
rect 1411 1442 1467 1476
rect 1411 1408 1422 1442
rect 1456 1408 1467 1442
rect 1411 1374 1467 1408
rect 1411 1340 1422 1374
rect 1456 1340 1467 1374
rect 1411 1306 1467 1340
rect 1411 1272 1422 1306
rect 1456 1272 1467 1306
rect 1411 1202 1467 1272
rect 1567 2190 1620 2202
rect 1567 2156 1575 2190
rect 1609 2156 1620 2190
rect 1567 2122 1620 2156
rect 1567 2088 1575 2122
rect 1609 2088 1620 2122
rect 1567 2054 1620 2088
rect 1567 2020 1575 2054
rect 1609 2020 1620 2054
rect 1567 1986 1620 2020
rect 1567 1952 1575 1986
rect 1609 1952 1620 1986
rect 1567 1918 1620 1952
rect 1567 1884 1575 1918
rect 1609 1884 1620 1918
rect 1567 1850 1620 1884
rect 1567 1816 1575 1850
rect 1609 1816 1620 1850
rect 1567 1782 1620 1816
rect 1567 1748 1575 1782
rect 1609 1748 1620 1782
rect 1567 1714 1620 1748
rect 1567 1680 1575 1714
rect 1609 1680 1620 1714
rect 1567 1646 1620 1680
rect 1567 1612 1575 1646
rect 1609 1612 1620 1646
rect 1567 1578 1620 1612
rect 1567 1544 1575 1578
rect 1609 1544 1620 1578
rect 1567 1510 1620 1544
rect 1567 1476 1575 1510
rect 1609 1476 1620 1510
rect 1567 1442 1620 1476
rect 1567 1408 1575 1442
rect 1609 1408 1620 1442
rect 1567 1374 1620 1408
rect 1567 1340 1575 1374
rect 1609 1340 1620 1374
rect 1567 1306 1620 1340
rect 1567 1272 1575 1306
rect 1609 1272 1620 1306
rect 1567 1202 1620 1272
rect 1720 2190 1773 2202
rect 1720 2156 1731 2190
rect 1765 2156 1773 2190
rect 1720 2122 1773 2156
rect 1720 2088 1731 2122
rect 1765 2088 1773 2122
rect 1720 2054 1773 2088
rect 1720 2020 1731 2054
rect 1765 2020 1773 2054
rect 1720 1986 1773 2020
rect 1847 2184 1900 2202
rect 1847 2150 1855 2184
rect 1889 2150 1900 2184
rect 1847 2116 1900 2150
rect 1847 2082 1855 2116
rect 1889 2082 1900 2116
rect 1847 2048 1900 2082
rect 1847 2014 1855 2048
rect 1889 2014 1900 2048
rect 1847 2002 1900 2014
rect 2080 2184 2133 2202
rect 2080 2150 2091 2184
rect 2125 2150 2133 2184
rect 2080 2116 2133 2150
rect 2080 2082 2091 2116
rect 2125 2082 2133 2116
rect 2080 2048 2133 2082
rect 2080 2014 2091 2048
rect 2125 2014 2133 2048
rect 2080 2002 2133 2014
rect 1720 1952 1731 1986
rect 1765 1952 1773 1986
rect 1720 1918 1773 1952
rect 1720 1884 1731 1918
rect 1765 1884 1773 1918
rect 1720 1850 1773 1884
rect 1720 1816 1731 1850
rect 1765 1816 1773 1850
rect 1720 1782 1773 1816
rect 1720 1748 1731 1782
rect 1765 1748 1773 1782
rect 1720 1714 1773 1748
rect 1847 1924 1900 1942
rect 1847 1890 1855 1924
rect 1889 1890 1900 1924
rect 1847 1856 1900 1890
rect 1847 1822 1855 1856
rect 1889 1822 1900 1856
rect 1847 1788 1900 1822
rect 1847 1754 1855 1788
rect 1889 1754 1900 1788
rect 1847 1742 1900 1754
rect 2080 1924 2133 1942
rect 2080 1890 2091 1924
rect 2125 1890 2133 1924
rect 2080 1856 2133 1890
rect 2080 1822 2091 1856
rect 2125 1822 2133 1856
rect 2080 1788 2133 1822
rect 2080 1754 2091 1788
rect 2125 1754 2133 1788
rect 2080 1742 2133 1754
rect 1720 1680 1731 1714
rect 1765 1680 1773 1714
rect 1720 1646 1773 1680
rect 1720 1612 1731 1646
rect 1765 1612 1773 1646
rect 1720 1578 1773 1612
rect 1720 1544 1731 1578
rect 1765 1544 1773 1578
rect 1720 1510 1773 1544
rect 1720 1476 1731 1510
rect 1765 1476 1773 1510
rect 1847 1664 1900 1682
rect 1847 1630 1855 1664
rect 1889 1630 1900 1664
rect 1847 1596 1900 1630
rect 1847 1562 1855 1596
rect 1889 1562 1900 1596
rect 1847 1528 1900 1562
rect 1847 1494 1855 1528
rect 1889 1494 1900 1528
rect 1847 1482 1900 1494
rect 2080 1664 2133 1682
rect 2080 1630 2091 1664
rect 2125 1630 2133 1664
rect 2080 1596 2133 1630
rect 2080 1562 2091 1596
rect 2125 1562 2133 1596
rect 2080 1528 2133 1562
rect 2080 1494 2091 1528
rect 2125 1494 2133 1528
rect 2080 1482 2133 1494
rect 1720 1442 1773 1476
rect 1720 1408 1731 1442
rect 1765 1408 1773 1442
rect 1720 1374 1773 1408
rect 1720 1340 1731 1374
rect 1765 1340 1773 1374
rect 1720 1306 1773 1340
rect 1720 1272 1731 1306
rect 1765 1272 1773 1306
rect 1720 1202 1773 1272
rect 1847 1404 1900 1422
rect 1847 1370 1855 1404
rect 1889 1370 1900 1404
rect 1847 1336 1900 1370
rect 1847 1302 1855 1336
rect 1889 1302 1900 1336
rect 1847 1268 1900 1302
rect 1847 1234 1855 1268
rect 1889 1234 1900 1268
rect 1847 1222 1900 1234
rect 2080 1404 2133 1422
rect 2080 1370 2091 1404
rect 2125 1370 2133 1404
rect 2080 1336 2133 1370
rect 2080 1302 2091 1336
rect 2125 1302 2133 1336
rect 2080 1268 2133 1302
rect 2080 1234 2091 1268
rect 2125 1234 2133 1268
rect 2080 1222 2133 1234
rect 1122 1142 1175 1176
rect 1122 1108 1133 1142
rect 1167 1108 1175 1142
rect 1122 1082 1175 1108
rect 1251 1090 1304 1108
rect 1251 1056 1259 1090
rect 1293 1056 1304 1090
rect 1251 1022 1304 1056
rect 1251 988 1259 1022
rect 1293 988 1304 1022
rect 1251 954 1304 988
rect 1251 920 1259 954
rect 1293 920 1304 954
rect 1251 908 1304 920
rect 1484 1090 1540 1108
rect 1484 1056 1495 1090
rect 1529 1056 1540 1090
rect 1484 1022 1540 1056
rect 1484 988 1495 1022
rect 1529 988 1540 1022
rect 1484 954 1540 988
rect 1484 920 1495 954
rect 1529 920 1540 954
rect 1484 908 1540 920
rect 1720 1090 1773 1108
rect 1720 1056 1731 1090
rect 1765 1056 1773 1090
rect 1720 1022 1773 1056
rect 1720 988 1731 1022
rect 1765 988 1773 1022
rect 1720 954 1773 988
rect 1720 920 1731 954
rect 1765 920 1773 954
rect 1720 908 1773 920
rect 1847 1090 1900 1108
rect 1847 1056 1855 1090
rect 1889 1056 1900 1090
rect 1847 1022 1900 1056
rect 1847 988 1855 1022
rect 1889 988 1900 1022
rect 1847 954 1900 988
rect 1847 920 1855 954
rect 1889 920 1900 954
rect 1847 908 1900 920
rect 2080 1090 2133 1108
rect 2080 1056 2091 1090
rect 2125 1056 2133 1090
rect 2080 1022 2133 1056
rect 2080 988 2091 1022
rect 2125 988 2133 1022
rect 2080 954 2133 988
rect 2080 920 2091 954
rect 2125 920 2133 954
rect 2080 908 2133 920
rect 1251 830 1304 848
rect 1251 796 1259 830
rect 1293 796 1304 830
rect 1251 762 1304 796
rect 1251 728 1259 762
rect 1293 728 1304 762
rect 1251 694 1304 728
rect 1251 660 1259 694
rect 1293 660 1304 694
rect 1251 648 1304 660
rect 1484 830 1540 848
rect 1484 796 1495 830
rect 1529 796 1540 830
rect 1484 762 1540 796
rect 1484 728 1495 762
rect 1529 728 1540 762
rect 1484 694 1540 728
rect 1484 660 1495 694
rect 1529 660 1540 694
rect 1484 648 1540 660
rect 1720 830 1773 848
rect 1720 796 1731 830
rect 1765 796 1773 830
rect 1720 762 1773 796
rect 1720 728 1731 762
rect 1765 728 1773 762
rect 1720 694 1773 728
rect 1720 660 1731 694
rect 1765 660 1773 694
rect 1720 648 1773 660
rect 1847 830 1900 848
rect 1847 796 1855 830
rect 1889 796 1900 830
rect 1847 762 1900 796
rect 1847 728 1855 762
rect 1889 728 1900 762
rect 1847 694 1900 728
rect 1847 660 1855 694
rect 1889 660 1900 694
rect 1847 648 1900 660
rect 2080 830 2133 848
rect 2080 796 2091 830
rect 2125 796 2133 830
rect 2080 762 2133 796
rect 2080 728 2091 762
rect 2125 728 2133 762
rect 2080 694 2133 728
rect 2080 660 2091 694
rect 2125 660 2133 694
rect 2080 648 2133 660
rect 1251 570 1304 588
rect 1251 536 1259 570
rect 1293 536 1304 570
rect 1251 502 1304 536
rect 1251 468 1259 502
rect 1293 468 1304 502
rect 1251 434 1304 468
rect 1251 400 1259 434
rect 1293 400 1304 434
rect 1251 388 1304 400
rect 1484 570 1540 588
rect 1484 536 1495 570
rect 1529 536 1540 570
rect 1484 502 1540 536
rect 1484 468 1495 502
rect 1529 468 1540 502
rect 1484 434 1540 468
rect 1484 400 1495 434
rect 1529 400 1540 434
rect 1484 388 1540 400
rect 1720 570 1773 588
rect 1720 536 1731 570
rect 1765 536 1773 570
rect 1720 502 1773 536
rect 1720 468 1731 502
rect 1765 468 1773 502
rect 1720 434 1773 468
rect 1720 400 1731 434
rect 1765 400 1773 434
rect 1720 388 1773 400
rect 1847 570 1900 588
rect 1847 536 1855 570
rect 1889 536 1900 570
rect 1847 502 1900 536
rect 1847 468 1855 502
rect 1889 468 1900 502
rect 1847 434 1900 468
rect 1847 400 1855 434
rect 1889 400 1900 434
rect 1847 388 1900 400
rect 2080 570 2133 588
rect 2080 536 2091 570
rect 2125 536 2133 570
rect 2080 502 2133 536
rect 2080 468 2091 502
rect 2125 468 2133 502
rect 2080 434 2133 468
rect 2080 400 2091 434
rect 2125 400 2133 434
rect 2080 388 2133 400
rect 1251 310 1304 328
rect 1251 276 1259 310
rect 1293 276 1304 310
rect 1251 242 1304 276
rect 1251 208 1259 242
rect 1293 208 1304 242
rect 1251 174 1304 208
rect 1251 140 1259 174
rect 1293 140 1304 174
rect 1251 128 1304 140
rect 1484 310 1540 328
rect 1484 276 1495 310
rect 1529 276 1540 310
rect 1484 242 1540 276
rect 1484 208 1495 242
rect 1529 208 1540 242
rect 1484 174 1540 208
rect 1484 140 1495 174
rect 1529 140 1540 174
rect 1484 128 1540 140
rect 1720 310 1773 328
rect 1720 276 1731 310
rect 1765 276 1773 310
rect 1720 242 1773 276
rect 1720 208 1731 242
rect 1765 208 1773 242
rect 1720 174 1773 208
rect 1720 140 1731 174
rect 1765 140 1773 174
rect 1720 128 1773 140
rect 1847 310 1900 328
rect 1847 276 1855 310
rect 1889 276 1900 310
rect 1847 242 1900 276
rect 1847 208 1855 242
rect 1889 208 1900 242
rect 1847 174 1900 208
rect 1847 140 1855 174
rect 1889 140 1900 174
rect 1847 128 1900 140
rect 2080 310 2133 328
rect 2080 276 2091 310
rect 2125 276 2133 310
rect 2080 242 2133 276
rect 2080 208 2091 242
rect 2125 208 2133 242
rect 2080 174 2133 208
rect 2080 140 2091 174
rect 2125 140 2133 174
rect 2080 128 2133 140
<< mvpdiff >>
rect -25 847 28 859
rect -25 813 -17 847
rect 17 813 28 847
rect -25 779 28 813
rect -25 745 -17 779
rect 17 745 28 779
rect -25 711 28 745
rect -25 677 -17 711
rect 17 677 28 711
rect -25 659 28 677
rect 128 847 181 859
rect 128 813 139 847
rect 173 813 181 847
rect 128 779 181 813
rect 128 745 139 779
rect 173 745 181 779
rect 128 711 181 745
rect 128 677 139 711
rect 173 677 181 711
rect 128 659 181 677
rect 261 720 314 732
rect 261 686 269 720
rect 303 686 314 720
rect 261 652 314 686
rect 261 618 269 652
rect 303 618 314 652
rect 261 584 314 618
rect 261 550 269 584
rect 303 550 314 584
rect 261 516 314 550
rect 261 482 269 516
rect 303 482 314 516
rect 261 448 314 482
rect -25 420 28 432
rect -25 386 -17 420
rect 17 386 28 420
rect -25 352 28 386
rect -25 318 -17 352
rect 17 318 28 352
rect -25 284 28 318
rect -25 250 -17 284
rect 17 250 28 284
rect -25 232 28 250
rect 128 420 181 432
rect 128 386 139 420
rect 173 386 181 420
rect 128 352 181 386
rect 128 318 139 352
rect 173 318 181 352
rect 128 284 181 318
rect 128 250 139 284
rect 173 250 181 284
rect 128 232 181 250
rect 261 414 269 448
rect 303 414 314 448
rect 261 380 314 414
rect 261 346 269 380
rect 303 346 314 380
rect 261 312 314 346
rect 261 278 269 312
rect 303 278 314 312
rect 261 244 314 278
rect 261 210 269 244
rect 303 210 314 244
rect 261 132 314 210
rect 414 720 470 732
rect 414 686 425 720
rect 459 686 470 720
rect 414 652 470 686
rect 414 618 425 652
rect 459 618 470 652
rect 414 584 470 618
rect 414 550 425 584
rect 459 550 470 584
rect 414 516 470 550
rect 414 482 425 516
rect 459 482 470 516
rect 414 448 470 482
rect 414 414 425 448
rect 459 414 470 448
rect 414 380 470 414
rect 414 346 425 380
rect 459 346 470 380
rect 414 312 470 346
rect 414 278 425 312
rect 459 278 470 312
rect 414 244 470 278
rect 414 210 425 244
rect 459 210 470 244
rect 414 132 470 210
rect 570 720 623 732
rect 570 686 581 720
rect 615 686 623 720
rect 570 652 623 686
rect 570 618 581 652
rect 615 618 623 652
rect 570 584 623 618
rect 570 550 581 584
rect 615 550 623 584
rect 570 516 623 550
rect 570 482 581 516
rect 615 482 623 516
rect 570 448 623 482
rect 570 414 581 448
rect 615 414 623 448
rect 570 380 623 414
rect 570 346 581 380
rect 615 346 623 380
rect 570 312 623 346
rect 570 278 581 312
rect 615 278 623 312
rect 570 244 623 278
rect 570 210 581 244
rect 615 210 623 244
rect 570 132 623 210
<< ndiffc >>
rect 2215 2150 2249 2184
rect 2215 2082 2249 2116
rect 2215 2014 2249 2048
rect 2301 2150 2335 2184
rect 2301 2082 2335 2116
rect 2301 2014 2335 2048
rect 2387 2150 2421 2184
rect 2387 2082 2421 2116
rect 2387 2014 2421 2048
rect 2215 1890 2249 1924
rect 2215 1822 2249 1856
rect 2215 1754 2249 1788
rect 2301 1890 2335 1924
rect 2301 1822 2335 1856
rect 2301 1754 2335 1788
rect 2387 1890 2421 1924
rect 2387 1822 2421 1856
rect 2387 1754 2421 1788
rect 2215 1630 2249 1664
rect 2215 1562 2249 1596
rect 2215 1494 2249 1528
rect 2301 1630 2335 1664
rect 2301 1562 2335 1596
rect 2301 1494 2335 1528
rect 2387 1630 2421 1664
rect 2387 1562 2421 1596
rect 2387 1494 2421 1528
rect 2215 1370 2249 1404
rect 2215 1302 2249 1336
rect 2215 1234 2249 1268
rect 2301 1370 2335 1404
rect 2301 1302 2335 1336
rect 2301 1234 2335 1268
rect 2387 1370 2421 1404
rect 2387 1302 2421 1336
rect 2387 1234 2421 1268
rect 2215 1056 2249 1090
rect 2215 988 2249 1022
rect 2215 920 2249 954
rect 2301 1056 2335 1090
rect 2301 988 2335 1022
rect 2301 920 2335 954
rect 2387 1056 2421 1090
rect 2387 988 2421 1022
rect 2387 920 2421 954
rect 2215 796 2249 830
rect 2215 728 2249 762
rect 2215 660 2249 694
rect 2301 796 2335 830
rect 2301 728 2335 762
rect 2301 660 2335 694
rect 2387 796 2421 830
rect 2387 728 2421 762
rect 2387 660 2421 694
rect 2634 972 2668 1006
rect 2634 904 2668 938
rect 2634 836 2668 870
rect 2740 972 2774 1006
rect 2740 904 2774 938
rect 2740 836 2774 870
rect 2846 972 2880 1006
rect 2846 904 2880 938
rect 2846 836 2880 870
rect 2952 972 2986 1006
rect 2952 904 2986 938
rect 2952 836 2986 870
rect 3058 972 3092 1006
rect 3058 904 3092 938
rect 3058 836 3092 870
rect 2215 536 2249 570
rect 2215 468 2249 502
rect 2215 400 2249 434
rect 2301 536 2335 570
rect 2301 468 2335 502
rect 2301 400 2335 434
rect 2387 536 2421 570
rect 2387 468 2421 502
rect 2387 400 2421 434
rect 2215 276 2249 310
rect 2215 208 2249 242
rect 2215 140 2249 174
rect 2301 276 2335 310
rect 2301 208 2335 242
rect 2301 140 2335 174
rect 2387 276 2421 310
rect 2387 208 2421 242
rect 2387 140 2421 174
<< pdiffc >>
rect 2779 1796 2813 1830
rect 2779 1728 2813 1762
rect 2779 1660 2813 1694
rect 2779 1592 2813 1626
rect 2779 1524 2813 1558
rect 2779 1456 2813 1490
rect 2779 1388 2813 1422
rect 2779 1320 2813 1354
rect 2885 1796 2919 1830
rect 2885 1728 2919 1762
rect 2885 1660 2919 1694
rect 2885 1592 2919 1626
rect 2885 1524 2919 1558
rect 2885 1456 2919 1490
rect 2885 1388 2919 1422
rect 2885 1320 2919 1354
rect 2991 1796 3025 1830
rect 2991 1728 3025 1762
rect 2991 1660 3025 1694
rect 2991 1592 3025 1626
rect 2991 1524 3025 1558
rect 2991 1456 3025 1490
rect 2991 1388 3025 1422
rect 2991 1320 3025 1354
<< mvndiffc >>
rect 1266 2156 1300 2190
rect 1266 2088 1300 2122
rect 781 1978 815 2012
rect 781 1910 815 1944
rect 781 1842 815 1876
rect 781 1774 815 1808
rect 781 1706 815 1740
rect 781 1638 815 1672
rect 781 1570 815 1604
rect 781 1502 815 1536
rect 957 1978 991 2012
rect 957 1910 991 1944
rect 957 1842 991 1876
rect 957 1774 991 1808
rect 957 1706 991 1740
rect 957 1638 991 1672
rect 957 1570 991 1604
rect 957 1502 991 1536
rect 1133 1978 1167 2012
rect 1133 1910 1167 1944
rect 1133 1842 1167 1876
rect 1133 1774 1167 1808
rect 1133 1706 1167 1740
rect 1133 1638 1167 1672
rect 1133 1570 1167 1604
rect 1133 1502 1167 1536
rect 1266 2020 1300 2054
rect 1266 1952 1300 1986
rect 1266 1884 1300 1918
rect 1266 1816 1300 1850
rect 1266 1748 1300 1782
rect 1266 1680 1300 1714
rect 1266 1612 1300 1646
rect 1266 1544 1300 1578
rect 1266 1476 1300 1510
rect 1266 1408 1300 1442
rect 1266 1340 1300 1374
rect 41 1236 75 1270
rect 41 1168 75 1202
rect 41 1100 75 1134
rect 217 1236 251 1270
rect 217 1168 251 1202
rect 217 1100 251 1134
rect 393 1236 427 1270
rect 1266 1272 1300 1306
rect 393 1168 427 1202
rect 393 1100 427 1134
rect 781 1176 815 1210
rect 781 1108 815 1142
rect 957 1176 991 1210
rect 957 1108 991 1142
rect 1133 1176 1167 1210
rect 1422 2156 1456 2190
rect 1422 2088 1456 2122
rect 1422 2020 1456 2054
rect 1422 1952 1456 1986
rect 1422 1884 1456 1918
rect 1422 1816 1456 1850
rect 1422 1748 1456 1782
rect 1422 1680 1456 1714
rect 1422 1612 1456 1646
rect 1422 1544 1456 1578
rect 1422 1476 1456 1510
rect 1422 1408 1456 1442
rect 1422 1340 1456 1374
rect 1422 1272 1456 1306
rect 1575 2156 1609 2190
rect 1575 2088 1609 2122
rect 1575 2020 1609 2054
rect 1575 1952 1609 1986
rect 1575 1884 1609 1918
rect 1575 1816 1609 1850
rect 1575 1748 1609 1782
rect 1575 1680 1609 1714
rect 1575 1612 1609 1646
rect 1575 1544 1609 1578
rect 1575 1476 1609 1510
rect 1575 1408 1609 1442
rect 1575 1340 1609 1374
rect 1575 1272 1609 1306
rect 1731 2156 1765 2190
rect 1731 2088 1765 2122
rect 1731 2020 1765 2054
rect 1855 2150 1889 2184
rect 1855 2082 1889 2116
rect 1855 2014 1889 2048
rect 2091 2150 2125 2184
rect 2091 2082 2125 2116
rect 2091 2014 2125 2048
rect 1731 1952 1765 1986
rect 1731 1884 1765 1918
rect 1731 1816 1765 1850
rect 1731 1748 1765 1782
rect 1855 1890 1889 1924
rect 1855 1822 1889 1856
rect 1855 1754 1889 1788
rect 2091 1890 2125 1924
rect 2091 1822 2125 1856
rect 2091 1754 2125 1788
rect 1731 1680 1765 1714
rect 1731 1612 1765 1646
rect 1731 1544 1765 1578
rect 1731 1476 1765 1510
rect 1855 1630 1889 1664
rect 1855 1562 1889 1596
rect 1855 1494 1889 1528
rect 2091 1630 2125 1664
rect 2091 1562 2125 1596
rect 2091 1494 2125 1528
rect 1731 1408 1765 1442
rect 1731 1340 1765 1374
rect 1731 1272 1765 1306
rect 1855 1370 1889 1404
rect 1855 1302 1889 1336
rect 1855 1234 1889 1268
rect 2091 1370 2125 1404
rect 2091 1302 2125 1336
rect 2091 1234 2125 1268
rect 1133 1108 1167 1142
rect 1259 1056 1293 1090
rect 1259 988 1293 1022
rect 1259 920 1293 954
rect 1495 1056 1529 1090
rect 1495 988 1529 1022
rect 1495 920 1529 954
rect 1731 1056 1765 1090
rect 1731 988 1765 1022
rect 1731 920 1765 954
rect 1855 1056 1889 1090
rect 1855 988 1889 1022
rect 1855 920 1889 954
rect 2091 1056 2125 1090
rect 2091 988 2125 1022
rect 2091 920 2125 954
rect 1259 796 1293 830
rect 1259 728 1293 762
rect 1259 660 1293 694
rect 1495 796 1529 830
rect 1495 728 1529 762
rect 1495 660 1529 694
rect 1731 796 1765 830
rect 1731 728 1765 762
rect 1731 660 1765 694
rect 1855 796 1889 830
rect 1855 728 1889 762
rect 1855 660 1889 694
rect 2091 796 2125 830
rect 2091 728 2125 762
rect 2091 660 2125 694
rect 1259 536 1293 570
rect 1259 468 1293 502
rect 1259 400 1293 434
rect 1495 536 1529 570
rect 1495 468 1529 502
rect 1495 400 1529 434
rect 1731 536 1765 570
rect 1731 468 1765 502
rect 1731 400 1765 434
rect 1855 536 1889 570
rect 1855 468 1889 502
rect 1855 400 1889 434
rect 2091 536 2125 570
rect 2091 468 2125 502
rect 2091 400 2125 434
rect 1259 276 1293 310
rect 1259 208 1293 242
rect 1259 140 1293 174
rect 1495 276 1529 310
rect 1495 208 1529 242
rect 1495 140 1529 174
rect 1731 276 1765 310
rect 1731 208 1765 242
rect 1731 140 1765 174
rect 1855 276 1889 310
rect 1855 208 1889 242
rect 1855 140 1889 174
rect 2091 276 2125 310
rect 2091 208 2125 242
rect 2091 140 2125 174
<< mvpdiffc >>
rect -17 813 17 847
rect -17 745 17 779
rect -17 677 17 711
rect 139 813 173 847
rect 139 745 173 779
rect 139 677 173 711
rect 269 686 303 720
rect 269 618 303 652
rect 269 550 303 584
rect 269 482 303 516
rect -17 386 17 420
rect -17 318 17 352
rect -17 250 17 284
rect 139 386 173 420
rect 139 318 173 352
rect 139 250 173 284
rect 269 414 303 448
rect 269 346 303 380
rect 269 278 303 312
rect 269 210 303 244
rect 425 686 459 720
rect 425 618 459 652
rect 425 550 459 584
rect 425 482 459 516
rect 425 414 459 448
rect 425 346 459 380
rect 425 278 459 312
rect 425 210 459 244
rect 581 686 615 720
rect 581 618 615 652
rect 581 550 615 584
rect 581 482 615 516
rect 581 414 615 448
rect 581 346 615 380
rect 581 278 615 312
rect 581 210 615 244
<< psubdiff >>
rect 2503 2145 2537 2169
rect 2503 2076 2537 2111
rect 2503 2007 2537 2042
rect 2503 1938 2537 1973
rect 2503 1869 2537 1904
rect 2503 1800 2537 1835
rect 2503 1731 2537 1766
rect 2503 1662 2537 1697
rect 2503 1594 2537 1628
rect 2503 1526 2537 1560
rect 2503 1458 2537 1492
rect 2503 1390 2537 1424
rect 2503 1322 2537 1356
rect 2503 1254 2537 1288
rect 2503 1186 2537 1220
rect 2503 1118 2537 1152
rect 2503 1050 2537 1084
rect 2503 982 2537 1016
rect 2503 914 2537 948
rect 2503 846 2537 880
rect 2503 778 2537 812
rect 2503 710 2537 744
rect 2503 642 2537 676
rect 2503 574 2537 608
rect 2503 506 2537 540
rect 2503 438 2537 472
rect 2503 370 2537 404
rect 2503 302 2537 336
rect 2503 234 2537 268
rect 2503 166 2537 200
rect 2503 108 2537 132
<< nsubdiff >>
rect 3131 1818 3165 1842
rect 3131 1750 3165 1784
rect 3131 1682 3165 1716
rect 3131 1614 3165 1648
rect 3131 1546 3165 1580
rect 3131 1478 3165 1512
rect 3131 1410 3165 1444
rect 3131 1342 3165 1376
rect 3131 1244 3165 1308
<< mvpsubdiff >>
rect 943 830 1161 854
rect 943 116 967 830
rect 1137 116 1161 830
rect 943 92 1161 116
<< mvnsubdiff >>
rect 717 708 751 732
rect 717 634 751 674
rect 717 560 751 600
rect 717 486 751 526
rect 717 412 751 452
rect 717 338 751 378
rect 717 264 751 304
rect 717 190 751 230
rect 717 132 751 156
<< psubdiffcont >>
rect 2503 2111 2537 2145
rect 2503 2042 2537 2076
rect 2503 1973 2537 2007
rect 2503 1904 2537 1938
rect 2503 1835 2537 1869
rect 2503 1766 2537 1800
rect 2503 1697 2537 1731
rect 2503 1628 2537 1662
rect 2503 1560 2537 1594
rect 2503 1492 2537 1526
rect 2503 1424 2537 1458
rect 2503 1356 2537 1390
rect 2503 1288 2537 1322
rect 2503 1220 2537 1254
rect 2503 1152 2537 1186
rect 2503 1084 2537 1118
rect 2503 1016 2537 1050
rect 2503 948 2537 982
rect 2503 880 2537 914
rect 2503 812 2537 846
rect 2503 744 2537 778
rect 2503 676 2537 710
rect 2503 608 2537 642
rect 2503 540 2537 574
rect 2503 472 2537 506
rect 2503 404 2537 438
rect 2503 336 2537 370
rect 2503 268 2537 302
rect 2503 200 2537 234
rect 2503 132 2537 166
<< nsubdiffcont >>
rect 3131 1784 3165 1818
rect 3131 1716 3165 1750
rect 3131 1648 3165 1682
rect 3131 1580 3165 1614
rect 3131 1512 3165 1546
rect 3131 1444 3165 1478
rect 3131 1376 3165 1410
rect 3131 1308 3165 1342
<< mvpsubdiffcont >>
rect 967 116 1137 830
<< mvnsubdiffcont >>
rect 717 674 751 708
rect 717 600 751 634
rect 717 526 751 560
rect 717 452 751 486
rect 717 378 751 412
rect 717 304 751 338
rect 717 230 751 264
rect 717 156 751 190
<< poly >>
rect 1311 2278 1720 2294
rect 1311 2244 1329 2278
rect 1363 2244 1397 2278
rect 1431 2244 1465 2278
rect 1499 2244 1533 2278
rect 1567 2244 1601 2278
rect 1635 2244 1669 2278
rect 1703 2244 1720 2278
rect 1311 2228 1720 2244
rect 1311 2202 1411 2228
rect 1620 2202 1720 2228
rect 1900 2278 2080 2294
rect 1900 2244 1939 2278
rect 1973 2244 2007 2278
rect 2041 2244 2080 2278
rect 1900 2202 2080 2244
rect 2251 2278 2385 2294
rect 2251 2244 2267 2278
rect 2301 2244 2335 2278
rect 2369 2244 2385 2278
rect 2251 2228 2385 2244
rect 2260 2202 2290 2228
rect 2346 2202 2376 2228
rect 812 2106 946 2122
rect 812 2072 828 2106
rect 862 2072 896 2106
rect 930 2072 946 2106
rect 812 2050 946 2072
rect 826 2024 946 2050
rect 1002 2106 1136 2122
rect 1002 2072 1018 2106
rect 1052 2072 1086 2106
rect 1120 2072 1136 2106
rect 1002 2050 1136 2072
rect 1002 2024 1122 2050
rect 826 1398 946 1424
rect 1002 1398 1122 1424
rect 86 1282 206 1308
rect 262 1282 382 1308
rect 826 1222 946 1248
rect 1002 1222 1122 1248
rect 1900 1942 2080 2002
rect 2260 1942 2290 2002
rect 2346 1942 2376 2002
rect 2824 1842 2874 1874
rect 2930 1842 2980 1874
rect 1900 1682 2080 1742
rect 2260 1682 2290 1742
rect 2346 1682 2376 1742
rect 1900 1422 2080 1482
rect 2260 1422 2290 1482
rect 2346 1422 2376 1482
rect 1311 1176 1411 1202
rect 1620 1176 1720 1202
rect 1900 1182 2080 1222
rect 2260 1196 2290 1222
rect 2346 1196 2376 1222
rect 1900 1148 1939 1182
rect 1973 1148 2007 1182
rect 2041 1148 2080 1182
rect 1304 1108 1484 1134
rect 1540 1108 1720 1134
rect 1900 1108 2080 1148
rect 2824 1210 2874 1242
rect 2260 1108 2290 1134
rect 2346 1108 2376 1134
rect 2740 1194 2874 1210
rect 2740 1160 2756 1194
rect 2790 1160 2824 1194
rect 2858 1160 2874 1194
rect 2740 1144 2874 1160
rect 2930 1210 2980 1242
rect 2930 1194 3064 1210
rect 2930 1160 2946 1194
rect 2980 1160 3014 1194
rect 3048 1160 3064 1194
rect 2930 1144 3064 1160
rect 2740 1119 2835 1144
rect 2930 1119 3049 1144
rect 86 1056 206 1082
rect 28 1030 206 1056
rect 28 928 67 1030
rect 169 928 206 1030
rect 28 885 206 928
rect 262 1056 382 1082
rect 262 1010 414 1056
rect 262 908 278 1010
rect 380 908 414 1010
rect 826 1040 946 1082
rect 826 1006 869 1040
rect 903 1006 946 1040
rect 826 972 946 1006
rect 826 938 869 972
rect 903 938 946 972
rect 826 922 946 938
rect 1002 1040 1122 1082
rect 1002 1006 1018 1040
rect 1052 1006 1122 1040
rect 1002 972 1122 1006
rect 1002 938 1018 972
rect 1052 938 1122 972
rect 1002 922 1122 938
rect 2679 1103 2835 1119
rect 2908 1104 3049 1119
rect 2679 1069 2695 1103
rect 2729 1069 2785 1103
rect 2819 1069 2835 1103
rect 2679 1053 2835 1069
rect 2679 1024 2729 1053
rect 2785 1024 2835 1053
rect 2891 1103 3049 1104
rect 2891 1069 2924 1103
rect 2958 1069 2999 1103
rect 3033 1069 3049 1103
rect 2891 1053 3049 1069
rect 2891 1024 2941 1053
rect 2997 1024 3047 1053
rect 28 859 128 885
rect 262 758 414 908
rect 1304 848 1484 908
rect 1540 848 1720 908
rect 1900 848 2080 908
rect 2260 848 2290 908
rect 2346 848 2376 908
rect 314 732 414 758
rect 470 732 570 758
rect 28 633 128 659
rect 28 432 128 458
rect 28 106 128 232
rect 314 106 414 132
rect 28 14 414 106
rect 470 106 570 132
rect 2679 798 2729 824
rect 2785 798 2835 824
rect 2891 798 2941 824
rect 2997 798 3047 824
rect 1304 588 1484 648
rect 1540 588 1720 648
rect 1900 588 2080 648
rect 2260 588 2290 648
rect 2346 588 2376 648
rect 1304 328 1484 388
rect 1540 328 1720 388
rect 1900 328 2080 388
rect 2260 328 2290 388
rect 2346 328 2376 388
rect 470 80 603 106
rect 1304 102 1484 128
rect 1540 102 1720 128
rect 1900 102 2080 128
rect 2260 102 2290 128
rect 2346 102 2376 128
rect 1304 86 2080 102
rect 470 64 604 80
rect 470 30 486 64
rect 520 30 554 64
rect 588 30 604 64
rect 1304 52 1328 86
rect 1362 52 1396 86
rect 1430 52 1464 86
rect 1498 52 1532 86
rect 1566 52 1600 86
rect 1634 52 1668 86
rect 1702 52 1736 86
rect 1770 52 1804 86
rect 1838 52 1872 86
rect 1906 52 1940 86
rect 1974 52 2008 86
rect 2042 52 2080 86
rect 1304 36 2080 52
rect 2251 86 2385 102
rect 2251 52 2267 86
rect 2301 52 2335 86
rect 2369 52 2385 86
rect 2251 36 2385 52
rect 470 14 604 30
<< polycont >>
rect 1329 2244 1363 2278
rect 1397 2244 1431 2278
rect 1465 2244 1499 2278
rect 1533 2244 1567 2278
rect 1601 2244 1635 2278
rect 1669 2244 1703 2278
rect 1939 2244 1973 2278
rect 2007 2244 2041 2278
rect 2267 2244 2301 2278
rect 2335 2244 2369 2278
rect 828 2072 862 2106
rect 896 2072 930 2106
rect 1018 2072 1052 2106
rect 1086 2072 1120 2106
rect 1939 1148 1973 1182
rect 2007 1148 2041 1182
rect 2756 1160 2790 1194
rect 2824 1160 2858 1194
rect 2946 1160 2980 1194
rect 3014 1160 3048 1194
rect 67 928 169 1030
rect 278 908 380 1010
rect 869 1006 903 1040
rect 869 938 903 972
rect 1018 1006 1052 1040
rect 1018 938 1052 972
rect 2695 1069 2729 1103
rect 2785 1069 2819 1103
rect 2924 1069 2958 1103
rect 2999 1069 3033 1103
rect 486 30 520 64
rect 554 30 588 64
rect 1328 52 1362 86
rect 1396 52 1430 86
rect 1464 52 1498 86
rect 1532 52 1566 86
rect 1600 52 1634 86
rect 1668 52 1702 86
rect 1736 52 1770 86
rect 1804 52 1838 86
rect 1872 52 1906 86
rect 1940 52 1974 86
rect 2008 52 2042 86
rect 2267 52 2301 86
rect 2335 52 2369 86
<< locali >>
rect 812 2106 946 2379
rect 812 2072 828 2106
rect 862 2072 896 2106
rect 930 2072 946 2106
rect 1002 2106 1136 2392
rect 2251 2354 2279 2388
rect 2313 2354 2351 2388
rect 2251 2278 2385 2354
rect 1313 2244 1329 2278
rect 1363 2244 1397 2278
rect 1431 2244 1465 2278
rect 1499 2244 1533 2278
rect 1567 2244 1601 2278
rect 1635 2244 1669 2278
rect 1703 2244 1719 2278
rect 1923 2244 1939 2278
rect 1973 2244 2007 2278
rect 2041 2244 2057 2278
rect 2251 2244 2267 2278
rect 2301 2244 2335 2278
rect 2369 2244 2385 2278
rect 1002 2072 1018 2106
rect 1052 2072 1086 2106
rect 1120 2072 1136 2106
rect 1266 2190 1300 2206
rect 1266 2122 1300 2156
rect 1266 2054 1300 2088
rect 781 2012 815 2028
rect 781 1944 815 1978
rect 781 1876 815 1910
rect 781 1808 815 1842
rect 781 1740 815 1771
rect 781 1672 815 1699
rect 781 1604 815 1638
rect 781 1536 815 1570
rect 217 1387 641 1443
rect 41 1270 75 1286
rect 41 1202 75 1236
rect 41 1134 75 1168
rect 41 1098 75 1100
rect 323 1382 641 1387
rect 323 1348 393 1382
rect 427 1348 465 1382
rect 323 1320 494 1348
rect 217 1270 323 1281
rect 251 1236 323 1270
rect 217 1202 323 1236
rect 251 1168 323 1202
rect 217 1134 323 1168
rect 251 1100 323 1134
rect 75 1064 113 1098
rect 217 1080 323 1100
rect 393 1270 448 1286
rect 427 1236 448 1270
rect 482 1276 494 1320
rect 571 1310 641 1382
rect 600 1276 641 1310
rect 482 1265 641 1276
rect 393 1202 448 1236
rect 427 1168 448 1202
rect 393 1134 448 1168
rect 427 1100 448 1134
rect 393 1084 448 1100
rect 781 1210 815 1502
rect 781 1142 815 1176
rect 51 928 67 1030
rect 169 1018 185 1030
rect 278 1010 380 1026
rect 169 928 185 984
rect -17 847 17 863
rect -17 779 17 813
rect -17 711 17 745
rect -17 420 17 677
rect -17 352 17 386
rect -17 294 17 318
rect -17 222 17 250
rect -17 150 17 188
rect 51 436 105 928
rect 274 908 278 910
rect 274 894 380 908
rect 139 857 380 894
rect 139 847 173 857
rect 414 823 448 1084
rect 139 779 173 813
rect 139 711 173 745
rect 139 661 173 677
rect 269 789 448 823
rect 516 1058 554 1092
rect 482 796 588 1058
rect 781 944 815 1108
rect 957 2012 991 2028
rect 957 1944 991 1978
rect 957 1876 991 1910
rect 957 1808 991 1842
rect 957 1740 991 1774
rect 957 1672 991 1706
rect 957 1604 991 1638
rect 957 1536 991 1570
rect 957 1443 991 1502
rect 957 1371 991 1409
rect 957 1299 991 1337
rect 957 1210 991 1265
rect 957 1142 991 1176
rect 957 1092 991 1108
rect 1133 2020 1266 2028
rect 1133 2012 1300 2020
rect 1167 1986 1300 2012
rect 1167 1978 1266 1986
rect 1133 1952 1266 1978
rect 1133 1944 1300 1952
rect 1167 1918 1300 1944
rect 1167 1910 1266 1918
rect 1133 1884 1266 1910
rect 1133 1876 1300 1884
rect 1167 1850 1300 1876
rect 1167 1842 1266 1850
rect 1133 1816 1266 1842
rect 1133 1808 1300 1816
rect 1167 1782 1300 1808
rect 1167 1774 1266 1782
rect 1133 1748 1266 1774
rect 1133 1740 1300 1748
rect 1167 1714 1300 1740
rect 1167 1706 1266 1714
rect 1133 1680 1266 1706
rect 1133 1672 1300 1680
rect 1167 1646 1300 1672
rect 1167 1638 1266 1646
rect 1133 1612 1266 1638
rect 1133 1604 1300 1612
rect 1167 1578 1300 1604
rect 1167 1570 1266 1578
rect 1133 1544 1266 1570
rect 1133 1536 1300 1544
rect 1167 1510 1300 1536
rect 1167 1502 1266 1510
rect 1133 1476 1266 1502
rect 1133 1442 1300 1476
rect 1133 1408 1266 1442
rect 1133 1374 1300 1408
rect 1133 1340 1266 1374
rect 1133 1306 1300 1340
rect 1133 1272 1266 1306
rect 1133 1256 1300 1272
rect 1422 2190 1456 2206
rect 1422 2122 1456 2156
rect 1422 2054 1456 2088
rect 1422 1986 1456 2020
rect 1422 1918 1456 1952
rect 1422 1850 1456 1884
rect 1422 1782 1456 1816
rect 1575 2190 1609 2206
rect 1575 2122 1609 2156
rect 1575 2054 1609 2088
rect 1575 1986 1609 2020
rect 1575 1918 1609 1952
rect 1575 1850 1609 1884
rect 1575 1811 1609 1816
rect 1731 2190 1889 2206
rect 1765 2184 1889 2190
rect 1765 2156 1855 2184
rect 1731 2150 1855 2156
rect 1731 2122 1889 2150
rect 1765 2116 1889 2122
rect 1765 2088 1855 2116
rect 1731 2082 1855 2088
rect 1731 2054 1889 2082
rect 1765 2048 1889 2054
rect 1765 2020 1855 2048
rect 1731 2014 1855 2020
rect 1731 1986 1889 2014
rect 1765 1952 1889 1986
rect 1731 1924 1889 1952
rect 1731 1918 1855 1924
rect 1765 1890 1855 1918
rect 1765 1884 1889 1890
rect 1731 1856 1889 1884
rect 1731 1850 1855 1856
rect 1765 1822 1855 1850
rect 1765 1816 1889 1822
rect 1553 1782 1591 1811
rect 1553 1777 1575 1782
rect 1731 1788 1889 1816
rect 1731 1782 1855 1788
rect 1422 1714 1456 1748
rect 1422 1646 1456 1680
rect 1422 1578 1456 1612
rect 1422 1510 1456 1544
rect 1422 1442 1456 1476
rect 1422 1374 1456 1408
rect 1422 1306 1456 1340
rect 1133 1210 1167 1256
rect 1422 1180 1456 1272
rect 1575 1714 1609 1748
rect 1575 1646 1609 1680
rect 1575 1578 1609 1612
rect 1575 1510 1609 1544
rect 1575 1442 1609 1476
rect 1575 1374 1609 1408
rect 1575 1306 1609 1340
rect 1575 1256 1609 1272
rect 1765 1754 1855 1782
rect 1765 1748 1889 1754
rect 1731 1714 1889 1748
rect 1765 1680 1889 1714
rect 1731 1664 1889 1680
rect 1731 1646 1855 1664
rect 1765 1630 1855 1646
rect 1765 1612 1889 1630
rect 1731 1596 1889 1612
rect 1731 1578 1855 1596
rect 1765 1562 1855 1578
rect 1765 1544 1889 1562
rect 1731 1528 1889 1544
rect 1731 1510 1855 1528
rect 1765 1494 1855 1510
rect 1765 1476 1889 1494
rect 1731 1442 1889 1476
rect 1765 1408 1889 1442
rect 1731 1404 1889 1408
rect 1731 1374 1855 1404
rect 1765 1370 1855 1374
rect 1765 1340 1889 1370
rect 1731 1336 1889 1340
rect 1731 1306 1855 1336
rect 1765 1302 1855 1306
rect 1765 1272 1889 1302
rect 1731 1268 1889 1272
rect 1731 1256 1855 1268
rect 1133 1142 1167 1176
rect 743 910 781 944
rect 853 1018 869 1040
rect 903 1018 919 1040
rect 903 1006 925 1018
rect 887 984 925 1006
rect 1002 1006 1018 1040
rect 1052 1006 1068 1040
rect 1133 1018 1167 1108
rect 1259 1140 1765 1180
rect 1259 1090 1293 1140
rect 1259 1022 1293 1056
rect 853 972 919 984
rect 853 938 869 972
rect 903 938 919 972
rect 1002 972 1068 1006
rect 1137 984 1175 1018
rect 1002 944 1018 972
rect 1052 944 1068 972
rect 1259 954 1293 988
rect 1052 938 1074 944
rect 1036 910 1074 938
rect 967 830 1137 846
rect 269 720 303 789
rect 482 762 615 796
rect 269 652 303 686
rect 269 584 303 618
rect 269 516 303 550
rect 269 448 303 482
rect 51 420 173 436
rect 51 386 139 420
rect 51 352 173 386
rect 51 318 139 352
rect 51 284 173 318
rect 51 250 139 284
rect 51 64 173 250
rect 269 380 303 414
rect 269 312 303 346
rect 269 244 303 278
rect 269 194 303 210
rect 425 720 459 736
rect 425 652 459 686
rect 425 584 459 618
rect 425 516 459 550
rect 425 448 459 482
rect 425 380 459 414
rect 425 312 459 346
rect 425 244 459 260
rect 581 720 615 762
rect 581 652 615 686
rect 581 584 615 618
rect 581 516 615 550
rect 581 448 615 482
rect 581 380 615 414
rect 581 312 615 346
rect 581 244 615 278
rect 581 194 615 210
rect 717 708 751 732
rect 717 634 751 674
rect 717 560 751 600
rect 717 486 751 526
rect 717 412 751 452
rect 717 338 751 378
rect 717 294 751 304
rect 717 222 751 230
rect 425 150 459 188
rect 717 150 751 156
rect 1259 830 1293 920
rect 1259 762 1293 796
rect 1259 694 1293 728
rect 1259 570 1293 660
rect 1259 502 1293 536
rect 1259 434 1293 468
rect 1259 310 1293 400
rect 1259 242 1293 276
rect 1259 174 1293 208
rect 1259 124 1293 140
rect 1495 1090 1529 1106
rect 1495 1022 1529 1056
rect 1495 954 1529 988
rect 1495 830 1529 916
rect 1495 762 1529 796
rect 1495 694 1529 728
rect 1495 570 1529 660
rect 1495 502 1529 536
rect 1495 434 1529 468
rect 1495 310 1529 400
rect 1495 242 1529 276
rect 1495 174 1529 208
rect 1495 124 1529 140
rect 1731 1090 1765 1140
rect 1731 1022 1765 1056
rect 1731 954 1765 988
rect 1731 830 1765 920
rect 1731 762 1765 796
rect 1731 694 1765 728
rect 1731 570 1765 660
rect 1731 502 1765 536
rect 1731 434 1765 468
rect 1731 310 1765 400
rect 1731 242 1765 276
rect 1731 174 1765 208
rect 1731 124 1765 140
rect 1855 1090 1889 1234
rect 1855 1022 1889 1056
rect 1855 954 1889 988
rect 1855 830 1889 920
rect 1855 762 1889 796
rect 1855 694 1889 728
rect 1855 570 1889 660
rect 1855 502 1889 536
rect 1855 434 1889 468
rect 1855 310 1889 400
rect 1855 242 1889 276
rect 1855 174 1889 208
rect 1855 124 1889 140
rect 1923 2090 2057 2244
rect 1923 1912 1937 2090
rect 2043 1912 2057 2090
rect 1923 1182 2057 1912
rect 1923 1148 1939 1182
rect 1973 1148 2007 1182
rect 2041 1148 2057 1182
rect 967 100 1137 116
rect 1923 90 2057 1148
rect 2091 2184 2125 2200
rect 2091 2116 2125 2150
rect 2091 2048 2125 2082
rect 2091 1924 2125 2014
rect 2091 1856 2125 1890
rect 2091 1788 2125 1822
rect 2091 1664 2125 1754
rect 2091 1596 2125 1630
rect 2091 1528 2125 1561
rect 2091 1404 2125 1489
rect 2091 1336 2125 1370
rect 2091 1268 2125 1302
rect 2091 1090 2125 1234
rect 2091 1022 2125 1056
rect 2091 954 2125 988
rect 2091 830 2125 920
rect 2091 762 2125 796
rect 2091 694 2125 728
rect 2091 570 2125 660
rect 2091 502 2125 536
rect 2091 434 2125 468
rect 2091 310 2125 400
rect 2091 242 2125 276
rect 2091 174 2125 208
rect 2091 124 2125 140
rect 2159 2184 2267 2200
rect 2159 2150 2215 2184
rect 2249 2150 2267 2184
rect 2159 2116 2267 2150
rect 2159 2082 2215 2116
rect 2249 2082 2267 2116
rect 2159 2048 2267 2082
rect 2159 2014 2215 2048
rect 2249 2014 2267 2048
rect 2159 1924 2267 2014
rect 2159 1890 2215 1924
rect 2249 1890 2267 1924
rect 2159 1856 2267 1890
rect 2159 1822 2215 1856
rect 2249 1822 2267 1856
rect 2159 1788 2267 1822
rect 2159 1754 2215 1788
rect 2249 1754 2267 1788
rect 2159 1664 2267 1754
rect 2159 1630 2215 1664
rect 2249 1630 2267 1664
rect 2159 1596 2267 1630
rect 2159 1562 2215 1596
rect 2249 1562 2267 1596
rect 2159 1528 2267 1562
rect 2159 1494 2215 1528
rect 2249 1494 2267 1528
rect 2159 1443 2267 1494
rect 2159 1409 2202 1443
rect 2236 1409 2267 1443
rect 2159 1404 2267 1409
rect 2159 1371 2215 1404
rect 2159 1337 2202 1371
rect 2249 1370 2267 1404
rect 2236 1337 2267 1370
rect 2159 1336 2267 1337
rect 2159 1302 2215 1336
rect 2249 1302 2267 1336
rect 2159 1299 2267 1302
rect 2159 1265 2202 1299
rect 2236 1268 2267 1299
rect 2159 1234 2215 1265
rect 2249 1234 2267 1268
rect 2159 1090 2267 1234
rect 2301 2184 2335 2200
rect 2301 2116 2335 2150
rect 2301 2048 2335 2082
rect 2301 1924 2335 2014
rect 2301 1856 2335 1890
rect 2301 1788 2335 1822
rect 2301 1664 2335 1754
rect 2301 1596 2335 1630
rect 2301 1528 2335 1561
rect 2301 1404 2335 1489
rect 2301 1336 2335 1370
rect 2301 1268 2335 1302
rect 2301 1218 2335 1234
rect 2369 2184 2537 2200
rect 2369 2150 2387 2184
rect 2421 2150 2537 2184
rect 2369 2145 2537 2150
rect 2369 2116 2503 2145
rect 2369 2082 2387 2116
rect 2421 2111 2503 2116
rect 2421 2082 2537 2111
rect 2369 2076 2537 2082
rect 2369 2048 2503 2076
rect 2369 2014 2387 2048
rect 2421 2042 2503 2048
rect 2421 2014 2537 2042
rect 2369 2007 2537 2014
rect 2369 1973 2503 2007
rect 2369 1938 2537 1973
rect 2369 1924 2503 1938
rect 2369 1890 2387 1924
rect 2421 1904 2503 1924
rect 2421 1890 2537 1904
rect 2369 1869 2537 1890
rect 2369 1856 2503 1869
rect 2369 1822 2387 1856
rect 2421 1835 2503 1856
rect 2848 1957 2956 1986
rect 2848 1923 2849 1957
rect 2883 1923 2922 1957
rect 2848 1885 2956 1923
rect 2848 1851 2849 1885
rect 2883 1851 2922 1885
rect 2421 1822 2537 1835
rect 2369 1800 2537 1822
rect 2369 1788 2503 1800
rect 2369 1754 2387 1788
rect 2421 1766 2503 1788
rect 2421 1754 2537 1766
rect 2369 1731 2537 1754
rect 2779 1830 2813 1846
rect 2779 1762 2813 1796
rect 2369 1697 2503 1731
rect 2369 1664 2537 1697
rect 2369 1630 2387 1664
rect 2421 1662 2537 1664
rect 2421 1630 2503 1662
rect 2369 1628 2503 1630
rect 2369 1596 2537 1628
rect 2369 1562 2387 1596
rect 2421 1594 2537 1596
rect 2421 1562 2503 1594
rect 2369 1560 2503 1562
rect 2369 1528 2537 1560
rect 2369 1494 2387 1528
rect 2421 1526 2537 1528
rect 2421 1494 2503 1526
rect 2369 1492 2503 1494
rect 2369 1458 2537 1492
rect 2369 1443 2503 1458
rect 2369 1409 2387 1443
rect 2421 1409 2503 1443
rect 2369 1404 2537 1409
rect 2369 1337 2387 1404
rect 2421 1390 2537 1404
rect 2421 1337 2503 1390
rect 2369 1336 2537 1337
rect 2369 1302 2387 1336
rect 2421 1322 2537 1336
rect 2421 1302 2503 1322
rect 2369 1299 2503 1302
rect 2369 1234 2387 1299
rect 2421 1265 2503 1299
rect 2421 1254 2537 1265
rect 2421 1234 2503 1254
rect 2369 1220 2503 1234
rect 2369 1186 2537 1220
rect 2369 1152 2503 1186
rect 2369 1118 2537 1152
rect 2159 1056 2215 1090
rect 2249 1056 2267 1090
rect 2159 1022 2267 1056
rect 2159 988 2215 1022
rect 2249 988 2267 1022
rect 2159 954 2267 988
rect 2159 920 2215 954
rect 2249 920 2267 954
rect 2159 830 2267 920
rect 2159 796 2215 830
rect 2249 796 2267 830
rect 2159 762 2267 796
rect 2159 728 2215 762
rect 2249 728 2267 762
rect 2159 694 2267 728
rect 2159 660 2215 694
rect 2249 660 2267 694
rect 2159 570 2267 660
rect 2159 536 2215 570
rect 2249 536 2267 570
rect 2159 502 2267 536
rect 2159 468 2215 502
rect 2249 468 2267 502
rect 2159 452 2267 468
rect 2159 418 2203 452
rect 2237 434 2267 452
rect 2159 400 2215 418
rect 2249 400 2267 434
rect 2159 380 2267 400
rect 2159 346 2203 380
rect 2237 346 2267 380
rect 2159 310 2267 346
rect 2159 276 2215 310
rect 2249 276 2267 310
rect 2159 242 2267 276
rect 2159 208 2215 242
rect 2249 208 2267 242
rect 2159 174 2267 208
rect 2159 140 2215 174
rect 2249 140 2267 174
rect 2159 124 2267 140
rect 2301 1090 2335 1106
rect 2301 1022 2335 1056
rect 2301 954 2335 988
rect 2301 830 2335 916
rect 2301 762 2335 796
rect 2301 694 2335 728
rect 2301 570 2335 660
rect 2301 502 2335 536
rect 2301 434 2335 468
rect 2301 310 2335 400
rect 2301 242 2335 276
rect 2301 174 2335 208
rect 2301 124 2335 140
rect 2369 1090 2503 1118
rect 2369 1056 2387 1090
rect 2421 1084 2503 1090
rect 2421 1056 2537 1084
rect 2600 1732 2745 1739
rect 2600 1698 2612 1732
rect 2646 1698 2699 1732
rect 2733 1698 2745 1732
rect 2600 1194 2745 1698
rect 2779 1694 2813 1728
rect 2779 1626 2813 1660
rect 2779 1558 2813 1569
rect 2779 1490 2813 1497
rect 2779 1422 2813 1456
rect 2779 1354 2813 1388
rect 2779 1304 2813 1320
rect 2848 1830 2956 1851
rect 2848 1796 2885 1830
rect 2919 1796 2956 1830
rect 2848 1762 2956 1796
rect 2848 1728 2885 1762
rect 2919 1728 2956 1762
rect 2848 1694 2956 1728
rect 2848 1660 2885 1694
rect 2919 1660 2956 1694
rect 2848 1626 2956 1660
rect 2848 1592 2885 1626
rect 2919 1592 2956 1626
rect 2848 1558 2956 1592
rect 2848 1524 2885 1558
rect 2919 1524 2956 1558
rect 2848 1490 2956 1524
rect 2848 1456 2885 1490
rect 2919 1456 2956 1490
rect 2848 1422 2956 1456
rect 2848 1388 2885 1422
rect 2919 1388 2956 1422
rect 2848 1354 2956 1388
rect 2848 1320 2885 1354
rect 2919 1320 2956 1354
rect 2848 1305 2956 1320
rect 2991 1830 3025 1846
rect 2991 1762 3025 1796
rect 2991 1694 3025 1728
rect 2991 1626 3025 1660
rect 2991 1558 3025 1586
rect 2991 1490 3025 1514
rect 2991 1422 3025 1456
rect 2991 1354 3025 1388
rect 2885 1304 2919 1305
rect 2991 1304 3025 1320
rect 3131 1830 3165 1842
rect 3131 1758 3165 1784
rect 3131 1686 3165 1716
rect 3131 1614 3165 1648
rect 3131 1546 3165 1580
rect 3131 1478 3165 1512
rect 3131 1410 3165 1444
rect 3131 1342 3165 1376
rect 3131 1244 3165 1308
rect 2971 1194 3009 1196
rect 2600 1160 2756 1194
rect 2790 1160 2824 1194
rect 2858 1160 2874 1194
rect 2930 1162 2937 1194
rect 2980 1162 3009 1194
rect 2930 1160 2946 1162
rect 2980 1160 3014 1162
rect 3048 1160 3064 1194
rect 2600 1103 2835 1160
rect 2930 1103 3049 1160
rect 2600 1069 2695 1103
rect 2729 1069 2785 1103
rect 2819 1069 2835 1103
rect 2908 1069 2924 1103
rect 2958 1069 2999 1103
rect 3033 1069 3049 1103
rect 2369 1050 2537 1056
rect 2369 1022 2503 1050
rect 2369 988 2387 1022
rect 2421 1016 2503 1022
rect 2421 988 2537 1016
rect 2369 982 2537 988
rect 2369 954 2503 982
rect 2369 920 2387 954
rect 2421 948 2503 954
rect 2421 920 2537 948
rect 2369 914 2537 920
rect 2369 880 2503 914
rect 2369 846 2537 880
rect 2369 830 2503 846
rect 2369 796 2387 830
rect 2421 812 2503 830
rect 2634 1006 2668 1022
rect 2740 1006 2778 1035
rect 2634 955 2668 972
rect 2634 883 2668 904
rect 2634 820 2668 836
rect 2774 1001 2778 1006
rect 2846 1006 2880 1022
rect 2740 938 2774 972
rect 2740 870 2774 904
rect 2740 820 2774 836
rect 2950 1006 2988 1035
rect 2950 1001 2952 1006
rect 2846 955 2880 972
rect 2846 883 2880 904
rect 2846 820 2880 836
rect 2986 1001 2988 1006
rect 3058 1006 3092 1022
rect 2952 938 2986 972
rect 2952 870 2986 904
rect 2952 820 2986 836
rect 3058 955 3092 972
rect 3058 883 3092 904
rect 3058 820 3092 836
rect 2421 796 2537 812
rect 2369 778 2537 796
rect 2369 762 2503 778
rect 2369 728 2387 762
rect 2421 744 2503 762
rect 2421 728 2537 744
rect 2369 710 2537 728
rect 2369 694 2503 710
rect 2369 660 2387 694
rect 2421 676 2503 694
rect 2421 660 2537 676
rect 2369 642 2537 660
rect 2369 608 2503 642
rect 2369 574 2537 608
rect 2369 570 2503 574
rect 2369 536 2387 570
rect 2421 540 2503 570
rect 2421 536 2537 540
rect 2369 506 2537 536
rect 2369 502 2503 506
rect 2369 468 2387 502
rect 2421 472 2503 502
rect 2421 468 2537 472
rect 2369 452 2537 468
rect 2369 400 2387 452
rect 2421 404 2503 452
rect 2421 400 2537 404
rect 2369 380 2537 400
rect 2369 346 2387 380
rect 2421 346 2503 380
rect 2369 336 2503 346
rect 2369 310 2537 336
rect 2369 276 2387 310
rect 2421 302 2537 310
rect 2421 276 2503 302
rect 2369 268 2503 276
rect 2369 242 2537 268
rect 2369 208 2387 242
rect 2421 234 2537 242
rect 2421 208 2503 234
rect 2369 200 2503 208
rect 2369 174 2537 200
rect 2369 140 2387 174
rect 2421 166 2537 174
rect 2421 140 2503 166
rect 2369 132 2503 140
rect 2369 124 2537 132
rect 2503 108 2537 124
rect 1312 86 2058 90
rect 51 30 486 64
rect 520 30 554 64
rect 588 30 604 64
rect 1312 52 1328 86
rect 1362 52 1396 86
rect 1430 52 1464 86
rect 1498 52 1532 86
rect 1566 52 1600 86
rect 1634 52 1668 86
rect 1702 52 1736 86
rect 1770 52 1804 86
rect 1838 52 1872 86
rect 1906 52 1940 86
rect 1974 52 2008 86
rect 2042 52 2058 86
rect 1312 26 2058 52
rect 2251 66 2267 86
rect 2301 66 2335 86
rect 2251 40 2262 66
rect 2301 52 2334 66
rect 2369 52 2385 86
rect 2296 32 2334 52
rect 2368 40 2385 52
<< viali >>
rect 2279 2354 2313 2388
rect 2351 2354 2385 2388
rect 781 1774 815 1805
rect 781 1771 815 1774
rect 781 1706 815 1733
rect 781 1699 815 1706
rect 217 1281 323 1387
rect 393 1348 427 1382
rect 465 1348 571 1382
rect 41 1064 75 1098
rect 113 1064 147 1098
rect 494 1310 571 1348
rect 494 1276 600 1310
rect 641 1265 747 1443
rect 88 984 122 1018
rect 160 984 169 1018
rect 169 984 194 1018
rect -17 284 17 294
rect -17 260 17 284
rect -17 188 17 222
rect -17 116 17 150
rect 274 910 278 944
rect 278 910 308 944
rect 346 910 380 944
rect 482 1058 516 1092
rect 554 1058 588 1092
rect 957 1409 991 1443
rect 957 1337 991 1371
rect 957 1265 991 1299
rect 1519 1777 1553 1811
rect 1591 1782 1625 1811
rect 1591 1777 1609 1782
rect 1609 1777 1625 1782
rect 709 910 743 944
rect 781 910 815 944
rect 853 1006 869 1018
rect 869 1006 887 1018
rect 853 984 887 1006
rect 925 984 959 1018
rect 1103 984 1137 1018
rect 1175 984 1209 1018
rect 1002 938 1018 944
rect 1018 938 1036 944
rect 1002 910 1036 938
rect 1074 910 1108 944
rect 425 278 459 294
rect 425 260 459 278
rect 425 210 459 222
rect 425 188 459 210
rect 959 346 967 452
rect 967 346 1137 452
rect 717 264 751 294
rect 717 260 751 264
rect 425 116 459 150
rect 717 190 751 222
rect 717 188 751 190
rect 717 116 751 150
rect 1495 988 1529 1022
rect 1495 920 1529 950
rect 1495 916 1529 920
rect 1937 1912 2043 2090
rect 2091 1562 2125 1595
rect 2091 1561 2125 1562
rect 2091 1494 2125 1523
rect 2091 1489 2125 1494
rect 2202 1409 2236 1443
rect 2202 1370 2215 1371
rect 2215 1370 2236 1371
rect 2202 1337 2236 1370
rect 2202 1268 2236 1299
rect 2202 1265 2215 1268
rect 2215 1265 2236 1268
rect 2301 1562 2335 1595
rect 2301 1561 2335 1562
rect 2301 1494 2335 1523
rect 2301 1489 2335 1494
rect 2849 1923 2883 1957
rect 2922 1923 2956 1957
rect 2849 1851 2883 1885
rect 2922 1851 2956 1885
rect 2387 1409 2421 1443
rect 2503 1424 2537 1443
rect 2503 1409 2537 1424
rect 2387 1370 2421 1371
rect 2387 1337 2421 1370
rect 2503 1356 2537 1371
rect 2503 1337 2537 1356
rect 2387 1268 2421 1299
rect 2387 1265 2421 1268
rect 2503 1288 2537 1299
rect 2503 1265 2537 1288
rect 2203 434 2237 452
rect 2203 418 2215 434
rect 2215 418 2237 434
rect 2203 346 2237 380
rect 2301 988 2335 1022
rect 2301 920 2335 950
rect 2301 916 2335 920
rect 2612 1698 2646 1732
rect 2699 1698 2733 1732
rect 2779 1592 2813 1603
rect 2779 1569 2813 1592
rect 2779 1524 2813 1531
rect 2779 1497 2813 1524
rect 2991 1592 3025 1620
rect 2991 1586 3025 1592
rect 2991 1524 3025 1548
rect 2991 1514 3025 1524
rect 3131 1818 3165 1830
rect 3131 1796 3165 1818
rect 3131 1750 3165 1758
rect 3131 1724 3165 1750
rect 3131 1682 3165 1686
rect 3131 1652 3165 1682
rect 3131 1580 3165 1614
rect 2937 1194 2971 1196
rect 3009 1194 3043 1196
rect 2937 1162 2946 1194
rect 2946 1162 2971 1194
rect 3009 1162 3014 1194
rect 3014 1162 3043 1194
rect 2706 1001 2740 1035
rect 2634 938 2668 955
rect 2634 921 2668 938
rect 2634 870 2668 883
rect 2634 849 2668 870
rect 2778 1001 2812 1035
rect 2916 1001 2950 1035
rect 2846 938 2880 955
rect 2846 921 2880 938
rect 2846 870 2880 883
rect 2846 849 2880 870
rect 2988 1001 3022 1035
rect 3058 938 3092 955
rect 3058 921 3092 938
rect 3058 870 3092 883
rect 3058 849 3092 870
rect 2387 434 2421 452
rect 2387 418 2421 434
rect 2503 438 2537 452
rect 2503 418 2537 438
rect 2387 346 2421 380
rect 2503 370 2537 380
rect 2503 346 2537 370
rect 2262 52 2267 66
rect 2267 52 2296 66
rect 2334 52 2335 66
rect 2335 52 2368 66
rect 2262 32 2296 52
rect 2334 32 2368 52
<< metal1 >>
rect 2267 2388 2354 2400
rect 2267 2354 2279 2388
rect 2313 2354 2351 2388
rect 2267 2348 2354 2354
rect 2406 2348 2418 2400
rect 2470 2348 2476 2400
rect 738 2090 3312 2246
rect 738 1912 1937 2090
rect 2043 1957 3312 2090
rect 2043 1923 2849 1957
rect 2883 1923 2922 1957
rect 2956 1923 3312 1957
rect 2043 1912 2525 1923
rect 738 1898 2525 1912
tri 2525 1898 2550 1923 nw
tri 2755 1839 2839 1923 ne
rect 2839 1885 3312 1923
rect 2839 1851 2849 1885
rect 2883 1851 2922 1885
rect 2956 1851 3312 1885
rect 2839 1839 3312 1851
rect 775 1811 1637 1817
rect 775 1805 1519 1811
rect 775 1771 781 1805
rect 815 1777 1519 1805
rect 1553 1777 1591 1811
rect 1625 1777 1637 1811
tri 3059 1779 3119 1839 ne
rect 3119 1830 3177 1839
rect 3119 1796 3131 1830
rect 3165 1796 3177 1830
rect 815 1771 1637 1777
rect 775 1733 821 1771
tri 821 1737 855 1771 nw
rect 3119 1758 3177 1796
tri 3177 1779 3237 1839 nw
rect 775 1699 781 1733
rect 815 1699 821 1733
rect 775 1687 821 1699
rect 2378 1733 2953 1739
rect 2378 1692 2395 1733
tri 2378 1675 2395 1692 ne
rect 2447 1681 2459 1733
rect 2511 1732 2953 1733
rect 2511 1698 2612 1732
rect 2646 1698 2699 1732
rect 2733 1728 2953 1732
tri 2953 1728 2964 1739 sw
rect 2733 1698 2964 1728
rect 2511 1692 2964 1698
rect 2395 1675 2511 1681
tri 2511 1675 2528 1692 nw
tri 2930 1658 2964 1692 ne
tri 2964 1658 3034 1728 sw
rect 681 1499 699 1642
tri 617 1455 661 1499 se
rect 661 1455 699 1499
tri 699 1455 886 1642 sw
tri 2964 1640 2982 1658 ne
rect 2982 1652 3034 1658
rect 2770 1609 2822 1615
rect 2079 1595 2347 1601
rect 2079 1561 2091 1595
rect 2125 1561 2301 1595
rect 2335 1561 2347 1595
rect 2079 1523 2347 1561
rect 2079 1489 2091 1523
rect 2125 1489 2301 1523
rect 2335 1489 2347 1523
rect 2079 1483 2347 1489
rect 2770 1543 2822 1557
rect 2982 1586 2991 1600
rect 3025 1586 3034 1600
rect 2982 1560 3034 1586
rect 3119 1724 3131 1758
rect 3165 1724 3177 1758
rect 3119 1686 3177 1724
rect 3119 1652 3131 1686
rect 3165 1652 3177 1686
rect 3119 1614 3177 1652
rect 3119 1580 3131 1614
rect 3165 1580 3177 1614
rect 3119 1511 3177 1580
rect 2982 1502 3034 1508
rect 2770 1485 2822 1491
rect -96 1443 3312 1455
rect -96 1387 641 1443
rect -96 1281 217 1387
rect 323 1382 641 1387
rect 323 1348 393 1382
rect 427 1348 465 1382
rect 323 1281 494 1348
rect 571 1310 641 1382
rect -96 1276 494 1281
rect 600 1276 641 1310
rect -96 1265 641 1276
rect 747 1409 957 1443
rect 991 1409 2202 1443
rect 2236 1409 2387 1443
rect 2421 1409 2503 1443
rect 2537 1409 3312 1443
rect 747 1371 3312 1409
rect 747 1337 957 1371
rect 991 1337 2202 1371
rect 2236 1337 2387 1371
rect 2421 1337 2503 1371
rect 2537 1337 3312 1371
rect 747 1299 3312 1337
rect 747 1265 957 1299
rect 991 1265 2202 1299
rect 2236 1265 2387 1299
rect 2421 1265 2503 1299
rect 2537 1265 3312 1299
rect -96 1253 3312 1265
rect 2843 1215 2895 1221
tri 2895 1202 2914 1221 sw
rect 2895 1196 3055 1202
rect 2895 1163 2937 1196
rect 2843 1162 2937 1163
rect 2971 1162 3009 1196
rect 3043 1162 3055 1196
rect 2843 1156 3055 1162
rect 2843 1151 2895 1156
rect 2731 1119 2783 1125
rect 29 1098 600 1104
rect 29 1064 41 1098
rect 75 1064 113 1098
rect 147 1092 600 1098
rect 147 1064 482 1092
rect 29 1058 482 1064
rect 516 1058 554 1092
rect 588 1058 600 1092
rect 29 1052 600 1058
tri 2695 1041 2731 1077 se
tri 2895 1130 2921 1156 nw
rect 2843 1093 2895 1099
rect 2943 1119 2995 1125
rect 2731 1053 2783 1067
rect 2694 1035 2731 1041
tri 2783 1041 2819 1077 sw
tri 2904 1041 2943 1080 se
rect 2943 1053 2995 1067
rect 2783 1035 2824 1041
rect 76 1018 1221 1024
rect 76 984 88 1018
rect 122 984 160 1018
rect 194 984 853 1018
rect 887 984 925 1018
rect 959 984 1103 1018
rect 1137 984 1175 1018
rect 1209 984 1221 1018
rect 76 978 1221 984
rect 1489 1022 2347 1034
rect 1489 988 1495 1022
rect 1529 988 2301 1022
rect 2335 988 2347 1022
rect 2694 1001 2706 1035
rect 2812 1001 2824 1035
rect 2694 995 2824 1001
rect 2904 1035 2943 1041
tri 2995 1041 3034 1080 sw
rect 2995 1035 3034 1041
rect 2904 1001 2916 1035
rect 3022 1001 3034 1035
rect 2904 995 3034 1001
rect 1489 950 2347 988
rect 262 944 1120 950
rect 262 910 274 944
rect 308 910 346 944
rect 380 910 709 944
rect 743 910 781 944
rect 815 910 1002 944
rect 1036 910 1074 944
rect 1108 910 1120 944
rect 262 904 1120 910
rect 1489 916 1495 950
rect 1529 916 2301 950
rect 2335 916 2347 950
rect 1489 904 2347 916
rect 2628 961 3148 967
rect 2628 955 2885 961
rect 2628 921 2634 955
rect 2668 921 2846 955
rect 2880 921 2885 955
rect 2628 909 2885 921
rect 2937 909 2993 961
rect 3045 955 3148 961
rect 3045 921 3058 955
rect 3092 921 3148 955
rect 3045 909 3148 921
rect 2628 889 3148 909
rect 2628 883 2885 889
rect 2628 849 2634 883
rect 2668 849 2846 883
rect 2880 849 2885 883
rect 2628 837 2885 849
rect 2937 837 2993 889
rect 3045 883 3148 889
rect 3045 849 3058 883
rect 3092 849 3148 883
rect 3045 837 3148 849
rect 50 452 2885 464
rect 50 346 959 452
rect 1137 418 2203 452
rect 2237 418 2387 452
rect 2421 418 2503 452
rect 2537 418 2885 452
rect 1137 412 2885 418
rect 2937 412 2993 464
rect 3045 412 3312 464
rect 1137 386 3312 412
rect 1137 380 2885 386
rect 1137 346 2203 380
rect 2237 346 2387 380
rect 2421 346 2503 380
rect 2537 346 2885 380
rect 50 334 2885 346
rect 2937 334 2993 386
rect 3045 334 3312 386
rect -179 294 3312 306
rect -179 260 -17 294
rect 17 260 425 294
rect 459 260 717 294
rect 751 260 3312 294
rect -179 222 3312 260
rect -179 188 -17 222
rect 17 188 425 222
rect 459 188 717 222
rect 751 188 3312 222
rect -179 150 3312 188
rect -179 116 -17 150
rect 17 116 425 150
rect 459 116 717 150
rect 751 116 3312 150
rect -179 104 3312 116
tri 2680 72 2683 75 se
rect 2683 72 2689 75
rect 2250 66 2689 72
rect 2250 32 2262 66
rect 2296 32 2334 66
rect 2368 32 2689 66
rect 2250 26 2689 32
tri 2680 23 2683 26 ne
rect 2683 23 2689 26
rect 2741 23 2755 75
rect 2807 23 2813 75
<< via1 >>
rect 2354 2388 2406 2400
rect 2354 2354 2385 2388
rect 2385 2354 2406 2388
rect 2354 2348 2406 2354
rect 2418 2348 2470 2400
rect 2395 1681 2447 1733
rect 2459 1681 2511 1733
rect 2982 1620 3034 1652
rect 2770 1603 2822 1609
rect 2770 1569 2779 1603
rect 2779 1569 2813 1603
rect 2813 1569 2822 1603
rect 2770 1557 2822 1569
rect 2770 1531 2822 1543
rect 2770 1497 2779 1531
rect 2779 1497 2813 1531
rect 2813 1497 2822 1531
rect 2982 1600 2991 1620
rect 2991 1600 3025 1620
rect 3025 1600 3034 1620
rect 2982 1548 3034 1560
rect 2982 1514 2991 1548
rect 2991 1514 3025 1548
rect 3025 1514 3034 1548
rect 2982 1508 3034 1514
rect 2770 1491 2822 1497
rect 2843 1163 2895 1215
rect 2731 1067 2783 1119
rect 2843 1099 2895 1151
rect 2731 1035 2783 1053
rect 2943 1067 2995 1119
rect 2731 1001 2740 1035
rect 2740 1001 2778 1035
rect 2778 1001 2783 1035
rect 2943 1035 2995 1053
rect 2943 1001 2950 1035
rect 2950 1001 2988 1035
rect 2988 1001 2995 1035
rect 2885 909 2937 961
rect 2993 909 3045 961
rect 2885 837 2937 889
rect 2993 837 3045 889
rect 2885 412 2937 464
rect 2993 412 3045 464
rect 2885 334 2937 386
rect 2993 334 3045 386
rect 2689 23 2741 75
rect 2755 23 2807 75
<< metal2 >>
rect 2348 2348 2354 2400
rect 2406 2348 2418 2400
rect 2470 2348 2482 2400
tri 2393 2323 2418 2348 ne
tri 2395 1739 2418 1762 se
rect 2418 1739 2482 2348
tri 2850 2240 2884 2274 ne
tri 2482 1739 2511 1768 sw
rect 2395 1733 2511 1739
rect 2447 1681 2459 1733
rect 2395 1675 2511 1681
rect 2770 1609 2822 1615
rect 2770 1543 2822 1557
tri 2731 1358 2770 1397 se
rect 2770 1383 2822 1491
rect 2770 1358 2783 1383
rect 2731 1119 2783 1358
tri 2783 1344 2822 1383 nw
tri 2843 1284 2884 1325 se
rect 2884 1303 2936 2326
rect 2884 1284 2895 1303
rect 2843 1215 2895 1284
tri 2895 1262 2936 1303 nw
rect 2982 1652 3034 1658
rect 2982 1560 3034 1600
rect 2843 1151 2895 1163
rect 2843 1093 2895 1099
tri 2943 1231 2982 1270 se
rect 2982 1256 3034 1508
rect 2982 1231 2995 1256
rect 2943 1119 2995 1231
tri 2995 1217 3034 1256 nw
rect 2731 1053 2783 1067
tri 2697 75 2731 109 se
rect 2731 75 2783 1001
rect 2943 1053 2995 1067
rect 2943 995 2995 1001
rect 2879 909 2885 961
rect 2937 909 2993 961
rect 3045 909 3051 961
rect 2879 889 3051 909
rect 2879 837 2885 889
rect 2937 837 2993 889
rect 3045 837 3051 889
rect 2879 464 3051 837
rect 2879 412 2885 464
rect 2937 412 2993 464
rect 3045 412 3051 464
rect 2879 386 3051 412
rect 2879 334 2885 386
rect 2937 334 2993 386
rect 3045 334 3051 386
tri 2783 75 2813 105 sw
rect 2683 23 2689 75
rect 2741 23 2755 75
rect 2807 23 2813 75
use sky130_fd_pr__nfet_01v8__example_55959141808375  sky130_fd_pr__nfet_01v8__example_55959141808375_0
timestamp 1676037725
transform 1 0 2679 0 1 824
box -1 0 369 1
use sky130_fd_pr__nfet_01v8__example_55959141808376  sky130_fd_pr__nfet_01v8__example_55959141808376_0
timestamp 1676037725
transform 1 0 1620 0 -1 2202
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808377  sky130_fd_pr__nfet_01v8__example_55959141808377_0
timestamp 1676037725
transform -1 0 1411 0 -1 2202
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808379  sky130_fd_pr__nfet_01v8__example_55959141808379_0
timestamp 1676037725
transform -1 0 206 0 -1 1282
box -1 0 121 1
use sky130_fd_pr__nfet_01v8__example_55959141808380  sky130_fd_pr__nfet_01v8__example_55959141808380_0
timestamp 1676037725
transform 1 0 262 0 -1 1282
box -1 0 121 1
use sky130_fd_pr__nfet_01v8__example_55959141808381  sky130_fd_pr__nfet_01v8__example_55959141808381_0
timestamp 1676037725
transform -1 0 946 0 -1 1222
box -1 0 121 1
use sky130_fd_pr__nfet_01v8__example_55959141808382  sky130_fd_pr__nfet_01v8__example_55959141808382_0
timestamp 1676037725
transform 1 0 1002 0 -1 2024
box -1 0 121 1
use sky130_fd_pr__nfet_01v8__example_55959141808383  sky130_fd_pr__nfet_01v8__example_55959141808383_0
timestamp 1676037725
transform -1 0 946 0 -1 2024
box -1 0 121 1
use sky130_fd_pr__nfet_01v8__example_55959141808384  sky130_fd_pr__nfet_01v8__example_55959141808384_0
timestamp 1676037725
transform 1 0 1002 0 -1 1222
box -1 0 121 1
use sky130_fd_pr__nfet_01v8__example_55959141808386  sky130_fd_pr__nfet_01v8__example_55959141808386_0
timestamp 1676037725
transform 1 0 1304 0 1 648
box -1 0 417 1
use sky130_fd_pr__nfet_01v8__example_55959141808386  sky130_fd_pr__nfet_01v8__example_55959141808386_1
timestamp 1676037725
transform 1 0 1304 0 1 128
box -1 0 417 1
use sky130_fd_pr__nfet_01v8__example_55959141808386  sky130_fd_pr__nfet_01v8__example_55959141808386_2
timestamp 1676037725
transform 1 0 1304 0 1 388
box -1 0 417 1
use sky130_fd_pr__nfet_01v8__example_55959141808386  sky130_fd_pr__nfet_01v8__example_55959141808386_3
timestamp 1676037725
transform 1 0 1304 0 1 908
box -1 0 417 1
use sky130_fd_pr__nfet_01v8__example_55959141808387  sky130_fd_pr__nfet_01v8__example_55959141808387_0
timestamp 1676037725
transform 1 0 1900 0 1 2002
box -1 0 181 1
use sky130_fd_pr__nfet_01v8__example_55959141808387  sky130_fd_pr__nfet_01v8__example_55959141808387_1
timestamp 1676037725
transform 1 0 1900 0 1 1222
box -1 0 181 1
use sky130_fd_pr__nfet_01v8__example_55959141808387  sky130_fd_pr__nfet_01v8__example_55959141808387_2
timestamp 1676037725
transform 1 0 1900 0 1 1742
box -1 0 181 1
use sky130_fd_pr__nfet_01v8__example_55959141808387  sky130_fd_pr__nfet_01v8__example_55959141808387_3
timestamp 1676037725
transform 1 0 1900 0 1 388
box -1 0 181 1
use sky130_fd_pr__nfet_01v8__example_55959141808387  sky130_fd_pr__nfet_01v8__example_55959141808387_4
timestamp 1676037725
transform 1 0 1900 0 1 1482
box -1 0 181 1
use sky130_fd_pr__nfet_01v8__example_55959141808387  sky130_fd_pr__nfet_01v8__example_55959141808387_5
timestamp 1676037725
transform 1 0 1900 0 1 128
box -1 0 181 1
use sky130_fd_pr__nfet_01v8__example_55959141808387  sky130_fd_pr__nfet_01v8__example_55959141808387_6
timestamp 1676037725
transform 1 0 1900 0 1 648
box -1 0 181 1
use sky130_fd_pr__nfet_01v8__example_55959141808387  sky130_fd_pr__nfet_01v8__example_55959141808387_7
timestamp 1676037725
transform 1 0 1900 0 1 908
box -1 0 181 1
use sky130_fd_pr__nfet_01v8__example_55959141808388  sky130_fd_pr__nfet_01v8__example_55959141808388_0
timestamp 1676037725
transform 1 0 2260 0 1 908
box -1 0 117 1
use sky130_fd_pr__nfet_01v8__example_55959141808388  sky130_fd_pr__nfet_01v8__example_55959141808388_1
timestamp 1676037725
transform 1 0 2260 0 1 648
box -1 0 117 1
use sky130_fd_pr__nfet_01v8__example_55959141808388  sky130_fd_pr__nfet_01v8__example_55959141808388_2
timestamp 1676037725
transform 1 0 2260 0 1 1482
box -1 0 117 1
use sky130_fd_pr__nfet_01v8__example_55959141808388  sky130_fd_pr__nfet_01v8__example_55959141808388_3
timestamp 1676037725
transform 1 0 2260 0 1 1222
box -1 0 117 1
use sky130_fd_pr__nfet_01v8__example_55959141808388  sky130_fd_pr__nfet_01v8__example_55959141808388_4
timestamp 1676037725
transform 1 0 2260 0 1 2002
box -1 0 117 1
use sky130_fd_pr__nfet_01v8__example_55959141808388  sky130_fd_pr__nfet_01v8__example_55959141808388_5
timestamp 1676037725
transform 1 0 2260 0 1 1742
box -1 0 117 1
use sky130_fd_pr__nfet_01v8__example_55959141808388  sky130_fd_pr__nfet_01v8__example_55959141808388_6
timestamp 1676037725
transform 1 0 2260 0 1 128
box -1 0 117 1
use sky130_fd_pr__nfet_01v8__example_55959141808388  sky130_fd_pr__nfet_01v8__example_55959141808388_7
timestamp 1676037725
transform 1 0 2260 0 1 388
box -1 0 117 1
use sky130_fd_pr__pfet_01v8__example_55959141808389  sky130_fd_pr__pfet_01v8__example_55959141808389_0
timestamp 1676037725
transform 1 0 2824 0 -1 1842
box -1 0 157 1
use sky130_fd_pr__pfet_01v8__example_55959141808390  sky130_fd_pr__pfet_01v8__example_55959141808390_0
timestamp 1676037725
transform 1 0 28 0 -1 432
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808391  sky130_fd_pr__pfet_01v8__example_55959141808391_0
timestamp 1676037725
transform 1 0 28 0 -1 859
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808392  sky130_fd_pr__pfet_01v8__example_55959141808392_0
timestamp 1676037725
transform 1 0 470 0 -1 732
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808393  sky130_fd_pr__pfet_01v8__example_55959141808393_0
timestamp 1676037725
transform -1 0 414 0 -1 732
box -1 0 101 1
use sky130_fd_pr__tpl1__example_55959141808374  sky130_fd_pr__tpl1__example_55959141808374_0
timestamp 1676037725
transform -1 0 1161 0 1 92
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_0
timestamp 1676037725
transform 0 -1 2335 -1 0 1022
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_1
timestamp 1676037725
transform 0 -1 1529 -1 0 1022
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_2
timestamp 1676037725
transform 1 0 1103 0 1 984
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_3
timestamp 1676037725
transform -1 0 815 0 1 910
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_4
timestamp 1676037725
transform 0 1 2203 -1 0 452
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_5
timestamp 1676037725
transform 0 1 2503 -1 0 452
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_6
timestamp 1676037725
transform -1 0 1108 0 1 910
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_7
timestamp 1676037725
transform 0 -1 2537 -1 0 452
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_8
timestamp 1676037725
transform -1 0 959 0 1 984
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_9
timestamp 1676037725
transform 1 0 482 0 1 1058
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_10
timestamp 1676037725
transform 0 1 2387 -1 0 452
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_11
timestamp 1676037725
transform -1 0 600 0 1 1276
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_12
timestamp 1676037725
transform -1 0 380 0 1 910
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_13
timestamp 1676037725
transform -1 0 147 0 -1 1098
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_14
timestamp 1676037725
transform 1 0 1519 0 -1 1811
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_15
timestamp 1676037725
transform 0 1 781 1 0 1699
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_16
timestamp 1676037725
transform -1 0 194 0 1 984
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_17
timestamp 1676037725
transform 1 0 2279 0 1 2354
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180857  sky130_fd_pr__via_l1m1__example_5595914180857_0
timestamp 1676037725
transform 0 -1 747 -1 0 1443
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180858  sky130_fd_pr__via_l1m1__example_5595914180858_0
timestamp 1676037725
transform 0 1 217 -1 0 1387
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180878  sky130_fd_pr__via_l1m1__example_5595914180878_0
timestamp 1676037725
transform 1 0 2091 0 -1 1595
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180878  sky130_fd_pr__via_l1m1__example_5595914180878_1
timestamp 1676037725
transform 1 0 2301 0 -1 1595
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_0
timestamp 1676037725
transform 0 -1 2236 -1 0 1443
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_1
timestamp 1676037725
transform 0 -1 2421 -1 0 1443
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_2
timestamp 1676037725
transform 0 -1 751 1 0 116
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_3
timestamp 1676037725
transform 0 1 2503 -1 0 1443
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_4
timestamp 1676037725
transform 0 -1 17 1 0 116
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_5
timestamp 1676037725
transform 0 -1 459 1 0 116
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_6
timestamp 1676037725
transform -1 0 571 0 -1 1382
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_7
timestamp 1676037725
transform 0 -1 991 -1 0 1443
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808264  sky130_fd_pr__via_l1m1__example_55959141808264_0
timestamp 1676037725
transform -1 0 2043 0 -1 2090
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808264  sky130_fd_pr__via_l1m1__example_55959141808264_1
timestamp 1676037725
transform 0 1 959 -1 0 452
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_0
timestamp 1676037725
transform 1 0 2348 0 1 2348
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808271  sky130_fd_pr__via_m1m2__example_55959141808271_0
timestamp 1676037725
transform 0 1 2395 -1 0 1739
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_0
timestamp 1676037725
transform 0 1 1002 1 0 922
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_1
timestamp 1676037725
transform 0 1 853 1 0 922
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_0
timestamp 1676037725
transform 0 1 1923 1 0 2228
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_1
timestamp 1676037725
transform 0 1 2251 1 0 36
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_2
timestamp 1676037725
transform 0 1 2251 1 0 2228
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_3
timestamp 1676037725
transform 0 1 1002 -1 0 2122
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_4
timestamp 1676037725
transform 0 1 812 -1 0 2122
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_5
timestamp 1676037725
transform 0 1 470 1 0 14
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_6
timestamp 1676037725
transform 0 1 1923 1 0 1132
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808272  sky130_fd_pr__via_pol1__example_55959141808272_0
timestamp 1676037725
transform 0 -1 1719 -1 0 2294
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808273  sky130_fd_pr__via_pol1__example_55959141808273_0
timestamp 1676037725
transform 0 1 1312 1 0 36
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808373  sky130_fd_pr__via_pol1__example_55959141808373_0
timestamp 1676037725
transform 1 0 262 0 -1 1026
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808373  sky130_fd_pr__via_pol1__example_55959141808373_1
timestamp 1676037725
transform 0 1 51 -1 0 1046
box 0 0 1 1
<< labels >>
flabel metal2 s 2885 2290 2935 2320 3 FreeSans 300 180 0 0 IN
port 1 nsew
flabel locali s 413 1105 448 1151 7 FreeSans 300 180 0 0 OUT_H_N
port 3 nsew
flabel locali s 812 2333 852 2379 3 FreeSans 300 180 0 0 RST_H
port 4 nsew
flabel locali s 1096 2333 1136 2379 7 FreeSans 300 180 0 0 SET_H
port 5 nsew
flabel locali s 1496 2245 1536 2277 0 FreeSans 200 0 0 0 HLD_H_N
port 6 nsew
flabel metal1 s 3277 104 3312 306 7 FreeSans 300 180 0 0 VCC_IO
port 7 nsew
flabel metal1 s 50 334 85 464 3 FreeSans 300 180 0 0 VGND
port 8 nsew
flabel metal1 s -179 104 -144 306 3 FreeSans 300 180 0 0 VCC_IO
port 7 nsew
flabel metal1 s 3277 334 3312 464 7 FreeSans 300 180 0 0 VGND
port 8 nsew
flabel metal1 s 543 1052 578 1104 7 FreeSans 400 180 0 0 OUT_H
port 9 nsew
flabel metal1 s 3277 1253 3312 1455 7 FreeSans 300 180 0 0 VGND
port 8 nsew
flabel metal1 s 3277 1898 3312 2246 7 FreeSans 300 0 0 0 VPWR_KA
port 10 nsew
flabel metal1 s 738 1898 773 2246 3 FreeSans 300 180 0 0 VPWR_KA
port 10 nsew
flabel metal1 s -96 1253 -56 1455 3 FreeSans 300 180 0 0 VGND
port 8 nsew
flabel comment s 870 1048 870 1048 0 FreeSans 300 0 0 0 FBK_N
flabel comment s 1065 1048 1065 1048 0 FreeSans 300 0 0 0 FBK
flabel comment s 766 836 766 836 0 FreeSans 300 180 0 0 IN_I
flabel comment s 1516 2251 1516 2251 0 FreeSans 200 180 0 0 HLD_H_N
flabel comment s 1405 1655 1405 1655 0 FreeSans 300 0 0 0 IN_I_N
flabel comment s 1512 1295 1512 1295 0 FreeSans 200 0 0 0 TO HVNATIVES
flabel comment s 1142 1338 1142 1338 0 FreeSans 300 90 0 0 FBK_N
flabel comment s 812 1318 812 1318 0 FreeSans 300 270 0 0 FBK
flabel comment s 388 727 388 727 0 FreeSans 200 0 0 0 OUT_H_N
flabel comment s 1197 1497 1197 1497 0 FreeSans 300 180 0 0 FBK
flabel comment s 2578 63 2578 63 0 FreeSans 400 0 0 0 IN_I
flabel comment s 1213 1832 1213 1832 0 FreeSans 300 180 0 0 FBK_N
<< properties >>
string GDS_END 48622460
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 48593242
<< end >>
