magic
tech sky130A
magscale 1 2
timestamp 1698769616
<< nwell >>
rect 1066 106885 108874 107451
rect 1066 105797 108874 106363
rect 1066 104709 108874 105275
rect 1066 103621 108874 104187
rect 1066 102533 108874 103099
rect 1066 101445 108874 102011
rect 1066 100357 108874 100923
rect 1066 99269 108874 99835
rect 1066 98181 108874 98747
rect 1066 97093 108874 97659
rect 1066 96005 108874 96571
rect 1066 94917 108874 95483
rect 1066 93829 108874 94395
rect 1066 92741 108874 93307
rect 1066 91653 108874 92219
rect 1066 90565 108874 91131
rect 1066 89477 108874 90043
rect 1066 88389 108874 88955
rect 1066 87301 108874 87867
rect 1066 86213 108874 86779
rect 1066 85125 108874 85691
rect 1066 84037 108874 84603
rect 1066 82949 108874 83515
rect 1066 81861 108874 82427
rect 1066 80773 108874 81339
rect 1066 79685 108874 80251
rect 1066 78597 108874 79163
rect 1066 77509 108874 78075
rect 1066 76421 108874 76987
rect 1066 75333 108874 75899
rect 1066 74245 108874 74811
rect 1066 73157 108874 73723
rect 1066 72069 108874 72635
rect 1066 70981 108874 71547
rect 1066 69893 108874 70459
rect 1066 68805 108874 69371
rect 1066 67717 108874 68283
rect 1066 66629 108874 67195
rect 1066 65541 108874 66107
rect 1066 64453 108874 65019
rect 1066 63365 108874 63931
rect 1066 62277 108874 62843
rect 1066 61189 108874 61755
rect 1066 60101 108874 60667
rect 1066 59013 108874 59579
rect 1066 57925 108874 58491
rect 1066 56837 108874 57403
rect 1066 55749 108874 56315
rect 1066 54661 108874 55227
rect 1066 53573 108874 54139
rect 1066 52485 108874 53051
rect 1066 51397 108874 51963
rect 1066 50309 108874 50875
rect 1066 49221 108874 49787
rect 1066 48133 108874 48699
rect 1066 47045 108874 47611
rect 1066 45957 108874 46523
rect 1066 44869 108874 45435
rect 1066 43781 108874 44347
rect 1066 42693 108874 43259
rect 1066 41605 108874 42171
rect 1066 40517 108874 41083
rect 1066 39429 108874 39995
rect 1066 38341 108874 38907
rect 1066 37253 108874 37819
rect 1066 36165 108874 36731
rect 1066 35077 108874 35643
rect 1066 33989 108874 34555
rect 1066 32901 108874 33467
rect 1066 31813 108874 32379
rect 1066 30725 108874 31291
rect 1066 29637 108874 30203
rect 1066 28549 108874 29115
rect 1066 27461 108874 28027
rect 1066 26373 108874 26939
rect 1066 25285 108874 25851
rect 1066 24197 108874 24763
rect 1066 23109 108874 23675
rect 1066 22021 108874 22587
rect 1066 20933 108874 21499
rect 1066 19845 108874 20411
rect 1066 18757 108874 19323
rect 1066 17669 108874 18235
rect 1066 16581 108874 17147
rect 1066 15493 108874 16059
rect 1066 14405 108874 14971
rect 1066 13317 108874 13883
rect 1066 12229 108874 12795
rect 1066 11141 108874 11707
rect 1066 10053 108874 10619
rect 1066 8965 108874 9531
rect 1066 7877 108874 8443
rect 1066 6789 108874 7355
rect 1066 5701 108874 6267
rect 1066 4613 108874 5179
rect 1066 3525 108874 4091
rect 1066 2437 108874 3003
<< obsli1 >>
rect 1104 2159 108836 107729
<< obsm1 >>
rect 1104 76 109098 109132
<< metal2 >>
rect 3054 109200 3110 110000
rect 7378 109200 7434 110000
rect 11702 109200 11758 110000
rect 16026 109200 16082 110000
rect 20350 109200 20406 110000
rect 24674 109200 24730 110000
rect 28998 109200 29054 110000
rect 33322 109200 33378 110000
rect 37646 109200 37702 110000
rect 41970 109200 42026 110000
rect 46294 109200 46350 110000
rect 50618 109200 50674 110000
rect 54942 109200 54998 110000
rect 59266 109200 59322 110000
rect 63590 109200 63646 110000
rect 67914 109200 67970 110000
rect 72238 109200 72294 110000
rect 76562 109200 76618 110000
rect 80886 109200 80942 110000
rect 85210 109200 85266 110000
rect 89534 109200 89590 110000
rect 93858 109200 93914 110000
rect 98182 109200 98238 110000
rect 102506 109200 102562 110000
rect 106830 109200 106886 110000
rect 1766 0 1822 800
rect 3330 0 3386 800
rect 4894 0 4950 800
rect 6458 0 6514 800
rect 8022 0 8078 800
rect 9586 0 9642 800
rect 11150 0 11206 800
rect 12714 0 12770 800
rect 14278 0 14334 800
rect 15842 0 15898 800
rect 17406 0 17462 800
rect 18970 0 19026 800
rect 20534 0 20590 800
rect 22098 0 22154 800
rect 23662 0 23718 800
rect 25226 0 25282 800
rect 26790 0 26846 800
rect 28354 0 28410 800
rect 29918 0 29974 800
rect 31482 0 31538 800
rect 33046 0 33102 800
rect 34610 0 34666 800
rect 36174 0 36230 800
rect 37738 0 37794 800
rect 39302 0 39358 800
rect 40866 0 40922 800
rect 42430 0 42486 800
rect 43994 0 44050 800
rect 45558 0 45614 800
rect 47122 0 47178 800
rect 48686 0 48742 800
rect 50250 0 50306 800
rect 51814 0 51870 800
rect 53378 0 53434 800
rect 54942 0 54998 800
rect 56506 0 56562 800
rect 58070 0 58126 800
rect 59634 0 59690 800
rect 61198 0 61254 800
rect 62762 0 62818 800
rect 64326 0 64382 800
rect 65890 0 65946 800
rect 67454 0 67510 800
rect 69018 0 69074 800
rect 70582 0 70638 800
rect 72146 0 72202 800
rect 73710 0 73766 800
rect 75274 0 75330 800
rect 76838 0 76894 800
rect 78402 0 78458 800
rect 79966 0 80022 800
rect 81530 0 81586 800
rect 83094 0 83150 800
rect 84658 0 84714 800
rect 86222 0 86278 800
rect 87786 0 87842 800
rect 89350 0 89406 800
rect 90914 0 90970 800
rect 92478 0 92534 800
rect 94042 0 94098 800
rect 95606 0 95662 800
rect 97170 0 97226 800
rect 98734 0 98790 800
rect 100298 0 100354 800
rect 101862 0 101918 800
rect 103426 0 103482 800
rect 104990 0 105046 800
rect 106554 0 106610 800
rect 108118 0 108174 800
<< obsm2 >>
rect 1768 109144 2998 109200
rect 3166 109144 7322 109200
rect 7490 109144 11646 109200
rect 11814 109144 15970 109200
rect 16138 109144 20294 109200
rect 20462 109144 24618 109200
rect 24786 109144 28942 109200
rect 29110 109144 33266 109200
rect 33434 109144 37590 109200
rect 37758 109144 41914 109200
rect 42082 109144 46238 109200
rect 46406 109144 50562 109200
rect 50730 109144 54886 109200
rect 55054 109144 59210 109200
rect 59378 109144 63534 109200
rect 63702 109144 67858 109200
rect 68026 109144 72182 109200
rect 72350 109144 76506 109200
rect 76674 109144 80830 109200
rect 80998 109144 85154 109200
rect 85322 109144 89478 109200
rect 89646 109144 93802 109200
rect 93970 109144 98126 109200
rect 98294 109144 102450 109200
rect 102618 109144 106774 109200
rect 106942 109144 109094 109200
rect 1768 856 109094 109144
rect 1878 70 3274 856
rect 3442 70 4838 856
rect 5006 70 6402 856
rect 6570 70 7966 856
rect 8134 70 9530 856
rect 9698 70 11094 856
rect 11262 70 12658 856
rect 12826 70 14222 856
rect 14390 70 15786 856
rect 15954 70 17350 856
rect 17518 70 18914 856
rect 19082 70 20478 856
rect 20646 70 22042 856
rect 22210 70 23606 856
rect 23774 70 25170 856
rect 25338 70 26734 856
rect 26902 70 28298 856
rect 28466 70 29862 856
rect 30030 70 31426 856
rect 31594 70 32990 856
rect 33158 70 34554 856
rect 34722 70 36118 856
rect 36286 70 37682 856
rect 37850 70 39246 856
rect 39414 70 40810 856
rect 40978 70 42374 856
rect 42542 70 43938 856
rect 44106 70 45502 856
rect 45670 70 47066 856
rect 47234 70 48630 856
rect 48798 70 50194 856
rect 50362 70 51758 856
rect 51926 70 53322 856
rect 53490 70 54886 856
rect 55054 70 56450 856
rect 56618 70 58014 856
rect 58182 70 59578 856
rect 59746 70 61142 856
rect 61310 70 62706 856
rect 62874 70 64270 856
rect 64438 70 65834 856
rect 66002 70 67398 856
rect 67566 70 68962 856
rect 69130 70 70526 856
rect 70694 70 72090 856
rect 72258 70 73654 856
rect 73822 70 75218 856
rect 75386 70 76782 856
rect 76950 70 78346 856
rect 78514 70 79910 856
rect 80078 70 81474 856
rect 81642 70 83038 856
rect 83206 70 84602 856
rect 84770 70 86166 856
rect 86334 70 87730 856
rect 87898 70 89294 856
rect 89462 70 90858 856
rect 91026 70 92422 856
rect 92590 70 93986 856
rect 94154 70 95550 856
rect 95718 70 97114 856
rect 97282 70 98678 856
rect 98846 70 100242 856
rect 100410 70 101806 856
rect 101974 70 103370 856
rect 103538 70 104934 856
rect 105102 70 106498 856
rect 106666 70 108062 856
rect 108230 70 109094 856
<< metal3 >>
rect 109200 106496 110000 106616
rect 109200 103368 110000 103488
rect 109200 100240 110000 100360
rect 109200 97112 110000 97232
rect 109200 93984 110000 94104
rect 109200 90856 110000 90976
rect 109200 87728 110000 87848
rect 109200 84600 110000 84720
rect 109200 81472 110000 81592
rect 109200 78344 110000 78464
rect 109200 75216 110000 75336
rect 109200 72088 110000 72208
rect 109200 68960 110000 69080
rect 109200 65832 110000 65952
rect 109200 62704 110000 62824
rect 109200 59576 110000 59696
rect 109200 56448 110000 56568
rect 109200 53320 110000 53440
rect 109200 50192 110000 50312
rect 109200 47064 110000 47184
rect 109200 43936 110000 44056
rect 109200 40808 110000 40928
rect 109200 37680 110000 37800
rect 109200 34552 110000 34672
rect 109200 31424 110000 31544
rect 109200 28296 110000 28416
rect 109200 25168 110000 25288
rect 109200 22040 110000 22160
rect 109200 18912 110000 19032
rect 109200 15784 110000 15904
rect 109200 12656 110000 12776
rect 109200 9528 110000 9648
rect 109200 6400 110000 6520
rect 109200 3272 110000 3392
<< obsm3 >>
rect 4210 106696 109200 107745
rect 4210 106416 109120 106696
rect 4210 103568 109200 106416
rect 4210 103288 109120 103568
rect 4210 100440 109200 103288
rect 4210 100160 109120 100440
rect 4210 97312 109200 100160
rect 4210 97032 109120 97312
rect 4210 94184 109200 97032
rect 4210 93904 109120 94184
rect 4210 91056 109200 93904
rect 4210 90776 109120 91056
rect 4210 87928 109200 90776
rect 4210 87648 109120 87928
rect 4210 84800 109200 87648
rect 4210 84520 109120 84800
rect 4210 81672 109200 84520
rect 4210 81392 109120 81672
rect 4210 78544 109200 81392
rect 4210 78264 109120 78544
rect 4210 75416 109200 78264
rect 4210 75136 109120 75416
rect 4210 72288 109200 75136
rect 4210 72008 109120 72288
rect 4210 69160 109200 72008
rect 4210 68880 109120 69160
rect 4210 66032 109200 68880
rect 4210 65752 109120 66032
rect 4210 62904 109200 65752
rect 4210 62624 109120 62904
rect 4210 59776 109200 62624
rect 4210 59496 109120 59776
rect 4210 56648 109200 59496
rect 4210 56368 109120 56648
rect 4210 53520 109200 56368
rect 4210 53240 109120 53520
rect 4210 50392 109200 53240
rect 4210 50112 109120 50392
rect 4210 47264 109200 50112
rect 4210 46984 109120 47264
rect 4210 44136 109200 46984
rect 4210 43856 109120 44136
rect 4210 41008 109200 43856
rect 4210 40728 109120 41008
rect 4210 37880 109200 40728
rect 4210 37600 109120 37880
rect 4210 34752 109200 37600
rect 4210 34472 109120 34752
rect 4210 31624 109200 34472
rect 4210 31344 109120 31624
rect 4210 28496 109200 31344
rect 4210 28216 109120 28496
rect 4210 25368 109200 28216
rect 4210 25088 109120 25368
rect 4210 22240 109200 25088
rect 4210 21960 109120 22240
rect 4210 19112 109200 21960
rect 4210 18832 109120 19112
rect 4210 15984 109200 18832
rect 4210 15704 109120 15984
rect 4210 12856 109200 15704
rect 4210 12576 109120 12856
rect 4210 9728 109200 12576
rect 4210 9448 109120 9728
rect 4210 6600 109200 9448
rect 4210 6320 109120 6600
rect 4210 3472 109200 6320
rect 4210 3192 109120 3472
rect 4210 1939 109200 3192
<< metal4 >>
rect 4208 2128 4528 107760
rect 19568 2128 19888 107760
rect 34928 2128 35248 107760
rect 50288 2128 50608 107760
rect 65648 2128 65968 107760
rect 81008 2128 81328 107760
rect 96368 2128 96688 107760
<< obsm4 >>
rect 22323 3299 34848 106317
rect 35328 3299 50208 106317
rect 50688 3299 65568 106317
rect 66048 3299 80928 106317
rect 81408 3299 96288 106317
rect 96768 3299 104085 106317
<< labels >>
rlabel metal2 s 3054 109200 3110 110000 6 buttons
port 1 nsew signal input
rlabel metal2 s 1766 0 1822 800 6 clk
port 2 nsew signal input
rlabel metal2 s 9586 0 9642 800 6 i_wb_addr[0]
port 3 nsew signal input
rlabel metal2 s 25226 0 25282 800 6 i_wb_addr[10]
port 4 nsew signal input
rlabel metal2 s 26790 0 26846 800 6 i_wb_addr[11]
port 5 nsew signal input
rlabel metal2 s 28354 0 28410 800 6 i_wb_addr[12]
port 6 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 i_wb_addr[13]
port 7 nsew signal input
rlabel metal2 s 31482 0 31538 800 6 i_wb_addr[14]
port 8 nsew signal input
rlabel metal2 s 33046 0 33102 800 6 i_wb_addr[15]
port 9 nsew signal input
rlabel metal2 s 34610 0 34666 800 6 i_wb_addr[16]
port 10 nsew signal input
rlabel metal2 s 36174 0 36230 800 6 i_wb_addr[17]
port 11 nsew signal input
rlabel metal2 s 37738 0 37794 800 6 i_wb_addr[18]
port 12 nsew signal input
rlabel metal2 s 39302 0 39358 800 6 i_wb_addr[19]
port 13 nsew signal input
rlabel metal2 s 11150 0 11206 800 6 i_wb_addr[1]
port 14 nsew signal input
rlabel metal2 s 40866 0 40922 800 6 i_wb_addr[20]
port 15 nsew signal input
rlabel metal2 s 42430 0 42486 800 6 i_wb_addr[21]
port 16 nsew signal input
rlabel metal2 s 43994 0 44050 800 6 i_wb_addr[22]
port 17 nsew signal input
rlabel metal2 s 45558 0 45614 800 6 i_wb_addr[23]
port 18 nsew signal input
rlabel metal2 s 47122 0 47178 800 6 i_wb_addr[24]
port 19 nsew signal input
rlabel metal2 s 48686 0 48742 800 6 i_wb_addr[25]
port 20 nsew signal input
rlabel metal2 s 50250 0 50306 800 6 i_wb_addr[26]
port 21 nsew signal input
rlabel metal2 s 51814 0 51870 800 6 i_wb_addr[27]
port 22 nsew signal input
rlabel metal2 s 53378 0 53434 800 6 i_wb_addr[28]
port 23 nsew signal input
rlabel metal2 s 54942 0 54998 800 6 i_wb_addr[29]
port 24 nsew signal input
rlabel metal2 s 12714 0 12770 800 6 i_wb_addr[2]
port 25 nsew signal input
rlabel metal2 s 56506 0 56562 800 6 i_wb_addr[30]
port 26 nsew signal input
rlabel metal2 s 58070 0 58126 800 6 i_wb_addr[31]
port 27 nsew signal input
rlabel metal2 s 14278 0 14334 800 6 i_wb_addr[3]
port 28 nsew signal input
rlabel metal2 s 15842 0 15898 800 6 i_wb_addr[4]
port 29 nsew signal input
rlabel metal2 s 17406 0 17462 800 6 i_wb_addr[5]
port 30 nsew signal input
rlabel metal2 s 18970 0 19026 800 6 i_wb_addr[6]
port 31 nsew signal input
rlabel metal2 s 20534 0 20590 800 6 i_wb_addr[7]
port 32 nsew signal input
rlabel metal2 s 22098 0 22154 800 6 i_wb_addr[8]
port 33 nsew signal input
rlabel metal2 s 23662 0 23718 800 6 i_wb_addr[9]
port 34 nsew signal input
rlabel metal2 s 4894 0 4950 800 6 i_wb_cyc
port 35 nsew signal input
rlabel metal2 s 59634 0 59690 800 6 i_wb_data[0]
port 36 nsew signal input
rlabel metal2 s 75274 0 75330 800 6 i_wb_data[10]
port 37 nsew signal input
rlabel metal2 s 76838 0 76894 800 6 i_wb_data[11]
port 38 nsew signal input
rlabel metal2 s 78402 0 78458 800 6 i_wb_data[12]
port 39 nsew signal input
rlabel metal2 s 79966 0 80022 800 6 i_wb_data[13]
port 40 nsew signal input
rlabel metal2 s 81530 0 81586 800 6 i_wb_data[14]
port 41 nsew signal input
rlabel metal2 s 83094 0 83150 800 6 i_wb_data[15]
port 42 nsew signal input
rlabel metal2 s 84658 0 84714 800 6 i_wb_data[16]
port 43 nsew signal input
rlabel metal2 s 86222 0 86278 800 6 i_wb_data[17]
port 44 nsew signal input
rlabel metal2 s 87786 0 87842 800 6 i_wb_data[18]
port 45 nsew signal input
rlabel metal2 s 89350 0 89406 800 6 i_wb_data[19]
port 46 nsew signal input
rlabel metal2 s 61198 0 61254 800 6 i_wb_data[1]
port 47 nsew signal input
rlabel metal2 s 90914 0 90970 800 6 i_wb_data[20]
port 48 nsew signal input
rlabel metal2 s 92478 0 92534 800 6 i_wb_data[21]
port 49 nsew signal input
rlabel metal2 s 94042 0 94098 800 6 i_wb_data[22]
port 50 nsew signal input
rlabel metal2 s 95606 0 95662 800 6 i_wb_data[23]
port 51 nsew signal input
rlabel metal2 s 97170 0 97226 800 6 i_wb_data[24]
port 52 nsew signal input
rlabel metal2 s 98734 0 98790 800 6 i_wb_data[25]
port 53 nsew signal input
rlabel metal2 s 100298 0 100354 800 6 i_wb_data[26]
port 54 nsew signal input
rlabel metal2 s 101862 0 101918 800 6 i_wb_data[27]
port 55 nsew signal input
rlabel metal2 s 103426 0 103482 800 6 i_wb_data[28]
port 56 nsew signal input
rlabel metal2 s 104990 0 105046 800 6 i_wb_data[29]
port 57 nsew signal input
rlabel metal2 s 62762 0 62818 800 6 i_wb_data[2]
port 58 nsew signal input
rlabel metal2 s 106554 0 106610 800 6 i_wb_data[30]
port 59 nsew signal input
rlabel metal2 s 108118 0 108174 800 6 i_wb_data[31]
port 60 nsew signal input
rlabel metal2 s 64326 0 64382 800 6 i_wb_data[3]
port 61 nsew signal input
rlabel metal2 s 65890 0 65946 800 6 i_wb_data[4]
port 62 nsew signal input
rlabel metal2 s 67454 0 67510 800 6 i_wb_data[5]
port 63 nsew signal input
rlabel metal2 s 69018 0 69074 800 6 i_wb_data[6]
port 64 nsew signal input
rlabel metal2 s 70582 0 70638 800 6 i_wb_data[7]
port 65 nsew signal input
rlabel metal2 s 72146 0 72202 800 6 i_wb_data[8]
port 66 nsew signal input
rlabel metal2 s 73710 0 73766 800 6 i_wb_data[9]
port 67 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 i_wb_stb
port 68 nsew signal input
rlabel metal2 s 8022 0 8078 800 6 i_wb_we
port 69 nsew signal input
rlabel metal2 s 7378 109200 7434 110000 6 led_enb[0]
port 70 nsew signal output
rlabel metal2 s 50618 109200 50674 110000 6 led_enb[10]
port 71 nsew signal output
rlabel metal2 s 54942 109200 54998 110000 6 led_enb[11]
port 72 nsew signal output
rlabel metal2 s 11702 109200 11758 110000 6 led_enb[1]
port 73 nsew signal output
rlabel metal2 s 16026 109200 16082 110000 6 led_enb[2]
port 74 nsew signal output
rlabel metal2 s 20350 109200 20406 110000 6 led_enb[3]
port 75 nsew signal output
rlabel metal2 s 24674 109200 24730 110000 6 led_enb[4]
port 76 nsew signal output
rlabel metal2 s 28998 109200 29054 110000 6 led_enb[5]
port 77 nsew signal output
rlabel metal2 s 33322 109200 33378 110000 6 led_enb[6]
port 78 nsew signal output
rlabel metal2 s 37646 109200 37702 110000 6 led_enb[7]
port 79 nsew signal output
rlabel metal2 s 41970 109200 42026 110000 6 led_enb[8]
port 80 nsew signal output
rlabel metal2 s 46294 109200 46350 110000 6 led_enb[9]
port 81 nsew signal output
rlabel metal2 s 59266 109200 59322 110000 6 leds[0]
port 82 nsew signal output
rlabel metal2 s 102506 109200 102562 110000 6 leds[10]
port 83 nsew signal output
rlabel metal2 s 106830 109200 106886 110000 6 leds[11]
port 84 nsew signal output
rlabel metal2 s 63590 109200 63646 110000 6 leds[1]
port 85 nsew signal output
rlabel metal2 s 67914 109200 67970 110000 6 leds[2]
port 86 nsew signal output
rlabel metal2 s 72238 109200 72294 110000 6 leds[3]
port 87 nsew signal output
rlabel metal2 s 76562 109200 76618 110000 6 leds[4]
port 88 nsew signal output
rlabel metal2 s 80886 109200 80942 110000 6 leds[5]
port 89 nsew signal output
rlabel metal2 s 85210 109200 85266 110000 6 leds[6]
port 90 nsew signal output
rlabel metal2 s 89534 109200 89590 110000 6 leds[7]
port 91 nsew signal output
rlabel metal2 s 93858 109200 93914 110000 6 leds[8]
port 92 nsew signal output
rlabel metal2 s 98182 109200 98238 110000 6 leds[9]
port 93 nsew signal output
rlabel metal3 s 109200 3272 110000 3392 6 o_wb_ack
port 94 nsew signal output
rlabel metal3 s 109200 9528 110000 9648 6 o_wb_data[0]
port 95 nsew signal output
rlabel metal3 s 109200 40808 110000 40928 6 o_wb_data[10]
port 96 nsew signal output
rlabel metal3 s 109200 43936 110000 44056 6 o_wb_data[11]
port 97 nsew signal output
rlabel metal3 s 109200 47064 110000 47184 6 o_wb_data[12]
port 98 nsew signal output
rlabel metal3 s 109200 50192 110000 50312 6 o_wb_data[13]
port 99 nsew signal output
rlabel metal3 s 109200 53320 110000 53440 6 o_wb_data[14]
port 100 nsew signal output
rlabel metal3 s 109200 56448 110000 56568 6 o_wb_data[15]
port 101 nsew signal output
rlabel metal3 s 109200 59576 110000 59696 6 o_wb_data[16]
port 102 nsew signal output
rlabel metal3 s 109200 62704 110000 62824 6 o_wb_data[17]
port 103 nsew signal output
rlabel metal3 s 109200 65832 110000 65952 6 o_wb_data[18]
port 104 nsew signal output
rlabel metal3 s 109200 68960 110000 69080 6 o_wb_data[19]
port 105 nsew signal output
rlabel metal3 s 109200 12656 110000 12776 6 o_wb_data[1]
port 106 nsew signal output
rlabel metal3 s 109200 72088 110000 72208 6 o_wb_data[20]
port 107 nsew signal output
rlabel metal3 s 109200 75216 110000 75336 6 o_wb_data[21]
port 108 nsew signal output
rlabel metal3 s 109200 78344 110000 78464 6 o_wb_data[22]
port 109 nsew signal output
rlabel metal3 s 109200 81472 110000 81592 6 o_wb_data[23]
port 110 nsew signal output
rlabel metal3 s 109200 84600 110000 84720 6 o_wb_data[24]
port 111 nsew signal output
rlabel metal3 s 109200 87728 110000 87848 6 o_wb_data[25]
port 112 nsew signal output
rlabel metal3 s 109200 90856 110000 90976 6 o_wb_data[26]
port 113 nsew signal output
rlabel metal3 s 109200 93984 110000 94104 6 o_wb_data[27]
port 114 nsew signal output
rlabel metal3 s 109200 97112 110000 97232 6 o_wb_data[28]
port 115 nsew signal output
rlabel metal3 s 109200 100240 110000 100360 6 o_wb_data[29]
port 116 nsew signal output
rlabel metal3 s 109200 15784 110000 15904 6 o_wb_data[2]
port 117 nsew signal output
rlabel metal3 s 109200 103368 110000 103488 6 o_wb_data[30]
port 118 nsew signal output
rlabel metal3 s 109200 106496 110000 106616 6 o_wb_data[31]
port 119 nsew signal output
rlabel metal3 s 109200 18912 110000 19032 6 o_wb_data[3]
port 120 nsew signal output
rlabel metal3 s 109200 22040 110000 22160 6 o_wb_data[4]
port 121 nsew signal output
rlabel metal3 s 109200 25168 110000 25288 6 o_wb_data[5]
port 122 nsew signal output
rlabel metal3 s 109200 28296 110000 28416 6 o_wb_data[6]
port 123 nsew signal output
rlabel metal3 s 109200 31424 110000 31544 6 o_wb_data[7]
port 124 nsew signal output
rlabel metal3 s 109200 34552 110000 34672 6 o_wb_data[8]
port 125 nsew signal output
rlabel metal3 s 109200 37680 110000 37800 6 o_wb_data[9]
port 126 nsew signal output
rlabel metal3 s 109200 6400 110000 6520 6 o_wb_stall
port 127 nsew signal output
rlabel metal2 s 3330 0 3386 800 6 reset
port 128 nsew signal input
rlabel metal4 s 4208 2128 4528 107760 6 vccd1
port 129 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 107760 6 vccd1
port 129 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 107760 6 vccd1
port 129 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 107760 6 vccd1
port 129 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 107760 6 vssd1
port 130 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 107760 6 vssd1
port 130 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 107760 6 vssd1
port 130 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 110000 110000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 27455834
string GDS_FILE /home/bignixon/unic-cass/caravel_tutorial/caravel_user_project/openlane/wb_buttons_leds/runs/23_10_31_13_17/results/signoff/wb_buttons_leds.magic.gds
string GDS_START 1509852
<< end >>

