magic
tech sky130A
timestamp 1676037725
<< properties >>
string GDS_END 229508
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_2kbyte_1rw1r_32x512_8.gds
string GDS_START 229184
<< end >>
