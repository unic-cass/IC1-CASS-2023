* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
X0 VPWR A2 a_469_443# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X1 X a_83_283# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X2 X a_83_283# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X3 a_631_107# A2 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X4 VGND B1 a_83_283# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X5 a_83_283# B1 a_469_443# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X6 a_83_283# A1 a_631_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X7 a_469_443# A1 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
X0 Y B1 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X1 VGND A2 a_271_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X2 a_56_443# A2 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X3 a_271_107# A1 Y VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X4 a_56_443# B1 Y VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X5 VPWR A1 a_56_443# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
X0 X a_83_81# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X1 a_822_107# A2 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X2 a_316_443# B2 a_83_81# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X3 X a_83_81# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X4 a_316_443# A1 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X5 VGND B2 a_519_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X6 a_519_107# B1 a_83_81# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X7 a_83_81# A1 a_822_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X8 a_83_81# B1 a_316_443# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X9 VPWR A2 a_316_443# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
X0 VGND B2 a_204_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X1 a_33_443# B2 Y VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X2 a_502_107# A2 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X3 a_204_107# B1 Y VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X4 Y B1 a_33_443# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X5 Y A1 a_502_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X6 VPWR A2 a_33_443# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X7 a_33_443# A1 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__and2_1 A B VGND VNB VPB VPWR X
X0 VGND a_30_107# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X1 VPWR a_30_107# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X2 a_30_107# A a_183_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X3 a_183_107# B VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X4 VPWR A a_30_107# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X5 a_30_107# B VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__and3_1 A B C VGND VNB VPB VPWR X
X0 VGND a_30_517# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X1 a_201_173# B a_343_173# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X2 a_30_517# C VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X3 VPWR a_30_517# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X4 a_30_517# A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X5 VPWR B a_30_517# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X6 a_30_517# A a_201_173# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X7 a_343_173# C VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__buf_1 A VGND VNB VPB VPWR X
X0 VPWR A a_84_81# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X1 X a_84_81# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X2 VGND A a_84_81# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X3 X a_84_81# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__buf_2 A VGND VNB VPB VPWR X
X0 VPWR A a_129_279# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X1 VPWR a_129_279# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X2 X a_129_279# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X3 VGND A a_129_279# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X4 X a_129_279# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X5 VGND a_129_279# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__buf_4 A VGND VNB VPB VPWR X
X0 X a_149_81# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X1 X a_149_81# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X2 X a_149_81# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X3 X a_149_81# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X4 VGND a_149_81# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X5 VGND A a_149_81# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X6 VPWR a_149_81# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X7 VPWR A a_149_81# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X8 VGND a_149_81# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X9 VPWR a_149_81# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__buf_8 A VGND VNB VPB VPWR X
X0 a_45_443# A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X1 X a_45_443# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X2 X a_45_443# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X3 X a_45_443# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X4 X a_45_443# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X5 VGND A a_45_443# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X6 VGND a_45_443# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X7 VGND a_45_443# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X8 a_45_443# A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X9 X a_45_443# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X10 VGND a_45_443# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X11 VGND a_45_443# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X12 X a_45_443# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X13 X a_45_443# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X14 a_45_443# A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X15 VPWR A a_45_443# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X16 a_45_443# A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X17 VPWR a_45_443# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X18 VPWR a_45_443# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X19 X a_45_443# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X20 VPWR a_45_443# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X21 VPWR a_45_443# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__buf_16 A VGND VNB VPB VPWR X
X0 X a_183_141# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X1 X a_183_141# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X2 a_183_141# A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X3 VGND a_183_141# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X4 X a_183_141# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X5 VPWR A a_183_141# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X6 X a_183_141# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X7 VPWR a_183_141# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X8 a_183_141# A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X9 VPWR A a_183_141# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X10 VPWR a_183_141# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X11 VGND a_183_141# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X12 X a_183_141# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X13 VPWR A a_183_141# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X14 VPWR a_183_141# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X15 VGND a_183_141# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X16 VPWR a_183_141# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X17 VGND a_183_141# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X18 a_183_141# A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X19 VGND a_183_141# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X20 a_183_141# A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X21 X a_183_141# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X22 a_183_141# A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X23 X a_183_141# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X24 VPWR a_183_141# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X25 X a_183_141# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X26 X a_183_141# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X27 X a_183_141# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X28 X a_183_141# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X29 X a_183_141# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X30 VPWR a_183_141# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X31 X a_183_141# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X32 VPWR a_183_141# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X33 VGND A a_183_141# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X34 VGND a_183_141# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X35 a_183_141# A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X36 VPWR a_183_141# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X37 VGND A a_183_141# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X38 VGND a_183_141# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X39 X a_183_141# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X40 VGND A a_183_141# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X41 X a_183_141# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X42 VGND a_183_141# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X43 X a_183_141# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__buf_32 A VGND VNB VPB VPWR X
X0 a_183_141# A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X1 X a_183_141# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X2 VPWR a_183_141# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X3 VGND a_183_141# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X4 X a_183_141# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X5 a_183_141# A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X6 VPWR a_183_141# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X7 X a_183_141# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X8 VGND a_183_141# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X9 VGND a_183_141# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X10 VPWR A a_183_141# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X11 X a_183_141# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X12 VPWR A a_183_141# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X13 a_183_141# A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X14 X a_183_141# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X15 VPWR a_183_141# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X16 X a_183_141# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X17 X a_183_141# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X18 VPWR A a_183_141# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X19 X a_183_141# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X20 VGND A a_183_141# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X21 VPWR a_183_141# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X22 X a_183_141# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X23 VPWR A a_183_141# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X24 VPWR a_183_141# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X25 X a_183_141# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X26 X a_183_141# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X27 X a_183_141# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X28 VPWR a_183_141# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X29 X a_183_141# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X30 VPWR a_183_141# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X31 X a_183_141# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X32 VPWR a_183_141# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X33 a_183_141# A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X34 VPWR a_183_141# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X35 VGND a_183_141# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X36 VPWR a_183_141# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X37 VGND a_183_141# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X38 a_183_141# A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X39 a_183_141# A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X40 X a_183_141# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X41 VGND a_183_141# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X42 VPWR A a_183_141# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X43 X a_183_141# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X44 VGND a_183_141# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X45 a_183_141# A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X46 X a_183_141# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X47 X a_183_141# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X48 X a_183_141# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X49 VGND a_183_141# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X50 VGND a_183_141# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X51 X a_183_141# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X52 a_183_141# A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X53 X a_183_141# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X54 VGND a_183_141# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X55 X a_183_141# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X56 X a_183_141# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X57 X a_183_141# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X58 X a_183_141# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X59 VGND a_183_141# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X60 X a_183_141# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X61 VGND A a_183_141# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X62 VGND A a_183_141# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X63 VPWR a_183_141# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X64 VGND a_183_141# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X65 X a_183_141# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X66 a_183_141# A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X67 VPWR a_183_141# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X68 X a_183_141# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X69 VGND A a_183_141# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X70 VPWR a_183_141# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X71 VGND A a_183_141# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X72 VGND a_183_141# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X73 X a_183_141# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X74 a_183_141# A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X75 VPWR a_183_141# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X76 VGND a_183_141# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X77 X a_183_141# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X78 X a_183_141# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X79 VPWR a_183_141# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X80 VGND a_183_141# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X81 X a_183_141# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X82 VPWR a_183_141# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X83 VGND a_183_141# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__conb_1 VGND VNB VPB VPWR HI LO
R0 HI VPWR sky130_fd_pr__res_generic_po w=510000u l=45000u
R1 VGND LO sky130_fd_pr__res_generic_po w=510000u l=45000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__decap_4 VGND VNB VPB VPWR
X0 VGND VPWR VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=1e+06u
X1 VPWR VGND VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=1e+06u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__decap_8 VGND VNB VPB VPWR
X0 VGND VPWR VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=1e+06u
X1 VPWR VGND VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=1e+06u
X2 VPWR VGND VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=1e+06u
X3 VGND VPWR VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=1e+06u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__dfrbp_1 CLK D RESET_B VGND VNB VPB VPWR Q Q_N
X0 a_1176_466# a_350_107# a_1900_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X1 a_37_107# CLK VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X2 VGND a_2937_443# Q VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X3 a_2122_348# a_1900_107# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X4 VPWR RESET_B a_978_608# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X5 VGND a_37_107# a_350_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X6 a_978_608# a_350_107# a_1215_173# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X7 VPWR a_2937_443# Q VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X8 a_2412_107# a_1900_107# a_2122_348# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X9 a_978_608# a_37_107# a_1134_608# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X10 VPWR a_37_107# a_350_107# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X11 a_2114_107# a_2122_348# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X12 a_2937_443# a_1900_107# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X13 a_1900_107# a_350_107# a_2079_462# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X14 VPWR a_1900_107# Q_N VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X15 a_2079_462# a_2122_348# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X16 a_509_608# a_37_107# a_978_608# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X17 VGND RESET_B a_2412_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X18 VGND a_1900_107# Q_N VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X19 a_1357_173# RESET_B VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X20 VPWR a_978_608# a_1176_466# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
X21 a_1215_173# a_1176_466# a_1357_173# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X22 a_509_608# RESET_B VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X23 VGND a_978_608# a_1176_466# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X24 a_2937_443# a_1900_107# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X25 a_509_608# a_350_107# a_978_608# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X26 VGND RESET_B a_728_173# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X27 a_37_107# CLK VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X28 a_728_173# D a_509_608# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X29 a_1900_107# a_37_107# a_2114_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X30 a_1134_608# a_1176_466# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X31 a_1176_466# a_37_107# a_1900_107# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
X32 VPWR RESET_B a_2122_348# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X33 VPWR D a_509_608# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
X0 a_1233_173# RESET_B VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X1 VGND RESET_B a_2387_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X2 VPWR a_921_632# a_1119_506# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
X3 a_1091_173# a_1119_506# a_1233_173# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X4 a_30_107# CLK VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X5 a_2089_107# a_2096_417# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X6 VPWR a_30_107# a_339_537# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X7 VGND RESET_B a_637_173# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X8 VPWR RESET_B a_921_632# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X9 VGND a_30_107# a_339_537# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X10 a_452_632# RESET_B VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X11 a_2054_543# a_2096_417# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X12 a_921_632# a_339_537# a_1091_173# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X13 VPWR a_2649_207# Q VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X14 a_1875_543# a_339_537# a_2054_543# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X15 a_1119_506# a_30_107# a_1875_543# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
X16 a_2387_107# a_1875_543# a_2096_417# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X17 a_2096_417# a_1875_543# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X18 a_1077_632# a_1119_506# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X19 a_30_107# CLK VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X20 a_1119_506# a_339_537# a_1875_543# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X21 VPWR D a_452_632# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X22 a_921_632# a_30_107# a_1077_632# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X23 VPWR RESET_B a_2096_417# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X24 a_637_173# D a_452_632# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X25 a_2649_207# a_1875_543# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X26 VGND a_921_632# a_1119_506# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X27 a_2649_207# a_1875_543# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X28 a_452_632# a_339_537# a_921_632# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X29 a_1875_543# a_30_107# a_2089_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X30 VGND a_2649_207# Q VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X31 a_452_632# a_30_107# a_921_632# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__dfsbp_1 CLK D SET_B VGND VNB VPB VPWR Q Q_N
X0 a_605_109# a_339_112# a_761_109# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X1 VPWR a_761_109# a_1732_543# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
X2 a_1755_153# a_30_112# a_1874_543# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X3 a_917_109# a_959_83# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X4 VGND a_761_109# a_1642_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X5 a_1325_107# SET_B VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X6 a_1874_543# a_339_112# a_1642_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X7 a_30_112# CLK VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X8 a_2427_107# SET_B VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X9 VPWR a_3129_479# Q VPB sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
X10 a_3129_479# a_1874_543# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X11 VPWR a_30_112# a_339_112# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X12 VPWR a_761_109# a_959_83# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X13 VPWR a_1874_543# Q_N VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X14 a_2156_417# a_1874_543# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X15 a_2053_543# a_2156_417# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X16 VGND a_30_112# a_339_112# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X17 VGND a_3129_479# Q VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X18 VGND D a_605_109# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X19 a_1874_543# a_339_112# a_2053_543# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X20 a_976_543# a_959_83# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X21 a_1732_543# a_30_112# a_1874_543# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
X22 a_761_109# a_339_112# a_917_109# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X23 a_959_83# SET_B VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X24 VPWR SET_B a_1874_543# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X25 a_959_83# a_761_109# a_1325_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X26 a_2156_417# a_1874_543# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X27 a_1755_153# a_2156_417# a_2427_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X28 VPWR D a_605_109# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X29 VGND a_1874_543# Q_N VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X30 a_761_109# a_30_112# a_976_543# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X31 a_605_109# a_30_112# a_761_109# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X32 a_3129_479# a_1874_543# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X33 a_30_112# CLK VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
X0 VPWR a_30_131# a_340_593# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X1 a_2553_203# a_1787_137# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X2 VPWR a_2553_203# Q VPB sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
X3 VGND a_798_107# a_1645_137# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X4 a_958_107# a_1000_81# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X5 a_1989_203# a_2031_177# a_2131_203# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X6 a_1268_251# SET_B VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X7 a_982_529# a_1000_81# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X8 VPWR a_798_107# a_1000_81# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X9 a_1653_515# a_30_131# a_1787_137# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
X10 VGND a_1787_137# a_2031_177# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X11 a_1787_137# a_340_593# a_1989_515# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X12 a_642_107# a_340_593# a_798_107# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X13 a_2553_203# a_1787_137# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X14 a_798_107# a_30_131# a_982_529# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X15 VPWR SET_B a_1787_137# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X16 a_642_107# a_30_131# a_798_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X17 a_1645_137# a_340_593# a_1787_137# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X18 VGND a_2553_203# Q VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X19 a_2031_177# a_1787_137# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X20 a_1000_81# a_798_107# a_1268_251# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X21 a_30_131# CLK VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X22 VGND D a_642_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X23 a_2131_203# SET_B VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X24 a_1989_515# a_2031_177# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X25 a_1000_81# SET_B VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X26 VGND a_30_131# a_340_593# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X27 VPWR D a_642_107# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X28 VPWR a_798_107# a_1653_515# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
X29 a_30_131# CLK VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X30 a_798_107# a_340_593# a_958_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X31 a_1787_137# a_30_131# a_1989_203# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__dfxbp_1 CLK D VGND VNB VPB VPWR Q Q_N
X0 a_1021_111# a_1063_85# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X1 a_1669_111# a_1711_85# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X2 VPWR a_865_111# a_1063_85# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
X3 a_865_111# a_339_112# a_1021_111# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X4 a_1494_539# a_30_112# a_1669_111# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X5 VPWR D a_709_111# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X6 VPWR a_1494_539# a_1711_85# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
X7 a_1063_85# a_339_112# a_1494_539# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X8 Q a_1711_85# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X9 VGND a_865_111# a_1063_85# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X10 a_1063_85# a_30_112# a_1494_539# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
X11 VGND a_30_112# a_339_112# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X12 a_30_112# CLK VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X13 Q a_1711_85# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X14 a_2365_443# a_1711_85# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X15 a_2365_443# a_1711_85# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X16 VGND D a_709_111# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X17 VPWR a_30_112# a_339_112# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X18 a_709_111# a_339_112# a_865_111# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X19 VGND a_1494_539# a_1711_85# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X20 VPWR a_2365_443# Q_N VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X21 a_1021_539# a_1063_85# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X22 a_1669_539# a_1711_85# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X23 a_865_111# a_30_112# a_1021_539# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X24 a_1494_539# a_339_112# a_1669_539# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X25 a_30_112# CLK VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X26 a_709_111# a_30_112# a_865_111# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X27 VGND a_2365_443# Q_N VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__dfxtp_1 CLK D VGND VNB VPB VPWR Q
X0 a_780_574# a_30_127# a_982_543# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X1 VPWR a_1455_543# a_1729_87# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
X2 VGND a_1729_87# Q VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X3 a_1015_113# a_1024_371# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X4 VPWR a_780_574# a_1024_371# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
X5 a_1455_543# a_339_559# a_1731_543# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X6 VGND a_1455_543# a_1729_87# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X7 a_780_574# a_339_559# a_1015_113# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X8 a_30_127# CLK VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X9 a_1455_543# a_30_127# a_1687_113# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X10 a_605_563# a_30_127# a_780_574# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X11 a_1024_371# a_30_127# a_1455_543# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
X12 a_1024_371# a_339_559# a_1455_543# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X13 a_605_563# a_339_559# a_780_574# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X14 a_30_127# CLK VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X15 VGND a_780_574# a_1024_371# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X16 VPWR a_1729_87# Q VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X17 VPWR D a_605_563# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X18 VGND a_30_127# a_339_559# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X19 VGND D a_605_563# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X20 a_982_543# a_1024_371# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X21 a_1687_113# a_1729_87# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X22 a_1731_543# a_1729_87# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X23 VPWR a_30_127# a_339_559# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__diode_2 DIODE VGND VNB VPB VPWR
D0 VNB DIODE sky130_fd_pr__diode_pw2nd_11v0 pj=3.16e+06 area=6.072e+11
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__dlclkp_1 CLK GATE VGND VNB VPB VPWR GCLK
X0 a_303_311# a_239_419# a_1027_159# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X1 a_189_159# a_231_71# a_303_311# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X2 VGND a_1438_171# GCLK VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X3 VGND GATE a_189_159# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X4 VGND a_303_311# a_1069_133# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X5 a_189_445# a_239_419# a_303_311# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X6 VPWR GATE a_189_445# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X7 a_239_419# a_231_71# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X8 VPWR a_1438_171# GCLK VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X9 a_1438_171# CLK VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X10 a_239_419# a_231_71# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X11 a_1027_457# a_1069_133# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X12 a_1591_171# CLK VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X13 VPWR a_1069_133# a_1438_171# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X14 VPWR CLK a_231_71# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X15 a_303_311# a_231_71# a_1027_457# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X16 VPWR a_303_311# a_1069_133# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X17 VGND CLK a_231_71# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X18 a_1438_171# a_1069_133# a_1591_171# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X19 a_1027_159# a_1069_133# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__dlrtp_1 D GATE RESET_B VGND VNB VPB VPWR Q
X0 a_1096_491# a_1138_81# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X1 a_775_491# a_345_107# a_917_107# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X2 a_1096_107# a_1138_81# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X3 a_917_107# a_462_107# a_1096_491# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X4 a_775_107# a_462_107# a_917_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X5 VPWR a_917_107# a_1138_81# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X6 a_462_107# a_345_107# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X7 a_1138_81# a_917_107# a_1512_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X8 a_917_107# a_345_107# a_1096_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X9 a_462_107# a_345_107# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X10 VPWR a_1138_81# Q VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X11 a_1138_81# RESET_B VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X12 a_32_107# D VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X13 VPWR a_32_107# a_775_491# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X14 VGND GATE a_345_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X15 a_32_107# D VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X16 VGND a_32_107# a_775_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X17 VGND a_1138_81# Q VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X18 VPWR GATE a_345_107# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X19 a_1512_107# RESET_B VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__dlxtp_1 D GATE VGND VNB VPB VPWR Q
X0 a_650_107# a_384_107# a_806_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X1 a_30_443# GATE VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X2 a_962_107# a_1004_81# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X3 VPWR D a_650_107# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X4 VGND D a_650_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X5 VGND a_806_107# Q VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X6 a_1014_587# a_1004_81# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X7 VPWR a_806_107# Q VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X8 a_806_107# a_30_443# a_962_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X9 a_1004_81# a_806_107# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X10 a_30_443# GATE VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X11 VPWR a_30_443# a_384_107# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X12 a_806_107# a_384_107# a_1014_587# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X13 a_650_107# a_30_443# a_806_107# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X14 a_1004_81# a_806_107# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X15 VGND a_30_443# a_384_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__einvn_1 A TE_B VGND VNB VPB VPWR Z
X0 VGND a_30_173# a_437_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X1 a_30_173# TE_B VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X2 a_437_107# A Z VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X3 VPWR TE_B a_413_443# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X4 a_30_173# TE_B VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X5 a_413_443# A Z VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__einvp_1 A TE VGND VNB VPB VPWR Z
X0 a_413_443# A Z VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X1 a_30_189# TE VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X2 a_30_189# TE VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X3 VGND TE a_413_123# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X4 a_413_123# A Z VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X5 VPWR a_30_189# a_413_443# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__fill_1 VGND VNB VPB VPWR
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__fill_2 VGND VNB VPB VPWR
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__fill_4 VGND VNB VPB VPWR
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__fill_8 VGND VNB VPB VPWR
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__inv_1 A VGND VNB VPB VPWR Y
X0 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X1 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__inv_2 A VGND VNB VPB VPWR Y
X0 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X2 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X3 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__inv_4 A VGND VNB VPB VPWR Y
X0 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X1 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X2 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X3 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X4 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X5 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X6 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X7 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__inv_8 A VGND VNB VPB VPWR Y
X0 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X1 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X2 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X3 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X4 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X5 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X6 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X7 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X8 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X9 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X10 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X11 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X12 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X13 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X14 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X15 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__inv_16 A VGND VNB VPB VPWR Y
X0 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X1 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X2 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X3 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X4 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X5 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X6 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X7 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X8 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X9 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X10 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X11 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X12 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X13 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X14 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X15 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X16 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X17 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X18 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X19 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X20 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X21 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X22 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X23 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X24 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X25 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X26 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X27 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X28 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X29 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X30 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X31 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__lsbufhv2hv_hl_1 A LOWHVPWR VGND VNB VPB VPWR X
X0 X a_662_81# LOWHVPWR LOWHVPWR sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X1 LOWHVPWR A a_662_81# LOWHVPWR sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X2 X a_662_81# a_762_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X3 a_762_107# A a_662_81# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__lsbufhv2hv_lh_1 A LOWHVPWR VGND VNB VPB VPWR X
X0 a_847_1221# a_626_141# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=500000u
X1 a_1353_107# a_935_141# a_779_141# VNB sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=500000u
X2 VPWR a_1353_107# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X3 a_847_1221# a_626_141# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=500000u
X4 a_1353_107# a_847_1221# a_1793_563# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=1e+06u
X5 a_1353_107# a_935_141# a_779_141# VNB sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=500000u
X6 a_626_141# A LOWHVPWR LOWHVPWR sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X7 VGND a_626_141# a_847_1221# VNB sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=500000u
X8 VGND a_1353_107# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X9 a_626_141# A a_779_141# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X10 LOWHVPWR a_626_141# a_935_141# LOWHVPWR sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X11 a_779_141# a_935_141# a_1353_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=500000u
X12 a_847_1221# a_1353_107# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=1e+06u
X13 a_779_141# a_935_141# a_1353_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=500000u
X14 VGND a_626_141# a_847_1221# VNB sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=500000u
X15 a_779_141# a_626_141# a_935_141# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__lsbufhv2lv_1 A LVPWR VGND VNB VPB VPWR X
X0 a_30_207# a_30_1337# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X1 VPWR a_30_1337# a_30_207# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X2 X a_389_141# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X3 a_389_1337# a_30_1337# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X4 a_389_1337# a_30_1337# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X5 X a_389_141# LVPWR LVPWR sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X6 a_389_141# a_389_1337# LVPWR LVPWR sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X7 VGND a_30_207# a_389_141# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X8 a_389_141# a_30_207# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X9 a_389_141# a_30_207# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X10 VPWR A a_30_1337# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X11 a_30_1337# A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X12 LVPWR a_389_141# a_389_1337# LVPWR sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X13 a_389_141# a_30_207# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X14 VGND a_30_1337# a_389_1337# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X15 VGND a_30_1337# a_389_1337# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__lsbufhv2lv_simple_1 A LVPWR VGND VNB VPB VPWR X
X0 X a_662_81# a_762_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X1 a_762_107# A a_662_81# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X2 X a_662_81# LVPWR LVPWR sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X3 LVPWR A a_662_81# LVPWR sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.subckt sky130_fd_sc_hvl__lsbuflv2hv_1 A LVPWR VGND VNB VPB VPWR X
X0 VGND a_404_1133# a_504_1221# VNB sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=500000u
X1 a_504_1221# a_404_1133# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=500000u
X2 X a_1711_885# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X3 X a_1711_885# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X4 VGND A a_404_1133# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X5 a_1197_107# a_772_151# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=500000u
X6 VPWR a_1197_107# a_504_1221# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=1e+06u
X7 a_504_1221# a_404_1133# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=500000u
X8 a_1197_107# a_772_151# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=500000u
X9 a_772_151# a_404_1133# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X10 a_504_1221# a_404_1133# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=500000u
X11 VGND a_404_1133# a_504_1221# VNB sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=500000u
X12 LVPWR A a_404_1133# LVPWR sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X13 VGND a_772_151# a_1197_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=500000u
X14 VPWR a_504_1221# a_1711_885# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X15 VGND a_504_1221# a_1711_885# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X16 VGND a_772_151# a_1197_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=500000u
X17 a_772_151# a_404_1133# LVPWR LVPWR sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X18 a_1197_107# a_772_151# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=500000u
X19 VPWR a_504_1221# a_1197_107# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=1e+06u
.ends



******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__lsbuflv2hv_clkiso_hlkg_3 A SLEEP_B LVPWR VGND VNB VPB VPWR
+ X
X0 VPWR a_262_107# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=3e+06u l=500000u
X1 VGND a_528_1171# a_362_1243# VNB sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X2 a_362_133# a_528_1171# a_1472_1171# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X3 a_362_1243# a_528_1171# VGND VNB sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X4 a_362_1243# a_840_107# a_1410_571# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X5 a_1472_1171# a_528_1171# a_362_133# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X6 a_940_485# a_2092_381# a_1410_571# VPB sky130_fd_pr__pfet_g5v0d10v5 w=3e+06u l=500000u
X7 a_1472_1171# a_528_1171# LVPWR LVPWR sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X8 a_840_107# a_1472_1171# VGND VNB sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X9 VGND a_1472_1171# a_840_107# VNB sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X10 a_940_485# a_2092_381# a_1410_571# VPB sky130_fd_pr__pfet_g5v0d10v5 w=3e+06u l=500000u
X11 a_528_1171# a_3617_1198# LVPWR LVPWR sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X12 VGND a_528_1171# a_362_1243# VNB sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X13 X a_262_107# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=3e+06u l=500000u
X14 LVPWR a_3617_1198# a_528_1171# LVPWR sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X15 a_362_133# a_528_1171# a_1472_1171# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X16 a_1472_1171# a_528_1171# a_362_133# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X17 a_3617_1198# A LVPWR LVPWR sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X18 a_362_133# a_840_107# a_262_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=1e+06u l=500000u
X19 X a_262_107# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=3e+06u l=500000u
X20 LVPWR a_3617_1198# a_528_1171# LVPWR sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X21 a_528_1171# a_3617_1198# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X22 a_262_107# a_840_107# a_362_133# VNB sky130_fd_pr__nfet_g5v0d10v5 w=1e+06u l=500000u
X23 a_1410_571# a_2092_381# a_940_485# VPB sky130_fd_pr__pfet_g5v0d10v5 w=3e+06u l=500000u
X24 a_840_107# a_2092_381# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X25 a_1472_1171# a_528_1171# LVPWR LVPWR sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X26 a_362_133# a_262_107# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=1e+06u l=500000u
X27 a_840_107# a_1472_1171# VGND VNB sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X28 VGND a_3617_1198# a_528_1171# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X29 LVPWR a_528_1171# a_1472_1171# LVPWR sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X30 a_2092_381# SLEEP_B VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X31 a_528_1171# a_3617_1198# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X32 VGND a_3617_1198# a_528_1171# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X33 LVPWR a_528_1171# a_1472_1171# LVPWR sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X34 a_940_485# a_840_107# a_262_107# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X35 a_362_1243# a_528_1171# VGND VNB sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X36 VGND VGND a_362_1243# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X37 VGND a_1472_1171# a_840_107# VNB sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X38 a_2092_381# SLEEP_B VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X39 a_528_1171# a_3617_1198# LVPWR LVPWR sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X40 a_3617_1198# A VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X41 LVPWR A a_3617_1198# LVPWR sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X42 VGND A a_3617_1198# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X43 X a_262_107# a_362_133# VNB sky130_fd_pr__nfet_g5v0d10v5 w=1e+06u l=500000u
X44 a_262_107# a_840_107# a_940_485# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X45 a_1410_571# a_362_1243# a_840_107# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X46 a_1410_571# a_2092_381# a_940_485# VPB sky130_fd_pr__pfet_g5v0d10v5 w=3e+06u l=500000u
X47 X a_262_107# a_362_133# VNB sky130_fd_pr__nfet_g5v0d10v5 w=1e+06u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__lsbuflv2hv_isosrchvaon_1 A SLEEP_B LVPWR VGND VNB VPB VPWR
+ X
X0 a_176_993# a_229_967# a_341_485# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=2e+06u
X1 a_341_183# SLEEP_B a_507_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X2 X a_229_967# a_341_485# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X3 a_188_1293# a_553_1225# a_229_967# VNB sky130_fd_pr__nfet_g5v0d10v5 w=1e+06u l=500000u
X4 a_341_183# A a_241_1225# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X5 a_188_1293# a_241_1225# a_176_993# VNB sky130_fd_pr__nfet_g5v0d10v5 w=1e+06u l=500000u
X6 a_341_485# SLEEP_B a_507_107# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X7 a_188_1293# SLEEP_B a_341_183# VNB sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=600000u
X8 a_553_1225# a_241_1225# LVPWR LVPWR sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X9 a_553_1225# a_241_1225# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X10 a_341_183# SLEEP_B a_188_1293# VNB sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=600000u
X11 a_176_993# a_241_1225# a_188_1293# VNB sky130_fd_pr__nfet_g5v0d10v5 w=1e+06u l=500000u
X12 a_341_485# a_176_993# a_229_967# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=2e+06u
X13 X a_229_967# a_341_183# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X14 a_176_993# a_507_107# a_341_183# VNB sky130_fd_pr__nfet_g5v0d10v5 w=1e+06u l=800000u
X15 LVPWR A a_241_1225# LVPWR sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X16 a_229_967# a_553_1225# a_188_1293# VNB sky130_fd_pr__nfet_g5v0d10v5 w=1e+06u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__lsbuflv2hv_symmetric_1 A LVPWR VGND VNB VPB VPWR X
X0 a_1400_777# a_1406_429# a_1197_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=500000u
X1 VGND a_1406_429# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X2 a_1406_429# a_816_1221# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X3 a_573_897# A a_686_151# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X4 a_573_897# A LVPWR LVPWR sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X5 a_1606_563# a_816_1221# a_1400_777# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=1e+06u
X6 VGND a_573_897# a_816_1221# VNB sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=500000u
X7 a_816_1221# a_1400_777# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X8 a_816_1221# a_573_897# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=500000u
X9 a_686_151# a_573_897# a_772_151# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X10 LVPWR a_573_897# a_772_151# LVPWR sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X11 a_686_151# a_772_151# a_1197_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=500000u
X12 a_816_1221# a_1406_429# a_1606_563# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=1e+06u
X13 VPWR a_1400_777# a_816_1221# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X14 VPWR a_1406_429# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X15 a_1406_429# a_816_1221# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X16 a_1197_107# a_772_151# a_686_151# VNB sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=500000u
X17 a_1400_777# a_1406_429# a_1606_563# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X18 a_1197_107# a_1406_429# a_1400_777# VNB sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__mux2_1 A0 A1 S VGND VNB VPB VPWR X
X0 X a_94_81# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X1 a_671_107# a_713_81# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X2 a_373_491# A0 a_94_81# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X3 X a_94_81# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X4 a_373_107# A1 a_94_81# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X5 a_94_81# A1 a_671_491# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X6 a_94_81# A0 a_671_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X7 VPWR S a_373_491# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X8 VPWR S a_713_81# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X9 a_671_491# a_713_81# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X10 VGND S a_373_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X11 VGND S a_713_81# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
X0 a_30_107# S0 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X1 a_30_107# S0 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X2 a_1097_627# a_1681_89# a_1669_615# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X3 a_1281_107# A0 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X4 a_955_627# a_30_107# a_1097_627# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X5 a_481_107# S0 a_637_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X6 a_1253_627# A0 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X7 a_983_107# S0 a_1097_627# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X8 VGND a_1669_615# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X9 a_481_107# a_30_107# a_637_627# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X10 a_637_627# A3 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X11 VPWR a_1669_615# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X12 a_1097_627# S1 a_1669_615# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X13 a_1681_89# S1 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X14 VGND A2 a_339_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X15 a_339_107# a_30_107# a_481_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X16 VGND A1 a_983_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X17 VPWR A1 a_955_627# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X18 VPWR A2 a_339_627# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X19 a_1669_615# a_1681_89# a_481_107# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X20 a_1097_627# a_30_107# a_1281_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X21 a_339_627# S0 a_481_107# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X22 a_1097_627# S0 a_1253_627# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X23 a_1681_89# S1 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X24 a_637_107# A3 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X25 a_1669_615# S1 a_481_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__nand2_1 A B VGND VNB VPB VPWR Y
X0 VPWR B Y VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X1 VGND B a_233_111# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X2 a_233_111# A Y VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X3 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__nand3_1 A B C VGND VNB VPB VPWR Y
X0 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X1 VGND C a_243_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X2 VPWR C Y VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X3 a_385_107# A Y VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X4 a_243_107# B a_385_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X5 Y B VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__nor2_1 A B VGND VNB VPB VPWR Y
X0 VPWR A a_251_443# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X1 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X2 Y B VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X3 a_251_443# B Y VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__nor3_1 A B C VGND VNB VPB VPWR Y
X0 a_347_443# C Y VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X1 Y B VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X2 a_205_443# B a_347_443# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X3 VGND C Y VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X4 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X5 VPWR A a_205_443# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
X0 a_83_87# A2 a_602_443# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X1 a_460_107# A2 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X2 a_83_87# B1 a_460_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X3 X a_83_87# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X4 VGND A1 a_460_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X5 X a_83_87# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X6 a_602_443# A1 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X7 VPWR B1 a_83_87# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
X0 a_30_107# A1 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X1 VGND A2 a_30_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X2 a_205_443# A2 Y VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X3 a_30_107# B1 Y VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X4 Y B1 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X5 VPWR A1 a_205_443# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
X0 a_354_107# A2 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X1 a_87_81# A2 a_831_443# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X2 X a_87_81# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X3 VGND A1 a_354_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X4 X a_87_81# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X5 VPWR B1 a_533_443# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X6 a_354_107# B1 a_87_81# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X7 a_831_443# A1 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X8 a_87_81# B2 a_354_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X9 a_533_443# B2 a_87_81# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
X0 a_207_443# B2 Y VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X1 a_520_443# A1 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X2 Y B2 a_36_113# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X3 VGND A1 a_36_113# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X4 VPWR B1 a_207_443# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X5 a_36_113# A2 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X6 a_36_113# B1 Y VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X7 Y A2 a_520_443# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__or2_1 A B VGND VNB VPB VPWR X
X0 VPWR a_84_443# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X1 a_241_443# A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X2 a_84_443# A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X3 VGND B a_84_443# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X4 a_84_443# B a_241_443# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X5 VGND a_84_443# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__or3_1 A B C VGND VNB VPB VPWR X
X0 VGND a_30_107# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X1 VPWR a_30_107# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X2 a_30_107# C VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X3 a_30_107# C a_190_464# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X4 a_341_464# A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X5 a_30_107# A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X6 VGND B a_30_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X7 a_190_464# B a_341_464# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__probe_p_8 A VGND VNB VPB VPWR X
X0 a_45_443# A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X1 X a_45_443# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X2 X a_45_443# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X3 X a_45_443# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X4 X a_45_443# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X5 VGND A a_45_443# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X6 VGND a_45_443# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X7 VGND a_45_443# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X8 a_45_443# A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X9 X a_45_443# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X10 VGND a_45_443# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X11 VGND a_45_443# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X12 X a_45_443# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X13 X a_45_443# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X14 a_45_443# A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X15 VPWR A a_45_443# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X16 a_45_443# A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X17 VPWR a_45_443# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X18 VPWR a_45_443# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X19 X a_45_443# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X20 VPWR a_45_443# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X21 VPWR a_45_443# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__probec_p_8 A VGND VNB VPB VPWR X
X0 a_45_443# A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X1 X a_45_443# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X2 X a_45_443# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X3 X a_45_443# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X4 X a_45_443# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X5 VGND A a_45_443# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X6 VGND a_45_443# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X7 VGND a_45_443# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X8 a_45_443# A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X9 X a_45_443# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X10 VGND a_45_443# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X11 VGND a_45_443# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X12 X a_45_443# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X13 X a_45_443# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X14 a_45_443# A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X15 VPWR A a_45_443# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X16 a_45_443# A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X17 VPWR a_45_443# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X18 VPWR a_45_443# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X19 X a_45_443# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X20 VPWR a_45_443# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X21 VPWR a_45_443# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__schmittbuf_1 A VGND VNB VPB VPWR X
X0 a_117_181# A a_231_463# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X1 a_117_181# A a_217_207# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X2 a_78_463# VGND VNB sky130_fd_pr__res_generic_nd__hv w=290000u l=1.355e+06u
X3 a_64_207# VPWR VPB sky130_fd_pr__res_generic_pd__hv w=290000u l=3.11e+06u
X4 a_231_463# A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X5 a_64_207# a_117_181# a_217_207# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X6 VGND a_117_181# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X7 VPWR a_117_181# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X8 a_217_207# A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X9 a_78_463# a_117_181# a_231_463# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__sdfrbp_1 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q Q_N
X0 a_3098_107# a_2624_107# a_2841_81# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X1 VPWR SCD a_794_655# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X2 a_1999_126# a_2014_537# a_2141_126# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X3 VGND a_2624_107# Q_N VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X4 a_1972_659# a_2014_537# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X5 a_2871_543# a_2841_81# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X6 VGND CLK a_1290_126# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X7 a_2799_107# a_2841_81# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X8 a_2624_107# a_1290_126# a_2799_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X9 VPWR a_1290_126# a_1569_126# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X10 a_339_655# D a_496_655# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X11 a_1816_659# a_1290_126# a_1972_659# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X12 VPWR a_1816_659# a_2014_537# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
X13 VPWR RESET_B a_2841_81# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X14 a_794_655# a_222_131# a_339_655# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X15 a_339_655# SCE a_816_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X16 VPWR CLK a_1290_126# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X17 VPWR RESET_B a_1816_659# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X18 VGND a_1816_659# a_2014_537# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X19 VGND SCE a_222_131# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X20 a_2841_81# a_2624_107# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X21 a_3613_443# a_2624_107# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X22 a_2141_126# RESET_B VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X23 a_361_107# D a_518_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X24 a_496_655# SCE VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X25 a_339_655# RESET_B VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X26 VGND a_1290_126# a_1569_126# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X27 a_2014_537# a_1569_126# a_2624_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X28 a_2624_107# a_1569_126# a_2871_543# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X29 a_518_107# a_222_131# a_339_655# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X30 a_2014_537# a_1290_126# a_2624_107# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
X31 a_361_107# RESET_B VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X32 VGND RESET_B a_3098_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X33 a_1816_659# a_1569_126# a_1999_126# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X34 a_3613_443# a_2624_107# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X35 VPWR a_3613_443# Q VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X36 VPWR SCE a_222_131# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X37 a_339_655# a_1290_126# a_1816_659# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X38 VPWR a_2624_107# Q_N VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X39 VGND a_3613_443# Q VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X40 a_339_655# a_1569_126# a_1816_659# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X41 a_816_107# SCD a_361_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__sdfrtp_1 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q
X0 VPWR SCE a_116_451# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X1 VGND SCE a_116_451# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X2 a_1510_100# a_1212_471# a_2360_115# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X3 a_2574_543# a_2616_417# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X4 VGND RESET_B a_2904_181# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X5 a_1212_100# CLK VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X6 VGND a_3417_443# Q VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X7 a_294_126# SCE a_65_649# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X8 VPWR a_3417_443# Q VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X9 a_1610_126# RESET_B VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X10 a_3417_443# a_2360_115# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X11 a_524_649# D a_65_649# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X12 a_2360_115# a_1212_100# a_2539_181# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X13 a_137_126# RESET_B VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X14 a_2539_181# a_2616_417# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X15 a_222_649# SCD VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X16 VPWR CLK a_1212_100# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X17 a_65_649# RESET_B VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X18 a_1468_641# a_1510_100# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X19 VPWR RESET_B a_2616_417# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X20 a_3417_443# a_2360_115# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X21 a_65_649# a_116_451# a_592_126# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X22 a_1312_126# a_1212_100# a_1468_641# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X23 VPWR a_1312_126# a_1510_100# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
X24 VGND a_1312_126# a_1510_100# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X25 a_1468_126# a_1510_100# a_1610_126# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X26 a_2904_181# a_2360_115# a_2616_417# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X27 VPWR SCE a_524_649# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X28 a_65_649# a_1212_471# a_1312_126# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X29 VPWR RESET_B a_1312_126# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X30 a_2360_115# a_1212_471# a_2574_543# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X31 a_1212_471# a_1212_100# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X32 a_1312_126# a_1212_471# a_1468_126# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X33 a_1212_471# a_1212_100# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X34 a_137_126# SCD a_294_126# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X35 a_65_649# a_116_451# a_222_649# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X36 a_2616_417# a_2360_115# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X37 a_65_649# a_1212_100# a_1312_126# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X38 a_592_126# D a_137_126# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X39 a_1510_100# a_1212_100# a_2360_115# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__sdfsbp_1 CLK D SCD SCE SET_B VGND VNB VPB VPWR Q Q_N
X0 a_641_569# SCD VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X1 VGND a_972_569# a_1243_116# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X2 a_2501_543# a_972_569# a_2715_173# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X3 a_485_569# a_1243_116# a_1513_120# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X4 a_1711_94# a_1513_120# a_2077_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X5 VGND D a_348_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X6 VPWR a_2501_543# Q_N VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X7 a_348_107# a_30_569# a_485_569# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X8 a_2857_173# SET_B VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X9 VPWR CLK a_972_569# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X10 a_343_569# D a_485_569# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X11 a_1513_120# a_972_569# a_1710_556# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X12 a_2394_107# a_1243_116# a_2501_543# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X13 a_2501_543# a_1243_116# a_2687_543# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X14 a_2729_463# a_2501_543# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X15 a_3609_173# a_2501_543# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X16 VPWR a_3609_173# Q VPB sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
X17 VPWR SET_B a_2501_543# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X18 a_646_107# SCD VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X19 a_3609_173# a_2501_543# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X20 a_485_569# a_30_569# a_641_569# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X21 a_30_569# SCE VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X22 VPWR a_972_569# a_1243_116# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X23 VGND a_3609_173# Q VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X24 a_2729_463# a_2501_543# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X25 VGND CLK a_972_569# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X26 a_1669_120# a_1711_94# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X27 a_2715_173# a_2729_463# a_2857_173# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X28 a_30_569# SCE VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X29 a_1711_94# SET_B VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X30 a_1513_120# a_1243_116# a_1669_120# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X31 VPWR SCE a_343_569# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X32 a_2687_543# a_2729_463# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X33 VGND a_2501_543# Q_N VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X34 a_2359_543# a_972_569# a_2501_543# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
X35 a_1710_556# a_1711_94# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X36 a_485_569# a_972_569# a_1513_120# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X37 a_485_569# SCE a_646_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X38 a_2077_107# SET_B VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X39 VPWR a_1513_120# a_1711_94# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X40 VPWR a_1513_120# a_2359_543# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
X41 VGND a_1513_120# a_2394_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__sdfstp_1 CLK D SCD SCE SET_B VGND VNB VPB VPWR Q
X0 VGND a_2477_543# a_2698_421# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X1 a_2352_107# a_1201_123# a_2477_543# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X2 VGND a_3321_173# Q VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X3 a_30_107# SCE VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X4 a_1471_113# a_1201_123# a_1627_113# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X5 VPWR SCE a_339_569# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X6 VPWR a_1471_113# a_1669_87# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X7 a_1471_113# a_935_107# a_1686_543# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X8 VGND CLK a_935_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X9 a_2477_543# a_935_107# a_2669_173# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X10 a_339_569# D a_481_107# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X11 a_481_107# a_1201_123# a_1471_113# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X12 VPWR a_1471_113# a_2335_543# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
X13 a_481_107# a_935_107# a_1471_113# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X14 a_1669_87# SET_B VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X15 a_481_107# SCE a_637_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X16 a_2812_173# SET_B VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X17 VPWR CLK a_935_107# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X18 a_637_569# SCD VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X19 a_2656_543# a_2698_421# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X20 VGND a_1471_113# a_2352_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X21 a_1686_543# a_1669_87# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X22 a_30_107# SCE VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X23 a_2035_107# SET_B VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X24 a_1627_113# a_1669_87# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X25 VPWR SET_B a_2477_543# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X26 VGND D a_339_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X27 a_1669_87# a_1471_113# a_2035_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X28 a_339_107# a_30_107# a_481_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X29 VPWR a_3321_173# Q VPB sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
X30 a_2698_421# a_2477_543# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X31 VGND a_935_107# a_1201_123# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X32 a_2669_173# a_2698_421# a_2812_173# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X33 a_3321_173# a_2477_543# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X34 a_3321_173# a_2477_543# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X35 a_481_107# a_30_107# a_637_569# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X36 VPWR a_935_107# a_1201_123# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X37 a_2477_543# a_1201_123# a_2656_543# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X38 a_2335_543# a_935_107# a_2477_543# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
X39 a_637_107# SCD VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__sdfxbp_1 CLK D SCD SCE VGND VNB VPB VPWR Q Q_N
X0 a_1528_579# a_1570_457# a_1124_81# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X1 a_425_107# SCE a_567_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X2 VGND a_2518_445# a_2789_147# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X3 a_2365_445# a_2789_147# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X4 VGND CLK a_1570_457# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X5 a_30_515# SCE VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X6 a_567_107# a_30_515# a_723_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X7 VPWR a_2789_147# a_3531_107# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X8 a_2518_445# a_1570_457# a_2747_173# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X9 a_268_659# a_30_515# a_567_107# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X10 VPWR CLK a_1570_457# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X11 a_567_107# a_1570_457# a_1124_81# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X12 VGND SCD a_425_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X13 a_567_107# D a_581_659# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X14 VGND a_1067_107# a_1454_173# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X15 VGND a_3531_107# Q_N VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X16 a_268_659# SCD VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X17 a_1067_107# a_1726_453# a_2518_445# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X18 a_1067_107# a_1124_81# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
X19 a_1124_81# a_1726_453# a_567_107# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X20 VPWR a_3531_107# Q_N VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X21 a_1726_453# a_1570_457# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X22 a_723_107# D VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X23 Q a_2789_147# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X24 a_1124_81# a_1726_453# a_1454_173# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X25 a_30_515# SCE VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X26 a_1067_107# a_1124_81# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X27 a_2747_173# a_2789_147# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X28 VGND a_2789_147# a_3531_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X29 VPWR a_2518_445# a_2789_147# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
X30 Q a_2789_147# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X31 a_2365_445# a_1726_453# a_2518_445# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X32 a_1726_453# a_1570_457# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X33 VPWR a_1067_107# a_1528_579# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X34 VPWR SCE a_581_659# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X35 a_2518_445# a_1570_457# a_1067_107# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__sdfxtp_1 CLK D SCD SCE VGND VNB VPB VPWR Q
X0 VPWR a_2123_543# a_2352_81# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
X1 VPWR CLK a_938_107# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X2 a_342_107# a_30_593# a_484_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X3 a_2123_543# a_938_107# a_2310_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X4 a_484_107# a_30_593# a_641_593# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X5 Q a_2352_81# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X6 a_1688_81# a_1204_107# a_2123_543# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X7 a_30_593# SCE VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X8 a_484_107# SCE a_640_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X9 a_1490_107# a_1204_107# a_1646_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X10 a_1490_107# a_938_107# a_1646_543# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X11 VPWR SCE a_343_593# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X12 a_2123_543# a_1204_107# a_2302_543# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X13 VGND a_938_107# a_1204_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X14 a_1688_81# a_938_107# a_2123_543# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
X15 a_30_593# SCE VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X16 VGND D a_342_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X17 VGND CLK a_938_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X18 a_484_107# a_938_107# a_1490_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X19 a_2310_107# a_2352_81# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X20 a_484_107# a_1204_107# a_1490_107# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X21 a_2302_543# a_2352_81# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X22 a_641_593# SCD VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X23 a_640_107# SCD VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X24 a_1646_107# a_1688_81# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X25 VGND a_1490_107# a_1688_81# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X26 VPWR a_1490_107# a_1688_81# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
X27 Q a_2352_81# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X28 a_1646_543# a_1688_81# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X29 a_343_593# D a_484_107# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X30 VPWR a_938_107# a_1204_107# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X31 VGND a_2123_543# a_2352_81# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__sdlclkp_1 CLK GATE SCE VGND VNB VPB VPWR GCLK
X0 VGND a_1630_171# GCLK VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X1 a_1783_171# CLK VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X2 a_58_159# a_423_71# a_495_311# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X3 VPWR a_1261_133# a_1630_171# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X4 VPWR SCE a_219_457# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X5 VPWR CLK a_423_71# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X6 VPWR a_1630_171# GCLK VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X7 a_431_431# a_423_71# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X8 VPWR a_495_311# a_1261_133# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X9 VGND CLK a_423_71# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X10 a_1630_171# a_1261_133# a_1783_171# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X11 a_58_159# SCE VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X12 a_219_457# GATE a_58_159# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X13 a_495_311# a_423_71# a_1219_457# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X14 a_1219_457# a_1261_133# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X15 VGND a_495_311# a_1261_133# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X16 a_58_159# a_431_431# a_495_311# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X17 a_1630_171# CLK VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X18 VGND GATE a_58_159# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X19 a_495_311# a_431_431# a_1219_159# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X20 a_431_431# a_423_71# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X21 a_1219_159# a_1261_133# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__sdlxtp_1 D GATE SCD SCE VGND VNB VPB VPWR Q
X0 a_1724_593# a_1678_81# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X1 a_1480_107# a_944_107# a_1636_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X2 a_489_107# SCE a_645_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X3 a_1678_81# a_1480_107# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X4 a_489_107# a_30_587# a_660_587# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X5 a_489_107# a_1214_107# a_1480_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X6 VGND D a_347_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X7 a_1480_107# a_1214_107# a_1724_593# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X8 VPWR a_944_107# a_1214_107# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X9 a_489_107# a_944_107# a_1480_107# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X10 VPWR SCE a_362_587# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X11 VPWR a_1480_107# Q VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X12 VPWR GATE a_944_107# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X13 a_1636_107# a_1678_81# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X14 VGND GATE a_944_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X15 VGND a_944_107# a_1214_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X16 a_660_587# SCD VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X17 a_645_107# SCD VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X18 a_30_587# SCE VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X19 a_30_587# SCE VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X20 a_347_107# a_30_587# a_489_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X21 a_1678_81# a_1480_107# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X22 VGND a_1480_107# Q VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X23 a_362_587# D a_489_107# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__xnor2_1 A B VGND VNB VPB VPWR Y
X0 VGND A a_523_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X1 VPWR A a_539_443# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X2 VPWR B a_30_107# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X3 a_539_443# B Y VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X4 a_222_107# A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X5 a_523_107# a_30_107# Y VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X6 a_523_107# B VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X7 Y a_30_107# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X8 a_30_107# B a_222_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X9 a_30_107# A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__xor2_1 A B VGND VNB VPB VPWR X
X0 X a_30_443# a_531_443# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X1 VGND B a_30_443# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X2 a_30_443# A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X3 a_30_443# B a_187_443# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X4 a_617_107# B X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X5 a_187_443# A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X6 a_531_443# B VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X7 X a_30_443# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X8 VPWR A a_531_443# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X9 VGND A a_617_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
.ends


******* EOF

