magic
tech sky130A
magscale 1 2
timestamp 1676037725
<< nwell >>
rect -38 261 2706 582
<< pwell >>
rect 1408 157 1759 201
rect 2198 157 2667 203
rect 1 21 2667 157
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 131
rect 151 47 181 131
rect 235 47 265 131
rect 319 47 349 131
rect 513 47 543 131
rect 701 47 731 131
rect 785 47 815 131
rect 973 47 1003 131
rect 1057 47 1087 131
rect 1129 47 1159 131
rect 1317 47 1347 131
rect 1389 47 1419 131
rect 1484 47 1514 175
rect 1653 47 1683 175
rect 1777 47 1807 131
rect 1849 47 1879 131
rect 1977 47 2007 131
rect 2088 47 2118 131
rect 2276 47 2306 177
rect 2464 47 2494 131
rect 2559 47 2589 177
<< scpmoshvt >>
rect 79 369 109 497
rect 163 369 193 497
rect 235 369 265 497
rect 319 369 349 497
rect 507 369 537 497
rect 695 369 725 497
rect 779 369 809 497
rect 967 413 997 497
rect 1051 413 1081 497
rect 1153 413 1183 497
rect 1271 413 1301 497
rect 1368 413 1398 497
rect 1484 329 1514 497
rect 1557 329 1587 497
rect 1682 413 1712 497
rect 1770 413 1800 497
rect 1899 413 1929 497
rect 2087 413 2117 497
rect 2276 297 2306 497
rect 2464 355 2494 483
rect 2559 297 2589 497
<< ndiff >>
rect 1434 131 1484 175
rect 27 103 79 131
rect 27 69 35 103
rect 69 69 79 103
rect 27 47 79 69
rect 109 47 151 131
rect 181 98 235 131
rect 181 64 191 98
rect 225 64 235 98
rect 181 47 235 64
rect 265 47 319 131
rect 349 93 407 131
rect 349 59 365 93
rect 399 59 407 93
rect 349 47 407 59
rect 461 105 513 131
rect 461 71 469 105
rect 503 71 513 105
rect 461 47 513 71
rect 543 93 595 131
rect 543 59 553 93
rect 587 59 595 93
rect 543 47 595 59
rect 649 105 701 131
rect 649 71 657 105
rect 691 71 701 105
rect 649 47 701 71
rect 731 89 785 131
rect 731 55 741 89
rect 775 55 785 89
rect 731 47 785 55
rect 815 101 867 131
rect 815 67 825 101
rect 859 67 867 101
rect 815 47 867 67
rect 921 101 973 131
rect 921 67 929 101
rect 963 67 973 101
rect 921 47 973 67
rect 1003 101 1057 131
rect 1003 67 1013 101
rect 1047 67 1057 101
rect 1003 47 1057 67
rect 1087 47 1129 131
rect 1159 93 1211 131
rect 1159 59 1169 93
rect 1203 59 1211 93
rect 1159 47 1211 59
rect 1265 119 1317 131
rect 1265 85 1273 119
rect 1307 85 1317 119
rect 1265 47 1317 85
rect 1347 47 1389 131
rect 1419 89 1484 131
rect 1419 55 1429 89
rect 1463 55 1484 89
rect 1419 47 1484 55
rect 1514 47 1653 175
rect 1683 131 1733 175
rect 2224 161 2276 177
rect 1683 89 1777 131
rect 1683 55 1698 89
rect 1732 55 1777 89
rect 1683 47 1777 55
rect 1807 47 1849 131
rect 1879 47 1977 131
rect 2007 89 2088 131
rect 2007 55 2044 89
rect 2078 55 2088 89
rect 2007 47 2088 55
rect 2118 101 2170 131
rect 2118 67 2128 101
rect 2162 67 2170 101
rect 2118 47 2170 67
rect 2224 127 2232 161
rect 2266 127 2276 161
rect 2224 93 2276 127
rect 2224 59 2232 93
rect 2266 59 2276 93
rect 2224 47 2276 59
rect 2306 161 2358 177
rect 2306 127 2316 161
rect 2350 127 2358 161
rect 2509 131 2559 177
rect 2306 93 2358 127
rect 2306 59 2316 93
rect 2350 59 2358 93
rect 2306 47 2358 59
rect 2412 105 2464 131
rect 2412 71 2420 105
rect 2454 71 2464 105
rect 2412 47 2464 71
rect 2494 103 2559 131
rect 2494 69 2515 103
rect 2549 69 2559 103
rect 2494 47 2559 69
rect 2589 165 2641 177
rect 2589 131 2599 165
rect 2633 131 2641 165
rect 2589 97 2641 131
rect 2589 63 2599 97
rect 2633 63 2641 97
rect 2589 47 2641 63
<< pdiff >>
rect 27 431 79 497
rect 27 397 35 431
rect 69 397 79 431
rect 27 369 79 397
rect 109 489 163 497
rect 109 455 119 489
rect 153 455 163 489
rect 109 369 163 455
rect 193 369 235 497
rect 265 411 319 497
rect 265 377 275 411
rect 309 377 319 411
rect 265 369 319 377
rect 349 485 401 497
rect 349 451 359 485
rect 393 451 401 485
rect 349 369 401 451
rect 455 415 507 497
rect 455 381 463 415
rect 497 381 507 415
rect 455 369 507 381
rect 537 485 589 497
rect 537 451 547 485
rect 581 451 589 485
rect 537 369 589 451
rect 643 449 695 497
rect 643 415 651 449
rect 685 415 695 449
rect 643 369 695 415
rect 725 489 779 497
rect 725 455 735 489
rect 769 455 779 489
rect 725 369 779 455
rect 809 477 861 497
rect 809 443 819 477
rect 853 443 861 477
rect 809 369 861 443
rect 915 477 967 497
rect 915 443 923 477
rect 957 443 967 477
rect 915 413 967 443
rect 997 477 1051 497
rect 997 443 1007 477
rect 1041 443 1051 477
rect 997 413 1051 443
rect 1081 413 1153 497
rect 1183 489 1271 497
rect 1183 455 1205 489
rect 1239 455 1271 489
rect 1183 413 1271 455
rect 1301 474 1368 497
rect 1301 440 1315 474
rect 1349 440 1368 474
rect 1301 413 1368 440
rect 1398 489 1484 497
rect 1398 455 1417 489
rect 1451 455 1484 489
rect 1398 413 1484 455
rect 1434 329 1484 413
rect 1514 329 1557 497
rect 1587 475 1682 497
rect 1587 441 1626 475
rect 1660 441 1682 475
rect 1587 413 1682 441
rect 1712 413 1770 497
rect 1800 489 1899 497
rect 1800 455 1855 489
rect 1889 455 1899 489
rect 1800 413 1899 455
rect 1929 474 1981 497
rect 1929 440 1939 474
rect 1973 440 1981 474
rect 1929 413 1981 440
rect 2035 485 2087 497
rect 2035 451 2043 485
rect 2077 451 2087 485
rect 2035 413 2087 451
rect 2117 474 2169 497
rect 2117 440 2127 474
rect 2161 440 2169 474
rect 2117 413 2169 440
rect 2224 485 2276 497
rect 2224 451 2232 485
rect 2266 451 2276 485
rect 2224 417 2276 451
rect 1587 329 1637 413
rect 2224 383 2232 417
rect 2266 383 2276 417
rect 2224 349 2276 383
rect 2224 315 2232 349
rect 2266 315 2276 349
rect 2224 297 2276 315
rect 2306 484 2358 497
rect 2306 450 2316 484
rect 2350 450 2358 484
rect 2509 483 2559 497
rect 2306 416 2358 450
rect 2306 382 2316 416
rect 2350 382 2358 416
rect 2306 348 2358 382
rect 2412 471 2464 483
rect 2412 437 2420 471
rect 2454 437 2464 471
rect 2412 403 2464 437
rect 2412 369 2420 403
rect 2454 369 2464 403
rect 2412 355 2464 369
rect 2494 465 2559 483
rect 2494 431 2515 465
rect 2549 431 2559 465
rect 2494 397 2559 431
rect 2494 363 2515 397
rect 2549 363 2559 397
rect 2494 355 2559 363
rect 2306 314 2316 348
rect 2350 314 2358 348
rect 2306 297 2358 314
rect 2509 297 2559 355
rect 2589 485 2641 497
rect 2589 451 2599 485
rect 2633 451 2641 485
rect 2589 417 2641 451
rect 2589 383 2599 417
rect 2633 383 2641 417
rect 2589 349 2641 383
rect 2589 315 2599 349
rect 2633 315 2641 349
rect 2589 297 2641 315
<< ndiffc >>
rect 35 69 69 103
rect 191 64 225 98
rect 365 59 399 93
rect 469 71 503 105
rect 553 59 587 93
rect 657 71 691 105
rect 741 55 775 89
rect 825 67 859 101
rect 929 67 963 101
rect 1013 67 1047 101
rect 1169 59 1203 93
rect 1273 85 1307 119
rect 1429 55 1463 89
rect 1698 55 1732 89
rect 2044 55 2078 89
rect 2128 67 2162 101
rect 2232 127 2266 161
rect 2232 59 2266 93
rect 2316 127 2350 161
rect 2316 59 2350 93
rect 2420 71 2454 105
rect 2515 69 2549 103
rect 2599 131 2633 165
rect 2599 63 2633 97
<< pdiffc >>
rect 35 397 69 431
rect 119 455 153 489
rect 275 377 309 411
rect 359 451 393 485
rect 463 381 497 415
rect 547 451 581 485
rect 651 415 685 449
rect 735 455 769 489
rect 819 443 853 477
rect 923 443 957 477
rect 1007 443 1041 477
rect 1205 455 1239 489
rect 1315 440 1349 474
rect 1417 455 1451 489
rect 1626 441 1660 475
rect 1855 455 1889 489
rect 1939 440 1973 474
rect 2043 451 2077 485
rect 2127 440 2161 474
rect 2232 451 2266 485
rect 2232 383 2266 417
rect 2232 315 2266 349
rect 2316 450 2350 484
rect 2316 382 2350 416
rect 2420 437 2454 471
rect 2420 369 2454 403
rect 2515 431 2549 465
rect 2515 363 2549 397
rect 2316 314 2350 348
rect 2599 451 2633 485
rect 2599 383 2633 417
rect 2599 315 2633 349
<< poly >>
rect 79 497 109 523
rect 163 497 193 523
rect 235 497 265 523
rect 319 497 349 523
rect 507 497 537 523
rect 695 497 725 523
rect 779 497 809 523
rect 967 497 997 523
rect 1051 497 1081 523
rect 1153 497 1183 523
rect 1271 497 1301 523
rect 1368 497 1398 523
rect 1484 497 1514 523
rect 1557 497 1587 523
rect 1682 497 1712 523
rect 1770 497 1800 523
rect 1899 497 1929 523
rect 2087 497 2117 523
rect 2276 497 2306 523
rect 967 398 997 413
rect 79 354 109 369
rect 49 324 109 354
rect 49 265 79 324
rect 163 283 193 369
rect 22 249 79 265
rect 22 215 35 249
rect 69 215 79 249
rect 121 267 193 283
rect 121 233 131 267
rect 165 253 193 267
rect 165 233 181 253
rect 121 217 181 233
rect 235 219 265 369
rect 319 265 349 369
rect 507 265 537 369
rect 695 354 725 369
rect 683 324 725 354
rect 683 284 713 324
rect 779 284 809 369
rect 908 368 997 398
rect 1051 381 1081 413
rect 1153 381 1183 413
rect 908 284 938 368
rect 1039 365 1093 381
rect 1039 331 1049 365
rect 1083 331 1093 365
rect 1039 315 1093 331
rect 1153 365 1229 381
rect 1153 331 1185 365
rect 1219 331 1229 365
rect 1153 315 1229 331
rect 659 268 713 284
rect 319 249 429 265
rect 22 199 79 215
rect 49 176 79 199
rect 49 146 109 176
rect 79 131 109 146
rect 151 131 181 217
rect 223 203 277 219
rect 223 169 233 203
rect 267 169 277 203
rect 223 153 277 169
rect 319 215 373 249
rect 407 215 429 249
rect 319 199 429 215
rect 480 249 543 265
rect 480 215 490 249
rect 524 215 543 249
rect 659 234 669 268
rect 703 234 713 268
rect 659 218 713 234
rect 755 268 812 284
rect 755 234 765 268
rect 799 234 812 268
rect 755 218 812 234
rect 854 268 938 284
rect 854 234 864 268
rect 898 248 938 268
rect 898 234 1087 248
rect 854 218 1087 234
rect 480 199 543 215
rect 235 131 265 153
rect 319 131 349 199
rect 513 131 543 199
rect 683 176 713 218
rect 782 176 812 218
rect 683 146 731 176
rect 782 146 1003 176
rect 701 131 731 146
rect 785 131 815 146
rect 973 131 1003 146
rect 1057 131 1087 218
rect 1153 213 1183 315
rect 1271 273 1301 413
rect 1368 369 1398 413
rect 1343 353 1398 369
rect 1343 319 1353 353
rect 1387 319 1398 353
rect 1682 381 1712 413
rect 1674 365 1728 381
rect 1674 345 1684 365
rect 1653 331 1684 345
rect 1718 331 1728 365
rect 1343 303 1398 319
rect 1237 270 1301 273
rect 1368 273 1398 303
rect 1237 263 1303 270
rect 1237 229 1253 263
rect 1287 229 1303 263
rect 1368 243 1419 273
rect 1484 265 1514 329
rect 1557 265 1587 329
rect 1653 315 1728 331
rect 1770 325 1800 413
rect 1899 397 1929 413
rect 1899 367 2007 397
rect 2087 375 2117 413
rect 1953 339 2007 367
rect 1237 219 1303 229
rect 1129 203 1195 213
rect 1129 169 1145 203
rect 1179 169 1195 203
rect 1129 159 1195 169
rect 1273 176 1303 219
rect 1129 131 1159 159
rect 1273 146 1347 176
rect 1317 131 1347 146
rect 1389 131 1419 243
rect 1461 249 1515 265
rect 1461 215 1471 249
rect 1505 215 1515 249
rect 1461 199 1515 215
rect 1557 249 1611 265
rect 1557 215 1567 249
rect 1601 215 1611 249
rect 1557 199 1611 215
rect 1484 175 1514 199
rect 1653 175 1683 315
rect 1770 295 1879 325
rect 1752 233 1807 249
rect 1752 199 1763 233
rect 1797 199 1807 233
rect 1752 183 1807 199
rect 1777 131 1807 183
rect 1849 237 1879 295
rect 1953 305 1963 339
rect 1997 305 2007 339
rect 1953 289 2007 305
rect 1849 221 1903 237
rect 1849 187 1859 221
rect 1893 187 1903 221
rect 1849 171 1903 187
rect 1849 131 1879 171
rect 1977 131 2007 289
rect 2049 355 2117 375
rect 2049 321 2059 355
rect 2093 321 2117 355
rect 2049 265 2117 321
rect 2464 483 2494 523
rect 2559 497 2589 523
rect 2276 265 2306 297
rect 2464 265 2494 355
rect 2559 265 2589 297
rect 2049 203 2494 265
rect 2049 169 2059 203
rect 2093 199 2494 203
rect 2536 249 2590 265
rect 2536 215 2546 249
rect 2580 215 2590 249
rect 2536 199 2590 215
rect 2093 169 2118 199
rect 2276 177 2306 199
rect 2049 153 2118 169
rect 2088 131 2118 153
rect 2464 131 2494 199
rect 2559 177 2589 199
rect 79 21 109 47
rect 151 21 181 47
rect 235 21 265 47
rect 319 21 349 47
rect 513 21 543 47
rect 701 21 731 47
rect 785 21 815 47
rect 973 21 1003 47
rect 1057 21 1087 47
rect 1129 21 1159 47
rect 1317 21 1347 47
rect 1389 21 1419 47
rect 1484 21 1514 47
rect 1653 21 1683 47
rect 1777 21 1807 47
rect 1849 21 1879 47
rect 1977 21 2007 47
rect 2088 21 2118 47
rect 2276 21 2306 47
rect 2464 21 2494 47
rect 2559 21 2589 47
<< polycont >>
rect 35 215 69 249
rect 131 233 165 267
rect 1049 331 1083 365
rect 1185 331 1219 365
rect 233 169 267 203
rect 373 215 407 249
rect 490 215 524 249
rect 669 234 703 268
rect 765 234 799 268
rect 864 234 898 268
rect 1353 319 1387 353
rect 1684 331 1718 365
rect 1253 229 1287 263
rect 1145 169 1179 203
rect 1471 215 1505 249
rect 1567 215 1601 249
rect 1763 199 1797 233
rect 1963 305 1997 339
rect 1859 187 1893 221
rect 2059 321 2093 355
rect 2059 169 2093 203
rect 2546 215 2580 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2668 561
rect 17 431 69 493
rect 103 489 153 527
rect 103 455 119 489
rect 103 439 153 455
rect 187 485 409 493
rect 187 451 359 485
rect 393 451 409 485
rect 17 397 35 431
rect 187 405 221 451
rect 454 417 504 493
rect 538 485 606 527
rect 538 451 547 485
rect 581 451 606 485
rect 719 489 785 527
rect 538 428 606 451
rect 651 449 685 465
rect 719 455 735 489
rect 769 455 785 489
rect 819 477 888 493
rect 373 415 504 417
rect 69 397 221 405
rect 17 369 221 397
rect 259 411 339 415
rect 259 377 275 411
rect 309 377 339 411
rect 259 374 339 377
rect 17 249 69 335
rect 17 215 35 249
rect 17 153 69 215
rect 109 267 165 335
rect 109 255 131 267
rect 109 221 122 255
rect 156 221 165 233
rect 109 153 165 221
rect 211 203 267 335
rect 211 169 233 203
rect 211 153 267 169
rect 301 323 339 374
rect 301 289 305 323
rect 301 141 339 289
rect 373 381 463 415
rect 497 381 504 415
rect 853 443 888 477
rect 819 427 888 443
rect 373 354 504 381
rect 373 249 440 354
rect 407 215 440 249
rect 474 255 540 320
rect 474 221 489 255
rect 523 249 540 255
rect 474 215 490 221
rect 524 215 540 249
rect 581 318 617 392
rect 651 391 685 415
rect 651 357 765 391
rect 651 355 799 357
rect 581 268 713 318
rect 581 234 669 268
rect 703 234 713 268
rect 373 181 440 215
rect 581 211 713 234
rect 747 268 799 355
rect 747 234 765 268
rect 373 143 503 181
rect 581 145 620 211
rect 747 177 799 234
rect 299 133 339 141
rect 295 131 339 133
rect 295 129 334 131
rect 292 127 334 129
rect 289 126 334 127
rect 288 124 334 126
rect 286 123 334 124
rect 284 122 332 123
rect 281 121 332 122
rect 279 120 332 121
rect 17 103 96 119
rect 276 118 332 120
rect 276 112 331 118
rect 17 69 35 103
rect 69 69 96 103
rect 17 17 96 69
rect 175 98 331 112
rect 175 64 191 98
rect 225 64 331 98
rect 175 56 331 64
rect 365 93 401 109
rect 399 59 401 93
rect 365 17 401 59
rect 452 105 503 143
rect 654 143 799 177
rect 833 284 888 427
rect 922 477 966 493
rect 922 443 923 477
rect 957 443 966 477
rect 922 323 966 443
rect 1006 477 1151 493
rect 1006 443 1007 477
rect 1041 443 1151 477
rect 1189 489 1255 527
rect 1189 455 1205 489
rect 1239 455 1255 489
rect 1310 474 1353 490
rect 1006 427 1151 443
rect 1075 365 1083 391
rect 1041 331 1049 357
rect 922 318 949 323
rect 932 289 949 318
rect 1041 315 1083 331
rect 833 268 898 284
rect 833 255 864 268
rect 833 221 857 255
rect 891 221 898 234
rect 833 218 898 221
rect 452 71 469 105
rect 452 51 503 71
rect 538 93 606 111
rect 538 59 553 93
rect 587 59 606 93
rect 538 17 606 59
rect 654 105 691 143
rect 833 117 867 218
rect 932 184 966 289
rect 1117 279 1151 427
rect 1310 440 1315 474
rect 1349 440 1353 474
rect 1310 421 1353 440
rect 1401 489 1592 527
rect 1401 455 1417 489
rect 1451 455 1592 489
rect 1401 425 1592 455
rect 1626 475 1787 492
rect 1660 441 1787 475
rect 1839 489 1905 527
rect 1839 455 1855 489
rect 1889 455 1905 489
rect 1839 447 1905 455
rect 1939 474 1982 490
rect 1626 425 1787 441
rect 1185 387 1353 421
rect 1753 413 1787 425
rect 1973 440 1982 474
rect 2027 485 2093 527
rect 2027 451 2043 485
rect 2077 451 2093 485
rect 2027 447 2093 451
rect 2127 474 2179 493
rect 1939 413 1982 440
rect 2161 440 2179 474
rect 1185 365 1219 387
rect 1438 357 1501 391
rect 1535 357 1601 391
rect 1185 315 1219 331
rect 1328 323 1353 353
rect 1387 319 1403 353
rect 1362 289 1403 319
rect 1438 299 1601 357
rect 1017 263 1287 279
rect 1017 255 1253 263
rect 654 71 657 105
rect 654 51 691 71
rect 726 89 788 109
rect 726 55 741 89
rect 775 55 788 89
rect 726 17 788 55
rect 822 101 867 117
rect 822 67 825 101
rect 859 67 867 101
rect 822 51 867 67
rect 901 101 966 184
rect 901 67 929 101
rect 963 67 966 101
rect 901 51 966 67
rect 1000 245 1253 255
rect 1000 101 1088 245
rect 1250 229 1253 245
rect 1460 255 1532 265
rect 1287 249 1532 255
rect 1287 229 1471 249
rect 1250 215 1471 229
rect 1505 215 1532 249
rect 1122 169 1145 203
rect 1179 169 1195 203
rect 1250 195 1532 215
rect 1567 249 1601 299
rect 1673 365 1719 381
rect 1753 379 2093 413
rect 1673 331 1684 365
rect 1718 331 1719 365
rect 2049 355 2093 379
rect 1673 255 1719 331
rect 1777 339 2015 345
rect 1777 323 1963 339
rect 1811 305 1963 323
rect 1997 305 2015 339
rect 2049 321 2059 355
rect 2049 305 2093 321
rect 1811 289 1822 305
rect 1777 283 1822 289
rect 2127 271 2179 440
rect 2224 485 2266 527
rect 2224 451 2232 485
rect 2224 417 2266 451
rect 2224 383 2232 417
rect 2224 349 2266 383
rect 2224 315 2232 349
rect 2224 297 2266 315
rect 2300 484 2366 493
rect 2300 450 2316 484
rect 2350 450 2366 484
rect 2300 416 2366 450
rect 2300 382 2316 416
rect 2350 382 2366 416
rect 2300 348 2366 382
rect 2300 314 2316 348
rect 2350 314 2366 348
rect 1673 221 1685 255
rect 1673 215 1719 221
rect 1762 233 1808 249
rect 1122 161 1195 169
rect 1567 179 1601 215
rect 1762 199 1763 233
rect 1797 199 1808 233
rect 1762 179 1808 199
rect 1122 127 1307 161
rect 1000 67 1013 101
rect 1047 67 1088 101
rect 1255 119 1307 127
rect 1000 51 1088 67
rect 1122 59 1169 93
rect 1203 59 1219 93
rect 1122 17 1219 59
rect 1255 85 1273 119
rect 1255 51 1307 85
rect 1347 89 1526 161
rect 1567 139 1808 179
rect 1858 237 2179 271
rect 1858 221 1893 237
rect 1858 187 1859 221
rect 1858 171 1893 187
rect 1931 169 2059 203
rect 2093 169 2109 203
rect 1931 89 1965 169
rect 1347 55 1429 89
rect 1463 55 1526 89
rect 1682 55 1698 89
rect 1732 55 1965 89
rect 2044 89 2078 109
rect 2143 108 2179 237
rect 1347 17 1526 55
rect 2044 17 2078 55
rect 2112 101 2179 108
rect 2112 67 2128 101
rect 2162 67 2179 101
rect 2112 51 2179 67
rect 2224 161 2266 177
rect 2224 127 2232 161
rect 2224 93 2266 127
rect 2224 59 2232 93
rect 2224 17 2266 59
rect 2300 161 2366 314
rect 2300 127 2316 161
rect 2350 127 2366 161
rect 2300 93 2366 127
rect 2300 59 2316 93
rect 2350 59 2366 93
rect 2300 51 2366 59
rect 2412 471 2454 493
rect 2412 437 2420 471
rect 2412 403 2454 437
rect 2412 369 2420 403
rect 2412 265 2454 369
rect 2515 465 2549 527
rect 2515 397 2549 431
rect 2515 315 2549 363
rect 2583 485 2651 490
rect 2583 451 2599 485
rect 2633 451 2651 485
rect 2583 417 2651 451
rect 2583 383 2599 417
rect 2633 383 2651 417
rect 2583 349 2651 383
rect 2583 315 2599 349
rect 2633 315 2651 349
rect 2583 299 2651 315
rect 2412 249 2580 265
rect 2412 215 2546 249
rect 2412 199 2580 215
rect 2412 105 2454 199
rect 2614 165 2651 299
rect 2412 71 2420 105
rect 2412 51 2454 71
rect 2508 103 2549 165
rect 2508 69 2515 103
rect 2508 17 2549 69
rect 2583 131 2599 165
rect 2633 131 2651 165
rect 2583 97 2651 131
rect 2583 63 2599 97
rect 2633 63 2651 97
rect 2583 55 2651 63
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2668 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 2237 527 2271 561
rect 2329 527 2363 561
rect 2421 527 2455 561
rect 2513 527 2547 561
rect 2605 527 2639 561
rect 122 233 131 255
rect 131 233 156 255
rect 122 221 156 233
rect 305 289 339 323
rect 489 249 523 255
rect 489 221 490 249
rect 490 221 523 249
rect 765 357 799 391
rect 1041 365 1075 391
rect 1041 357 1049 365
rect 1049 357 1075 365
rect 949 289 983 323
rect 857 234 864 255
rect 864 234 891 255
rect 857 221 891 234
rect 1501 357 1535 391
rect 1328 319 1353 323
rect 1353 319 1362 323
rect 1328 289 1362 319
rect 1777 289 1811 323
rect 1685 221 1719 255
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
rect 2329 -17 2363 17
rect 2421 -17 2455 17
rect 2513 -17 2547 17
rect 2605 -17 2639 17
<< metal1 >>
rect 0 561 2668 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2668 561
rect 0 496 2668 527
rect 753 391 811 397
rect 753 357 765 391
rect 799 388 811 391
rect 1029 391 1087 397
rect 1029 388 1041 391
rect 799 360 1041 388
rect 799 357 811 360
rect 753 351 811 357
rect 1029 357 1041 360
rect 1075 388 1087 391
rect 1489 391 1547 397
rect 1489 388 1501 391
rect 1075 360 1501 388
rect 1075 357 1087 360
rect 1029 351 1087 357
rect 1489 357 1501 360
rect 1535 357 1547 391
rect 1489 351 1547 357
rect 293 323 351 329
rect 293 289 305 323
rect 339 320 351 323
rect 937 323 995 329
rect 937 320 949 323
rect 339 292 949 320
rect 339 289 351 292
rect 293 283 351 289
rect 937 289 949 292
rect 983 289 995 323
rect 937 283 995 289
rect 1316 323 1374 329
rect 1316 289 1328 323
rect 1362 320 1374 323
rect 1765 323 1823 329
rect 1765 320 1777 323
rect 1362 292 1777 320
rect 1362 289 1374 292
rect 1316 283 1374 289
rect 1765 289 1777 292
rect 1811 289 1823 323
rect 1765 283 1823 289
rect 110 255 168 261
rect 110 221 122 255
rect 156 252 168 255
rect 477 255 535 261
rect 477 252 489 255
rect 156 224 489 252
rect 156 221 168 224
rect 110 215 168 221
rect 477 221 489 224
rect 523 221 535 255
rect 477 215 535 221
rect 845 255 903 261
rect 845 221 857 255
rect 891 252 903 255
rect 1673 255 1731 261
rect 1673 252 1685 255
rect 891 224 1685 252
rect 891 221 903 224
rect 845 215 903 221
rect 1673 221 1685 224
rect 1719 221 1731 255
rect 1673 215 1731 221
rect 0 17 2668 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2668 17
rect 0 -48 2668 -17
<< labels >>
flabel locali s 30 153 64 187 0 FreeSans 200 0 0 0 SCD
port 3 nsew signal input
flabel locali s 581 357 615 391 0 FreeSans 200 0 0 0 CLK
port 1 nsew clock input
flabel locali s 2329 357 2363 391 0 FreeSans 200 0 0 0 Q_N
port 11 nsew signal output
flabel locali s 214 289 248 323 0 FreeSans 200 0 0 0 D
port 2 nsew signal input
flabel locali s 2329 425 2363 459 0 FreeSans 200 0 0 0 Q_N
port 11 nsew signal output
flabel locali s 30 289 64 323 0 FreeSans 200 0 0 0 SCD
port 3 nsew signal input
flabel locali s 2329 289 2363 323 0 FreeSans 200 0 0 0 Q_N
port 11 nsew signal output
flabel locali s 2329 221 2363 255 0 FreeSans 200 0 0 0 Q_N
port 11 nsew signal output
flabel locali s 2329 153 2363 187 0 FreeSans 200 0 0 0 Q_N
port 11 nsew signal output
flabel locali s 2329 85 2363 119 0 FreeSans 200 0 0 0 Q_N
port 11 nsew signal output
flabel locali s 1328 289 1362 323 0 FreeSans 200 0 0 0 SET_B
port 5 nsew signal input
flabel locali s 122 221 156 255 0 FreeSans 200 0 0 0 SCE
port 4 nsew signal input
flabel locali s 214 153 248 187 0 FreeSans 200 0 0 0 D
port 2 nsew signal input
flabel locali s 581 221 615 255 0 FreeSans 200 0 0 0 CLK
port 1 nsew clock input
flabel locali s 581 153 615 187 0 FreeSans 200 0 0 0 CLK
port 1 nsew clock input
flabel locali s 673 221 707 255 0 FreeSans 200 0 0 0 CLK
port 1 nsew clock input
flabel locali s 2614 357 2648 391 0 FreeSans 200 0 0 0 Q
port 10 nsew signal output
flabel locali s 2614 425 2648 459 0 FreeSans 200 0 0 0 Q
port 10 nsew signal output
flabel locali s 2614 221 2648 255 0 FreeSans 200 0 0 0 Q
port 10 nsew signal output
flabel locali s 2614 153 2648 187 0 FreeSans 200 0 0 0 Q
port 10 nsew signal output
flabel locali s 2614 85 2648 119 0 FreeSans 200 0 0 0 Q
port 10 nsew signal output
flabel locali s 2614 289 2648 323 0 FreeSans 200 0 0 0 Q
port 10 nsew signal output
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 9 nsew power bidirectional abutment
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 6 nsew ground bidirectional abutment
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel comment s 2092 225 2092 225 0 FreeSans 200 0 0 0 no_jumper_check
rlabel comment s 0 0 0 0 4 sdfsbp_1
flabel comment s 1165 297 1165 297 0 FreeSans 200 0 0 0 no_jumper_check
rlabel locali s 474 215 540 320 1 SCE
port 4 nsew signal input
rlabel metal1 s 477 252 535 261 1 SCE
port 4 nsew signal input
rlabel metal1 s 477 215 535 224 1 SCE
port 4 nsew signal input
rlabel metal1 s 110 252 168 261 1 SCE
port 4 nsew signal input
rlabel metal1 s 110 224 535 252 1 SCE
port 4 nsew signal input
rlabel metal1 s 110 215 168 224 1 SCE
port 4 nsew signal input
rlabel locali s 1777 305 2015 345 1 SET_B
port 5 nsew signal input
rlabel locali s 1777 283 1822 305 1 SET_B
port 5 nsew signal input
rlabel metal1 s 1765 320 1823 329 1 SET_B
port 5 nsew signal input
rlabel metal1 s 1765 283 1823 292 1 SET_B
port 5 nsew signal input
rlabel metal1 s 1316 320 1374 329 1 SET_B
port 5 nsew signal input
rlabel metal1 s 1316 292 1823 320 1 SET_B
port 5 nsew signal input
rlabel metal1 s 1316 283 1374 292 1 SET_B
port 5 nsew signal input
rlabel metal1 s 0 -48 2668 48 1 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 496 2668 592 1 VPWR
port 9 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 2668 544
string GDS_END 53504
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 31832
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 2.720 13.340 2.720 
<< end >>
