magic
tech sky130B
magscale 1 2
timestamp 1676037725
<< locali >>
rect 243 1369 559 1388
rect 243 1335 255 1369
rect 289 1335 337 1369
rect 371 1335 431 1369
rect 465 1335 513 1369
rect 547 1335 559 1369
rect 243 1297 559 1335
rect 243 1263 255 1297
rect 289 1263 337 1297
rect 371 1263 431 1297
rect 465 1263 513 1297
rect 547 1263 559 1297
rect 243 1249 559 1263
rect 243 125 559 139
rect 243 91 255 125
rect 289 91 337 125
rect 371 91 431 125
rect 465 91 513 125
rect 547 91 559 125
rect 243 53 559 91
rect 243 19 255 53
rect 289 19 337 53
rect 371 19 431 53
rect 465 19 513 53
rect 547 19 559 53
rect 243 0 559 19
<< viali >>
rect 255 1335 289 1369
rect 337 1335 371 1369
rect 431 1335 465 1369
rect 513 1335 547 1369
rect 255 1263 289 1297
rect 337 1263 371 1297
rect 431 1263 465 1297
rect 513 1263 547 1297
rect 255 91 289 125
rect 337 91 371 125
rect 431 91 465 125
rect 513 91 547 125
rect 255 19 289 53
rect 337 19 371 53
rect 431 19 465 53
rect 513 19 547 53
<< obsli1 >>
rect 120 1231 186 1297
rect 616 1231 682 1297
rect 120 1203 160 1231
rect 642 1203 682 1231
rect 41 1179 160 1203
rect 41 1145 60 1179
rect 94 1145 160 1179
rect 41 1107 160 1145
rect 41 1073 60 1107
rect 94 1073 160 1107
rect 41 1035 160 1073
rect 41 1001 60 1035
rect 94 1001 160 1035
rect 41 963 160 1001
rect 41 929 60 963
rect 94 929 160 963
rect 41 891 160 929
rect 41 857 60 891
rect 94 857 160 891
rect 41 819 160 857
rect 41 785 60 819
rect 94 785 160 819
rect 41 747 160 785
rect 41 713 60 747
rect 94 713 160 747
rect 41 675 160 713
rect 41 641 60 675
rect 94 641 160 675
rect 41 603 160 641
rect 41 569 60 603
rect 94 569 160 603
rect 41 531 160 569
rect 41 497 60 531
rect 94 497 160 531
rect 41 459 160 497
rect 41 425 60 459
rect 94 425 160 459
rect 41 387 160 425
rect 41 353 60 387
rect 94 353 160 387
rect 41 315 160 353
rect 41 281 60 315
rect 94 281 160 315
rect 41 243 160 281
rect 41 209 60 243
rect 94 209 160 243
rect 41 185 160 209
rect 212 185 246 1203
rect 298 185 332 1203
rect 384 185 418 1203
rect 470 185 504 1203
rect 556 185 590 1203
rect 642 1179 761 1203
rect 642 1145 708 1179
rect 742 1145 761 1179
rect 642 1107 761 1145
rect 642 1073 708 1107
rect 742 1073 761 1107
rect 642 1035 761 1073
rect 642 1001 708 1035
rect 742 1001 761 1035
rect 642 963 761 1001
rect 642 929 708 963
rect 742 929 761 963
rect 642 891 761 929
rect 642 857 708 891
rect 742 857 761 891
rect 642 819 761 857
rect 642 785 708 819
rect 742 785 761 819
rect 642 747 761 785
rect 642 713 708 747
rect 742 713 761 747
rect 642 675 761 713
rect 642 641 708 675
rect 742 641 761 675
rect 642 603 761 641
rect 642 569 708 603
rect 742 569 761 603
rect 642 531 761 569
rect 642 497 708 531
rect 742 497 761 531
rect 642 459 761 497
rect 642 425 708 459
rect 742 425 761 459
rect 642 387 761 425
rect 642 353 708 387
rect 742 353 761 387
rect 642 315 761 353
rect 642 281 708 315
rect 742 281 761 315
rect 642 243 761 281
rect 642 209 708 243
rect 742 209 761 243
rect 642 185 761 209
rect 120 157 160 185
rect 642 157 682 185
rect 120 91 186 157
rect 616 91 682 157
<< obsli1c >>
rect 60 1145 94 1179
rect 60 1073 94 1107
rect 60 1001 94 1035
rect 60 929 94 963
rect 60 857 94 891
rect 60 785 94 819
rect 60 713 94 747
rect 60 641 94 675
rect 60 569 94 603
rect 60 497 94 531
rect 60 425 94 459
rect 60 353 94 387
rect 60 281 94 315
rect 60 209 94 243
rect 708 1145 742 1179
rect 708 1073 742 1107
rect 708 1001 742 1035
rect 708 929 742 963
rect 708 857 742 891
rect 708 785 742 819
rect 708 713 742 747
rect 708 641 742 675
rect 708 569 742 603
rect 708 497 742 531
rect 708 425 742 459
rect 708 353 742 387
rect 708 281 742 315
rect 708 209 742 243
<< metal1 >>
rect 243 1369 559 1388
rect 243 1335 255 1369
rect 289 1335 337 1369
rect 371 1335 431 1369
rect 465 1335 513 1369
rect 547 1335 559 1369
rect 243 1297 559 1335
rect 243 1263 255 1297
rect 289 1263 337 1297
rect 371 1263 431 1297
rect 465 1263 513 1297
rect 547 1263 559 1297
rect 243 1251 559 1263
rect 41 1179 100 1191
rect 41 1145 60 1179
rect 94 1145 100 1179
rect 41 1107 100 1145
rect 41 1073 60 1107
rect 94 1073 100 1107
rect 41 1035 100 1073
rect 41 1001 60 1035
rect 94 1001 100 1035
rect 41 963 100 1001
rect 41 929 60 963
rect 94 929 100 963
rect 41 891 100 929
rect 41 857 60 891
rect 94 857 100 891
rect 41 819 100 857
rect 41 785 60 819
rect 94 785 100 819
rect 41 747 100 785
rect 41 713 60 747
rect 94 713 100 747
rect 41 675 100 713
rect 41 641 60 675
rect 94 641 100 675
rect 41 603 100 641
rect 41 569 60 603
rect 94 569 100 603
rect 41 531 100 569
rect 41 497 60 531
rect 94 497 100 531
rect 41 459 100 497
rect 41 425 60 459
rect 94 425 100 459
rect 41 387 100 425
rect 41 353 60 387
rect 94 353 100 387
rect 41 315 100 353
rect 41 281 60 315
rect 94 281 100 315
rect 41 243 100 281
rect 41 209 60 243
rect 94 209 100 243
rect 41 197 100 209
rect 702 1179 761 1191
rect 702 1145 708 1179
rect 742 1145 761 1179
rect 702 1107 761 1145
rect 702 1073 708 1107
rect 742 1073 761 1107
rect 702 1035 761 1073
rect 702 1001 708 1035
rect 742 1001 761 1035
rect 702 963 761 1001
rect 702 929 708 963
rect 742 929 761 963
rect 702 891 761 929
rect 702 857 708 891
rect 742 857 761 891
rect 702 819 761 857
rect 702 785 708 819
rect 742 785 761 819
rect 702 747 761 785
rect 702 713 708 747
rect 742 713 761 747
rect 702 675 761 713
rect 702 641 708 675
rect 742 641 761 675
rect 702 603 761 641
rect 702 569 708 603
rect 742 569 761 603
rect 702 531 761 569
rect 702 497 708 531
rect 742 497 761 531
rect 702 459 761 497
rect 702 425 708 459
rect 742 425 761 459
rect 702 387 761 425
rect 702 353 708 387
rect 742 353 761 387
rect 702 315 761 353
rect 702 281 708 315
rect 742 281 761 315
rect 702 243 761 281
rect 702 209 708 243
rect 742 209 761 243
rect 702 197 761 209
rect 243 125 559 137
rect 243 91 255 125
rect 289 91 337 125
rect 371 91 431 125
rect 465 91 513 125
rect 547 91 559 125
rect 243 53 559 91
rect 243 19 255 53
rect 289 19 337 53
rect 371 19 431 53
rect 465 19 513 53
rect 547 19 559 53
rect 243 0 559 19
<< obsm1 >>
rect 203 197 255 1191
rect 289 197 341 1191
rect 375 197 427 1191
rect 461 197 513 1191
rect 547 197 599 1191
<< metal2 >>
rect 14 719 788 1191
rect 14 197 788 669
<< labels >>
rlabel metal1 s 702 197 761 1191 6 BULK
port 4 nsew
rlabel metal1 s 41 197 100 1191 6 BULK
port 4 nsew
rlabel metal2 s 14 719 788 1191 6 DRAIN
port 1 nsew
rlabel viali s 513 1335 547 1369 6 GATE
port 2 nsew
rlabel viali s 513 1263 547 1297 6 GATE
port 2 nsew
rlabel viali s 513 91 547 125 6 GATE
port 2 nsew
rlabel viali s 513 19 547 53 6 GATE
port 2 nsew
rlabel viali s 431 1335 465 1369 6 GATE
port 2 nsew
rlabel viali s 431 1263 465 1297 6 GATE
port 2 nsew
rlabel viali s 431 91 465 125 6 GATE
port 2 nsew
rlabel viali s 431 19 465 53 6 GATE
port 2 nsew
rlabel viali s 337 1335 371 1369 6 GATE
port 2 nsew
rlabel viali s 337 1263 371 1297 6 GATE
port 2 nsew
rlabel viali s 337 91 371 125 6 GATE
port 2 nsew
rlabel viali s 337 19 371 53 6 GATE
port 2 nsew
rlabel viali s 255 1335 289 1369 6 GATE
port 2 nsew
rlabel viali s 255 1263 289 1297 6 GATE
port 2 nsew
rlabel viali s 255 91 289 125 6 GATE
port 2 nsew
rlabel viali s 255 19 289 53 6 GATE
port 2 nsew
rlabel locali s 243 1249 559 1388 6 GATE
port 2 nsew
rlabel locali s 243 0 559 139 6 GATE
port 2 nsew
rlabel metal1 s 243 1251 559 1388 6 GATE
port 2 nsew
rlabel metal1 s 243 0 559 137 6 GATE
port 2 nsew
rlabel metal2 s 14 197 788 669 6 SOURCE
port 3 nsew
<< properties >>
string FIXED_BBOX 0 0 802 1388
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 9817484
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 9789886
string device primitive
<< end >>