magic
tech sky130A
magscale 1 2
timestamp 1676037725
<< locali >>
rect 161 1160 173 1194
rect 207 1160 245 1194
rect 279 1160 317 1194
rect 351 1160 363 1194
rect 48 1020 82 1058
rect 48 948 82 986
rect 48 876 82 914
rect 48 804 82 842
rect 48 732 82 770
rect 48 660 82 698
rect 48 588 82 626
rect 48 516 82 554
rect 48 444 82 482
rect 48 372 82 410
rect 48 300 82 338
rect 48 228 82 266
rect 48 122 82 194
rect 442 1020 476 1058
rect 442 948 476 986
rect 442 876 476 914
rect 442 804 476 842
rect 442 732 476 770
rect 442 660 476 698
rect 442 588 476 626
rect 442 516 476 554
rect 442 444 476 482
rect 442 372 476 410
rect 442 300 476 338
rect 442 228 476 266
rect 442 122 476 194
rect 161 20 173 54
rect 207 20 245 54
rect 279 20 317 54
rect 351 20 363 54
<< viali >>
rect 173 1160 207 1194
rect 245 1160 279 1194
rect 317 1160 351 1194
rect 48 1058 82 1092
rect 48 986 82 1020
rect 48 914 82 948
rect 48 842 82 876
rect 48 770 82 804
rect 48 698 82 732
rect 48 626 82 660
rect 48 554 82 588
rect 48 482 82 516
rect 48 410 82 444
rect 48 338 82 372
rect 48 266 82 300
rect 48 194 82 228
rect 442 1058 476 1092
rect 442 986 476 1020
rect 442 914 476 948
rect 442 842 476 876
rect 442 770 476 804
rect 442 698 476 732
rect 442 626 476 660
rect 442 554 476 588
rect 442 482 476 516
rect 442 410 476 444
rect 442 338 476 372
rect 442 266 476 300
rect 442 194 476 228
rect 173 20 207 54
rect 245 20 279 54
rect 317 20 351 54
<< obsli1 >>
rect 159 98 193 1116
rect 245 98 279 1116
rect 331 98 365 1116
<< metal1 >>
rect 161 1194 363 1214
rect 161 1160 173 1194
rect 207 1160 245 1194
rect 279 1160 317 1194
rect 351 1160 363 1194
rect 161 1148 363 1160
rect 36 1092 94 1104
rect 36 1058 48 1092
rect 82 1058 94 1092
rect 36 1020 94 1058
rect 36 986 48 1020
rect 82 986 94 1020
rect 36 948 94 986
rect 36 914 48 948
rect 82 914 94 948
rect 36 876 94 914
rect 36 842 48 876
rect 82 842 94 876
rect 36 804 94 842
rect 36 770 48 804
rect 82 770 94 804
rect 36 732 94 770
rect 36 698 48 732
rect 82 698 94 732
rect 36 660 94 698
rect 36 626 48 660
rect 82 626 94 660
rect 36 588 94 626
rect 36 554 48 588
rect 82 554 94 588
rect 36 516 94 554
rect 36 482 48 516
rect 82 482 94 516
rect 36 444 94 482
rect 36 410 48 444
rect 82 410 94 444
rect 36 372 94 410
rect 36 338 48 372
rect 82 338 94 372
rect 36 300 94 338
rect 36 266 48 300
rect 82 266 94 300
rect 36 228 94 266
rect 36 194 48 228
rect 82 194 94 228
rect 36 110 94 194
rect 430 1092 488 1104
rect 430 1058 442 1092
rect 476 1058 488 1092
rect 430 1020 488 1058
rect 430 986 442 1020
rect 476 986 488 1020
rect 430 948 488 986
rect 430 914 442 948
rect 476 914 488 948
rect 430 876 488 914
rect 430 842 442 876
rect 476 842 488 876
rect 430 804 488 842
rect 430 770 442 804
rect 476 770 488 804
rect 430 732 488 770
rect 430 698 442 732
rect 476 698 488 732
rect 430 660 488 698
rect 430 626 442 660
rect 476 626 488 660
rect 430 588 488 626
rect 430 554 442 588
rect 476 554 488 588
rect 430 516 488 554
rect 430 482 442 516
rect 476 482 488 516
rect 430 444 488 482
rect 430 410 442 444
rect 476 410 488 444
rect 430 372 488 410
rect 430 338 442 372
rect 476 338 488 372
rect 430 300 488 338
rect 430 266 442 300
rect 476 266 488 300
rect 430 228 488 266
rect 430 194 442 228
rect 476 194 488 228
rect 430 110 488 194
rect 161 54 363 66
rect 161 20 173 54
rect 207 20 245 54
rect 279 20 317 54
rect 351 20 363 54
rect 161 0 363 20
<< obsm1 >>
rect 150 110 202 1104
rect 236 110 288 1104
rect 322 110 374 1104
<< metal2 >>
rect 10 632 514 1104
rect 10 110 514 582
<< labels >>
rlabel viali s 442 1058 476 1092 6 BULK
port 1 nsew
rlabel viali s 442 986 476 1020 6 BULK
port 1 nsew
rlabel viali s 442 914 476 948 6 BULK
port 1 nsew
rlabel viali s 442 842 476 876 6 BULK
port 1 nsew
rlabel viali s 442 770 476 804 6 BULK
port 1 nsew
rlabel viali s 442 698 476 732 6 BULK
port 1 nsew
rlabel viali s 442 626 476 660 6 BULK
port 1 nsew
rlabel viali s 442 554 476 588 6 BULK
port 1 nsew
rlabel viali s 442 482 476 516 6 BULK
port 1 nsew
rlabel viali s 442 410 476 444 6 BULK
port 1 nsew
rlabel viali s 442 338 476 372 6 BULK
port 1 nsew
rlabel viali s 442 266 476 300 6 BULK
port 1 nsew
rlabel viali s 442 194 476 228 6 BULK
port 1 nsew
rlabel viali s 48 1058 82 1092 6 BULK
port 1 nsew
rlabel viali s 48 986 82 1020 6 BULK
port 1 nsew
rlabel viali s 48 914 82 948 6 BULK
port 1 nsew
rlabel viali s 48 842 82 876 6 BULK
port 1 nsew
rlabel viali s 48 770 82 804 6 BULK
port 1 nsew
rlabel viali s 48 698 82 732 6 BULK
port 1 nsew
rlabel viali s 48 626 82 660 6 BULK
port 1 nsew
rlabel viali s 48 554 82 588 6 BULK
port 1 nsew
rlabel viali s 48 482 82 516 6 BULK
port 1 nsew
rlabel viali s 48 410 82 444 6 BULK
port 1 nsew
rlabel viali s 48 338 82 372 6 BULK
port 1 nsew
rlabel viali s 48 266 82 300 6 BULK
port 1 nsew
rlabel viali s 48 194 82 228 6 BULK
port 1 nsew
rlabel locali s 442 122 476 1092 6 BULK
port 1 nsew
rlabel locali s 48 122 82 1092 6 BULK
port 1 nsew
rlabel metal1 s 430 110 488 1104 6 BULK
port 1 nsew
rlabel metal1 s 36 110 94 1104 6 BULK
port 1 nsew
rlabel metal2 s 10 632 514 1104 6 DRAIN
port 2 nsew
rlabel viali s 317 1160 351 1194 6 GATE
port 3 nsew
rlabel viali s 317 20 351 54 6 GATE
port 3 nsew
rlabel viali s 245 1160 279 1194 6 GATE
port 3 nsew
rlabel viali s 245 20 279 54 6 GATE
port 3 nsew
rlabel viali s 173 1160 207 1194 6 GATE
port 3 nsew
rlabel viali s 173 20 207 54 6 GATE
port 3 nsew
rlabel locali s 161 1160 363 1194 6 GATE
port 3 nsew
rlabel locali s 161 20 363 54 6 GATE
port 3 nsew
rlabel metal1 s 161 1148 363 1214 6 GATE
port 3 nsew
rlabel metal1 s 161 0 363 66 6 GATE
port 3 nsew
rlabel metal2 s 10 110 514 582 6 SOURCE
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 524 1214
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 9307698
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 9292238
<< end >>
