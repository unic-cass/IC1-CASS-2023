magic
tech sky130A
magscale 1 2
timestamp 1676037725
<< nwell >>
rect -38 261 682 582
<< pwell >>
rect 1 67 641 203
rect 30 21 641 67
rect 30 -17 64 21
<< locali >>
rect 207 401 273 493
rect 456 401 527 493
rect 207 367 527 401
rect 91 199 160 265
rect 306 181 362 367
rect 398 255 436 331
rect 472 299 527 367
rect 398 215 627 255
rect 306 161 371 181
rect 305 127 371 161
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 22 333 82 372
rect 116 367 167 527
rect 307 435 422 527
rect 22 299 272 333
rect 22 168 56 299
rect 206 215 272 299
rect 561 299 627 527
rect 22 102 69 168
rect 103 17 169 165
rect 216 93 271 181
rect 405 139 627 181
rect 405 93 455 139
rect 216 51 455 93
rect 489 17 523 105
rect 557 51 627 139
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
rlabel locali s 91 199 160 265 6 A_N
port 1 nsew signal input
rlabel locali s 398 215 627 255 6 B
port 2 nsew signal input
rlabel locali s 398 255 436 331 6 B
port 2 nsew signal input
rlabel metal1 s 0 -48 644 48 8 VGND
port 3 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 4 nsew ground bidirectional
rlabel pwell s 30 21 641 67 6 VNB
port 4 nsew ground bidirectional
rlabel pwell s 1 67 641 203 6 VNB
port 4 nsew ground bidirectional
rlabel nwell s -38 261 682 582 6 VPB
port 5 nsew power bidirectional
rlabel metal1 s 0 496 644 592 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 305 127 371 161 6 Y
port 7 nsew signal output
rlabel locali s 306 161 371 181 6 Y
port 7 nsew signal output
rlabel locali s 472 299 527 367 6 Y
port 7 nsew signal output
rlabel locali s 306 181 362 367 6 Y
port 7 nsew signal output
rlabel locali s 207 367 527 401 6 Y
port 7 nsew signal output
rlabel locali s 456 401 527 493 6 Y
port 7 nsew signal output
rlabel locali s 207 401 273 493 6 Y
port 7 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 644 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 1811168
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1804606
<< end >>
