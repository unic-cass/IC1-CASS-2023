magic
tech sky130B
magscale 1 2
timestamp 1676037725
<< nwell >>
rect 0 0 472 240
<< pmos >>
rect 95 36 125 204
rect 181 36 211 204
rect 267 36 297 204
rect 353 36 383 204
<< pdiff >>
rect 42 173 95 204
rect 42 139 50 173
rect 84 139 95 173
rect 42 101 95 139
rect 42 67 50 101
rect 84 67 95 101
rect 42 36 95 67
rect 125 173 181 204
rect 125 139 136 173
rect 170 139 181 173
rect 125 101 181 139
rect 125 67 136 101
rect 170 67 181 101
rect 125 36 181 67
rect 211 173 267 204
rect 211 139 222 173
rect 256 139 267 173
rect 211 101 267 139
rect 211 67 222 101
rect 256 67 267 101
rect 211 36 267 67
rect 297 173 353 204
rect 297 139 308 173
rect 342 139 353 173
rect 297 101 353 139
rect 297 67 308 101
rect 342 67 353 101
rect 297 36 353 67
rect 383 173 436 204
rect 383 139 394 173
rect 428 139 436 173
rect 383 101 436 139
rect 383 67 394 101
rect 428 67 436 101
rect 383 36 436 67
<< pdiffc >>
rect 50 139 84 173
rect 50 67 84 101
rect 136 139 170 173
rect 136 67 170 101
rect 222 139 256 173
rect 222 67 256 101
rect 308 139 342 173
rect 308 67 342 101
rect 394 139 428 173
rect 394 67 428 101
<< poly >>
rect 95 287 383 303
rect 95 253 120 287
rect 154 253 188 287
rect 222 253 256 287
rect 290 253 324 287
rect 358 253 383 287
rect 95 230 383 253
rect 95 204 125 230
rect 181 204 211 230
rect 267 204 297 230
rect 353 204 383 230
rect 95 10 125 36
rect 181 10 211 36
rect 267 10 297 36
rect 353 10 383 36
<< polycont >>
rect 120 253 154 287
rect 188 253 222 287
rect 256 253 290 287
rect 324 253 358 287
<< locali >>
rect 104 287 374 303
rect 104 253 114 287
rect 154 253 186 287
rect 222 253 256 287
rect 292 253 324 287
rect 364 253 374 287
rect 104 235 374 253
rect 50 173 84 189
rect 50 101 84 139
rect 50 51 84 67
rect 136 173 170 189
rect 136 101 170 139
rect 136 51 170 67
rect 222 173 256 189
rect 222 101 256 139
rect 222 51 256 67
rect 308 173 342 189
rect 308 101 342 139
rect 308 51 342 67
rect 394 173 428 189
rect 394 101 428 139
rect 394 51 428 67
<< viali >>
rect 114 253 120 287
rect 120 253 148 287
rect 186 253 188 287
rect 188 253 220 287
rect 258 253 290 287
rect 290 253 292 287
rect 330 253 358 287
rect 358 253 364 287
rect 50 139 84 173
rect 50 67 84 101
rect 136 139 170 173
rect 136 67 170 101
rect 222 139 256 173
rect 222 67 256 101
rect 308 139 342 173
rect 308 67 342 101
rect 394 139 428 173
rect 394 67 428 101
<< metal1 >>
rect 102 287 376 299
rect 102 253 114 287
rect 148 253 186 287
rect 220 253 258 287
rect 292 253 330 287
rect 364 253 376 287
rect 102 241 376 253
rect 44 173 90 189
rect 44 139 50 173
rect 84 139 90 173
rect 44 101 90 139
rect 44 67 50 101
rect 84 67 90 101
rect 44 -29 90 67
rect 127 178 179 189
rect 127 114 179 126
rect 127 51 179 62
rect 216 173 262 189
rect 216 139 222 173
rect 256 139 262 173
rect 216 101 262 139
rect 216 67 222 101
rect 256 67 262 101
rect 216 -29 262 67
rect 299 178 351 189
rect 299 114 351 126
rect 299 51 351 62
rect 388 173 434 189
rect 388 139 394 173
rect 428 139 434 173
rect 388 101 434 139
rect 388 67 394 101
rect 428 67 434 101
rect 388 -29 434 67
rect 44 -89 434 -29
<< via1 >>
rect 127 173 179 178
rect 127 139 136 173
rect 136 139 170 173
rect 170 139 179 173
rect 127 126 179 139
rect 127 101 179 114
rect 127 67 136 101
rect 136 67 170 101
rect 170 67 179 101
rect 127 62 179 67
rect 299 173 351 178
rect 299 139 308 173
rect 308 139 342 173
rect 342 139 351 173
rect 299 126 351 139
rect 299 101 351 114
rect 299 67 308 101
rect 308 67 342 101
rect 342 67 351 101
rect 299 62 351 67
<< metal2 >>
rect 120 188 186 197
rect 120 132 125 188
rect 181 132 186 188
rect 120 126 127 132
rect 179 126 186 132
rect 120 114 186 126
rect 120 108 127 114
rect 179 108 186 114
rect 120 52 125 108
rect 181 52 186 108
rect 120 43 186 52
rect 292 188 358 197
rect 292 132 297 188
rect 353 132 358 188
rect 292 126 299 132
rect 351 126 358 132
rect 292 114 358 126
rect 292 108 299 114
rect 351 108 358 114
rect 292 52 297 108
rect 353 52 358 108
rect 292 43 358 52
<< via2 >>
rect 125 178 181 188
rect 125 132 127 178
rect 127 132 179 178
rect 179 132 181 178
rect 125 62 127 108
rect 127 62 179 108
rect 179 62 181 108
rect 125 52 181 62
rect 297 178 353 188
rect 297 132 299 178
rect 299 132 351 178
rect 351 132 353 178
rect 297 62 299 108
rect 299 62 351 108
rect 351 62 353 108
rect 297 52 353 62
<< metal3 >>
rect 120 188 358 197
rect 120 132 125 188
rect 181 132 297 188
rect 353 132 358 188
rect 120 131 358 132
rect 120 108 186 131
rect 120 52 125 108
rect 181 52 186 108
rect 120 43 186 52
rect 292 108 358 131
rect 292 52 297 108
rect 353 52 358 108
rect 292 43 358 52
<< labels >>
flabel metal3 s 120 131 358 197 0 FreeSans 400 0 0 0 DRAIN
port 2 nsew
flabel metal1 s 44 -89 434 -29 0 FreeSans 400 0 0 0 SOURCE
port 3 nsew
flabel metal1 s 102 241 376 299 0 FreeSans 400 0 0 0 GATE
port 4 nsew
flabel nwell s 64 232 90 238 0 FreeSans 400 0 0 0 BULK
port 5 nsew
<< properties >>
string GDS_END 9129470
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 9122662
string path 8.125 4.725 8.125 1.275 
<< end >>
