magic
tech sky130B
magscale 1 2
timestamp 1676037725
<< locali >>
rect 11923 32808 11954 32846
rect 18056 32815 18086 32844
rect 18234 32813 18269 32838
rect 18234 32803 18242 32813
rect 16799 32751 16831 32795
rect 16965 32758 16996 32798
rect 18216 32779 18242 32781
rect 18420 32797 18456 32833
rect 18276 32779 18282 32781
rect 18216 32741 18282 32779
rect 19211 32744 19267 32788
rect 18216 32707 18242 32741
rect 18276 32707 18282 32741
<< viali >>
rect 18242 32779 18276 32813
rect 18242 32707 18276 32741
<< metal1 >>
rect 18522 33471 19108 33673
rect 17266 33331 17272 33383
rect 17324 33331 17336 33383
rect 17388 33331 17394 33383
rect 17875 33269 18003 33399
tri 27460 33067 27488 33095 ne
rect 18228 32814 18282 32825
rect 18280 32762 18282 32814
rect 18228 32750 18282 32762
rect 18280 32698 18282 32750
rect 18228 32692 18282 32698
rect 11513 32365 11551 32404
rect 18581 32317 19176 32472
rect 27140 32164 27192 32197
tri 27665 32194 27698 32227 ne
tri 27750 32194 27783 32227 nw
rect 19853 31506 19905 31512
rect 19853 31442 19905 31454
rect 19853 31384 19905 31390
rect 24432 30637 24634 30679
rect 25923 30641 26053 30683
rect 26335 30641 26537 30683
rect 26861 30641 27063 30683
rect 27575 30646 27721 30683
rect 27321 30418 27352 30562
tri 26781 29926 26787 29932 se
rect 26787 29926 26833 30165
rect 26781 29920 26833 29926
tri 27359 29893 27365 29899 nw
rect 26781 29856 26833 29868
rect 26781 29798 26833 29804
rect 24184 29706 24386 29748
rect 27091 24877 27137 24917
rect 27091 24740 27137 24781
rect 26721 23039 26752 23133
rect 27171 22975 27217 23015
rect 27289 22777 27335 22823
rect 26650 22321 26674 22407
rect 27289 21535 27335 21581
rect 25465 20856 25511 20902
rect 27247 20545 27293 20585
rect 25923 17881 26053 17923
rect 26335 17905 26537 17947
rect 24184 17775 24386 17817
rect 24710 17775 24912 17817
rect 25307 17775 25437 17817
rect 26861 17775 27063 17817
rect 27575 17775 27721 17812
<< via1 >>
rect 17272 33331 17324 33383
rect 17336 33331 17388 33383
rect 18228 32813 18280 32814
rect 18228 32779 18242 32813
rect 18242 32779 18276 32813
rect 18276 32779 18280 32813
rect 18228 32762 18280 32779
rect 18228 32741 18280 32750
rect 18228 32707 18242 32741
rect 18242 32707 18276 32741
rect 18276 32707 18280 32741
rect 18228 32698 18280 32707
rect 19853 31454 19905 31506
rect 19853 31390 19905 31442
rect 26781 29868 26833 29920
rect 26781 29804 26833 29856
<< metal2 >>
rect 11274 33500 11643 33685
rect 17260 33453 17269 33509
rect 17325 33453 17349 33509
rect 17405 33453 17414 33509
rect 17266 33383 17394 33453
tri 17394 33433 17414 33453 nw
rect 17266 33331 17272 33383
rect 17324 33331 17336 33383
rect 17388 33331 17394 33383
rect 20036 33327 20045 33383
rect 20101 33327 20125 33383
rect 20181 33327 20190 33383
tri 20037 33322 20042 33327 ne
tri 15704 33201 15760 33257 se
rect 15760 33201 16206 33257
rect 16262 33201 16307 33257
rect 16363 33201 16408 33257
rect 16464 33201 16473 33257
tri 15658 33155 15704 33201 se
rect 15704 33155 15712 33201
tri 15580 33077 15658 33155 se
rect 15658 33131 15712 33155
tri 15712 33131 15782 33201 nw
tri 15658 33077 15712 33131 nw
tri 15502 32999 15580 33077 se
tri 15580 32999 15658 33077 nw
tri 15787 33053 15865 33131 se
rect 15865 33075 16206 33131
rect 16262 33075 16307 33131
rect 16363 33075 16408 33131
rect 16464 33075 16473 33131
tri 15865 33053 15887 33075 nw
tri 15424 32921 15502 32999 se
tri 15502 32921 15580 32999 nw
tri 15709 32975 15787 33053 se
tri 15787 32975 15865 33053 nw
tri 15402 32899 15424 32921 se
rect 14766 32843 14775 32899
rect 14831 32843 14876 32899
rect 14932 32843 14977 32899
rect 15033 32843 15424 32899
tri 15424 32843 15502 32921 nw
tri 15631 32897 15709 32975 se
tri 15709 32897 15787 32975 nw
tri 15553 32819 15631 32897 se
tri 15631 32819 15709 32897 nw
rect 16933 32823 16942 32879
rect 16998 32823 17022 32879
rect 17078 32823 17087 32879
tri 15507 32773 15553 32819 se
rect 15553 32773 15565 32819
rect 14766 32717 14775 32773
rect 14831 32717 14876 32773
rect 14932 32717 14977 32773
rect 15033 32753 15565 32773
tri 15565 32753 15631 32819 nw
rect 16951 32805 17003 32823
rect 18228 32814 18280 32820
rect 18228 32753 18280 32762
rect 15033 32717 15529 32753
tri 15529 32717 15565 32753 nw
rect 18129 32697 18138 32753
rect 18194 32697 18218 32753
rect 18274 32750 18283 32753
rect 18280 32698 18283 32750
rect 18274 32697 18283 32698
rect 18228 32692 18280 32697
tri 19968 31516 20042 31590 se
rect 20042 31516 20097 33327
tri 20097 33292 20132 33327 nw
rect 19853 31506 20097 31516
rect 19905 31454 20097 31506
rect 19853 31442 20097 31454
rect 19905 31390 20097 31442
rect 19853 31384 20097 31390
rect 24402 29926 24458 29929
tri 24458 29926 24461 29929 sw
rect 24402 29920 26833 29926
tri 23413 29842 23444 29873 sw
rect 24458 29868 26781 29920
rect 24458 29864 26833 29868
rect 24402 29856 26833 29864
rect 24402 29840 26781 29856
tri 23409 29751 23443 29785 ne
rect 24458 29804 26781 29840
rect 24458 29798 26833 29804
rect 24402 29775 24458 29784
tri 24458 29775 24481 29798 nw
rect 2214 29431 2333 29489
rect 5497 29432 5506 29488
rect 5562 29432 5586 29488
rect 5642 29432 5651 29488
rect 2028 29282 2200 29364
rect 5291 29332 5300 29388
rect 5356 29332 5380 29388
rect 5436 29332 5445 29388
rect 4839 28595 4994 28884
rect 18919 27043 19027 27411
rect 22701 27039 22809 27407
rect 26693 23756 26745 23808
rect 25722 23272 25873 23315
rect 25032 21231 25088 21240
rect 25032 21151 25088 21175
rect 25032 21086 25088 21095
rect 25159 21137 25465 21146
rect 25215 21081 25465 21137
rect 25159 21057 25465 21081
rect 25215 21018 25465 21057
rect 25159 20992 25215 21001
rect 24780 20822 24836 20831
rect 25098 20781 25150 20828
rect 24780 20742 24836 20766
rect 24780 20677 24836 20686
rect 26781 20301 26833 20359
tri 27553 20199 27585 20231 ne
rect 24906 20105 24962 20114
tri 24962 20081 24995 20114 sw
rect 24962 20064 26751 20081
tri 26751 20064 26768 20081 sw
tri 27573 20064 27585 20076 se
rect 27585 20064 27671 20231
tri 27671 20199 27703 20231 nw
rect 24962 20049 26768 20064
rect 24906 20025 26768 20049
rect 24962 19995 26768 20025
rect 24906 19960 24962 19969
tri 24962 19961 24996 19995 nw
tri 26715 19942 26768 19995 ne
tri 26768 19942 26890 20064 sw
tri 27451 19942 27573 20064 se
rect 27573 20040 27671 20064
tri 27573 19942 27671 20040 nw
tri 26768 19856 26854 19942 ne
rect 26854 19856 27487 19942
tri 27487 19856 27573 19942 nw
tri 24644 18588 24654 18598 se
rect 24654 18589 24710 18598
tri 24710 18588 24720 18598 sw
tri 25406 18588 25410 18592 se
rect 25410 18588 25468 18592
tri 25468 18588 25472 18592 sw
rect 24654 18509 24710 18533
tri 24638 18444 24654 18460 ne
rect 24654 18444 24710 18453
tri 24710 18444 24726 18460 nw
tri 25376 18438 25410 18472 ne
tri 25466 18438 25500 18472 nw
rect 26621 17940 26673 17987
<< via2 >>
rect 17269 33453 17325 33509
rect 17349 33453 17405 33509
rect 20045 33327 20101 33383
rect 20125 33327 20181 33383
rect 16206 33201 16262 33257
rect 16307 33201 16363 33257
rect 16408 33201 16464 33257
rect 16206 33075 16262 33131
rect 16307 33075 16363 33131
rect 16408 33075 16464 33131
rect 14775 32843 14831 32899
rect 14876 32843 14932 32899
rect 14977 32843 15033 32899
rect 16942 32823 16998 32879
rect 17022 32823 17078 32879
rect 14775 32717 14831 32773
rect 14876 32717 14932 32773
rect 14977 32717 15033 32773
rect 18138 32697 18194 32753
rect 18218 32750 18274 32753
rect 18218 32698 18228 32750
rect 18228 32698 18274 32750
rect 18218 32697 18274 32698
rect 24402 29864 24458 29920
rect 24402 29784 24458 29840
rect 5506 29432 5562 29488
rect 5586 29432 5642 29488
rect 5300 29332 5356 29388
rect 5380 29332 5436 29388
rect 25032 21175 25088 21231
rect 25032 21095 25088 21151
rect 25159 21081 25215 21137
rect 25159 21001 25215 21057
rect 24780 20766 24836 20822
rect 24780 20686 24836 20742
rect 24906 20049 24962 20105
rect 24906 19969 24962 20025
rect 24654 18533 24710 18589
rect 24654 18453 24710 18509
<< metal3 >>
rect 17264 33509 23690 33514
rect 17264 33453 17269 33509
rect 17325 33453 17349 33509
rect 17405 33488 23690 33509
tri 23690 33488 23716 33514 sw
rect 17405 33453 23716 33488
rect 17264 33448 23716 33453
tri 23662 33394 23716 33448 ne
tri 23716 33394 23810 33488 sw
rect 20040 33383 23635 33388
rect 20040 33327 20045 33383
rect 20101 33327 20125 33383
rect 20181 33333 23635 33383
tri 23635 33333 23690 33388 sw
tri 23716 33333 23777 33394 ne
rect 23777 33333 23810 33394
rect 20181 33327 23690 33333
rect 20040 33322 23690 33327
rect 16183 33257 23581 33262
rect 16183 33201 16206 33257
rect 16262 33201 16307 33257
rect 16363 33201 16408 33257
rect 16464 33246 23581 33257
tri 23581 33246 23597 33262 sw
tri 23607 33246 23683 33322 ne
rect 23683 33246 23690 33322
tri 23690 33246 23777 33333 sw
tri 23777 33300 23810 33333 ne
tri 23810 33300 23904 33394 sw
rect 16464 33201 23597 33246
rect 16183 33196 23597 33201
tri 23553 33168 23581 33196 ne
rect 23581 33192 23597 33196
tri 23597 33192 23651 33246 sw
rect 23581 33168 23651 33192
rect 16183 33131 23527 33136
rect 16183 33075 16206 33131
rect 16262 33075 16307 33131
rect 16363 33075 16408 33131
rect 16464 33098 23527 33131
tri 23527 33098 23565 33136 sw
tri 23581 33098 23651 33168 ne
tri 23651 33160 23683 33192 sw
tri 23683 33160 23769 33246 ne
rect 23769 33239 23777 33246
tri 23777 33239 23784 33246 sw
tri 23810 33239 23871 33300 ne
rect 23871 33239 23904 33300
rect 23769 33160 23784 33239
rect 23651 33098 23683 33160
tri 23683 33098 23745 33160 sw
tri 23769 33152 23777 33160 ne
rect 23777 33152 23784 33160
tri 23784 33152 23871 33239 sw
tri 23871 33206 23904 33239 ne
tri 23904 33206 23998 33300 sw
rect 16464 33075 23565 33098
rect 16183 33070 23565 33075
tri 23499 33042 23527 33070 ne
rect 23527 33044 23565 33070
tri 23565 33044 23619 33098 sw
rect 23527 33042 23619 33044
rect 16649 32982 23473 33010
tri 23473 32982 23501 33010 sw
tri 23527 32982 23587 33042 ne
rect 23587 33012 23619 33042
tri 23619 33012 23651 33044 sw
tri 23651 33012 23737 33098 ne
rect 23737 33066 23745 33098
tri 23745 33066 23777 33098 sw
tri 23777 33066 23863 33152 ne
rect 23863 33145 23871 33152
tri 23871 33145 23878 33152 sw
tri 23904 33145 23965 33206 ne
rect 23965 33145 23998 33206
rect 23863 33066 23878 33145
rect 23737 33012 23777 33066
rect 23587 32982 23651 33012
rect 16649 32944 23501 32982
tri 5485 32776 5613 32904 se
rect 5613 32899 15041 32904
rect 5613 32843 14775 32899
rect 14831 32843 14876 32899
rect 14932 32843 14977 32899
rect 15033 32843 15041 32899
tri 23445 32896 23493 32944 ne
rect 23493 32896 23501 32944
tri 23501 32896 23587 32982 sw
tri 23587 32950 23619 32982 ne
rect 23619 32950 23651 32982
tri 23651 32950 23713 33012 sw
tri 23737 33004 23745 33012 ne
rect 23745 33004 23777 33012
tri 23777 33004 23839 33066 sw
tri 23863 33058 23871 33066 ne
rect 23871 33058 23878 33066
tri 23878 33058 23965 33145 sw
tri 23965 33112 23998 33145 ne
tri 23998 33112 24092 33206 sw
rect 5613 32838 15041 32843
rect 16937 32879 23419 32884
tri 5613 32776 5675 32838 nw
rect 16937 32823 16942 32879
rect 16998 32823 17022 32879
rect 17078 32834 23419 32879
tri 23419 32834 23469 32884 sw
tri 23493 32834 23555 32896 ne
rect 23555 32888 23587 32896
tri 23587 32888 23595 32896 sw
tri 23619 32888 23681 32950 ne
rect 23681 32918 23713 32950
tri 23713 32918 23745 32950 sw
tri 23745 32918 23831 33004 ne
rect 23831 32972 23839 33004
tri 23839 32972 23871 33004 sw
tri 23871 32972 23957 33058 ne
rect 23957 33051 23965 33058
tri 23965 33051 23972 33058 sw
tri 23998 33051 24059 33112 ne
rect 24059 33051 24092 33112
rect 23957 32972 23972 33051
rect 23831 32918 23871 32972
rect 23681 32888 23745 32918
rect 23555 32834 23595 32888
rect 17078 32823 23469 32834
rect 16937 32818 23469 32823
tri 5747 32776 5749 32778 se
rect 5749 32776 15041 32778
tri 5375 32666 5485 32776 se
rect 5485 32666 5503 32776
tri 5503 32666 5613 32776 nw
tri 5637 32666 5747 32776 se
rect 5747 32773 15041 32776
rect 5747 32717 14775 32773
rect 14831 32717 14876 32773
rect 14932 32717 14977 32773
rect 15033 32717 15041 32773
rect 5747 32712 15041 32717
rect 18133 32753 23365 32758
rect 5747 32666 5749 32712
tri 5295 29393 5375 29473 se
rect 5375 29393 5441 32666
tri 5441 32604 5503 32666 nw
tri 5598 32627 5637 32666 se
rect 5637 32627 5749 32666
tri 5749 32627 5834 32712 nw
rect 18133 32697 18138 32753
rect 18194 32697 18218 32753
rect 18274 32748 23365 32753
tri 23365 32748 23375 32758 sw
tri 23391 32748 23461 32818 ne
rect 23461 32748 23469 32818
tri 23469 32748 23555 32834 sw
tri 23555 32802 23587 32834 ne
rect 23587 32802 23595 32834
tri 23595 32802 23681 32888 sw
tri 23681 32856 23713 32888 ne
rect 23713 32856 23745 32888
tri 23745 32856 23807 32918 sw
tri 23831 32910 23839 32918 ne
rect 23839 32910 23871 32918
tri 23871 32910 23933 32972 sw
tri 23957 32964 23965 32972 ne
rect 23965 32964 23972 32972
tri 23972 32964 24059 33051 sw
tri 24059 33018 24092 33051 ne
tri 24092 33018 24186 33112 sw
rect 18274 32697 23375 32748
rect 18133 32694 23375 32697
tri 23375 32694 23429 32748 sw
rect 18133 32692 23429 32694
tri 5575 32604 5598 32627 se
rect 5598 32604 5602 32627
tri 5501 32530 5575 32604 se
rect 5575 32530 5602 32604
rect 5501 32480 5602 32530
tri 5602 32480 5749 32627 nw
tri 23337 32600 23429 32692 ne
tri 23429 32686 23437 32694 sw
tri 23461 32686 23523 32748 ne
rect 23523 32740 23555 32748
tri 23555 32740 23563 32748 sw
tri 23587 32740 23649 32802 ne
rect 23649 32794 23681 32802
tri 23681 32794 23689 32802 sw
tri 23713 32794 23775 32856 ne
rect 23775 32824 23807 32856
tri 23807 32824 23839 32856 sw
tri 23839 32824 23925 32910 ne
rect 23925 32878 23933 32910
tri 23933 32878 23965 32910 sw
tri 23965 32878 24051 32964 ne
rect 24051 32957 24059 32964
tri 24059 32957 24066 32964 sw
tri 24092 32957 24153 33018 ne
rect 24153 32957 24186 33018
rect 24051 32878 24066 32957
rect 23925 32824 23965 32878
rect 23775 32794 23839 32824
rect 23649 32740 23689 32794
rect 23523 32686 23563 32740
rect 23429 32600 23437 32686
tri 23437 32600 23523 32686 sw
tri 23523 32654 23555 32686 ne
rect 23555 32654 23563 32686
tri 23563 32654 23649 32740 sw
tri 23649 32708 23681 32740 ne
rect 23681 32708 23689 32740
tri 23689 32708 23775 32794 sw
tri 23775 32762 23807 32794 ne
rect 23807 32762 23839 32794
tri 23839 32762 23901 32824 sw
tri 23925 32816 23933 32824 ne
rect 23933 32816 23965 32824
tri 23965 32816 24027 32878 sw
tri 24051 32870 24059 32878 ne
rect 24059 32870 24066 32878
tri 24066 32870 24153 32957 sw
tri 24153 32924 24186 32957 ne
tri 24186 32924 24280 33018 sw
tri 23429 32506 23523 32600 ne
tri 23523 32592 23531 32600 sw
tri 23555 32592 23617 32654 ne
rect 23617 32646 23649 32654
tri 23649 32646 23657 32654 sw
tri 23681 32646 23743 32708 ne
rect 23743 32700 23775 32708
tri 23775 32700 23783 32708 sw
tri 23807 32700 23869 32762 ne
rect 23869 32730 23901 32762
tri 23901 32730 23933 32762 sw
tri 23933 32730 24019 32816 ne
rect 24019 32784 24027 32816
tri 24027 32784 24059 32816 sw
tri 24059 32784 24145 32870 ne
rect 24145 32863 24153 32870
tri 24153 32863 24160 32870 sw
tri 24186 32863 24247 32924 ne
rect 24247 32863 24280 32924
rect 24145 32784 24160 32863
rect 24019 32730 24059 32784
rect 23869 32700 23933 32730
rect 23743 32646 23783 32700
rect 23617 32592 23657 32646
rect 23523 32506 23531 32592
tri 23531 32506 23617 32592 sw
tri 23617 32560 23649 32592 ne
rect 23649 32560 23657 32592
tri 23657 32560 23743 32646 sw
tri 23743 32614 23775 32646 ne
rect 23775 32614 23783 32646
tri 23783 32614 23869 32700 sw
tri 23869 32668 23901 32700 ne
rect 23901 32668 23933 32700
tri 23933 32668 23995 32730 sw
tri 24019 32722 24027 32730 ne
rect 24027 32722 24059 32730
tri 24059 32722 24121 32784 sw
tri 24145 32776 24153 32784 ne
rect 24153 32776 24160 32784
tri 24160 32776 24247 32863 sw
tri 24247 32830 24280 32863 ne
tri 24280 32830 24374 32924 sw
rect 5501 29493 5567 32480
tri 5567 32445 5602 32480 nw
tri 23523 32412 23617 32506 ne
tri 23617 32498 23625 32506 sw
tri 23649 32498 23711 32560 ne
rect 23711 32552 23743 32560
tri 23743 32552 23751 32560 sw
tri 23775 32552 23837 32614 ne
rect 23837 32606 23869 32614
tri 23869 32606 23877 32614 sw
tri 23901 32606 23963 32668 ne
rect 23963 32636 23995 32668
tri 23995 32636 24027 32668 sw
tri 24027 32636 24113 32722 ne
rect 24113 32690 24121 32722
tri 24121 32690 24153 32722 sw
tri 24153 32690 24239 32776 ne
rect 24239 32769 24247 32776
tri 24247 32769 24254 32776 sw
tri 24280 32769 24341 32830 ne
rect 24341 32769 24374 32830
rect 24239 32690 24254 32769
rect 24113 32636 24153 32690
rect 23963 32606 24027 32636
rect 23837 32552 23877 32606
rect 23711 32498 23751 32552
rect 23617 32412 23625 32498
tri 23625 32412 23711 32498 sw
tri 23711 32466 23743 32498 ne
rect 23743 32466 23751 32498
tri 23751 32466 23837 32552 sw
tri 23837 32520 23869 32552 ne
rect 23869 32520 23877 32552
tri 23877 32520 23963 32606 sw
tri 23963 32574 23995 32606 ne
rect 23995 32574 24027 32606
tri 24027 32574 24089 32636 sw
tri 24113 32628 24121 32636 ne
rect 24121 32628 24153 32636
tri 24153 32628 24215 32690 sw
tri 24239 32682 24247 32690 ne
rect 24247 32682 24254 32690
tri 24254 32682 24341 32769 sw
tri 24341 32736 24374 32769 ne
tri 24374 32736 24468 32830 sw
tri 23617 32318 23711 32412 ne
tri 23711 32404 23719 32412 sw
tri 23743 32404 23805 32466 ne
rect 23805 32458 23837 32466
tri 23837 32458 23845 32466 sw
tri 23869 32458 23931 32520 ne
rect 23931 32512 23963 32520
tri 23963 32512 23971 32520 sw
tri 23995 32512 24057 32574 ne
rect 24057 32542 24089 32574
tri 24089 32542 24121 32574 sw
tri 24121 32542 24207 32628 ne
rect 24207 32596 24215 32628
tri 24215 32596 24247 32628 sw
tri 24247 32596 24333 32682 ne
rect 24333 32675 24341 32682
tri 24341 32675 24348 32682 sw
tri 24374 32675 24435 32736 ne
rect 24435 32675 24468 32736
rect 24333 32596 24348 32675
rect 24207 32542 24247 32596
rect 24057 32512 24121 32542
rect 23931 32458 23971 32512
rect 23805 32404 23845 32458
rect 23711 32318 23719 32404
tri 23719 32318 23805 32404 sw
tri 23805 32372 23837 32404 ne
rect 23837 32372 23845 32404
tri 23845 32372 23931 32458 sw
tri 23931 32426 23963 32458 ne
rect 23963 32426 23971 32458
tri 23971 32426 24057 32512 sw
tri 24057 32480 24089 32512 ne
rect 24089 32480 24121 32512
tri 24121 32480 24183 32542 sw
tri 24207 32534 24215 32542 ne
rect 24215 32534 24247 32542
tri 24247 32534 24309 32596 sw
tri 24333 32588 24341 32596 ne
rect 24341 32588 24348 32596
tri 24348 32588 24435 32675 sw
tri 24435 32642 24468 32675 ne
tri 24468 32642 24562 32736 sw
tri 23711 32224 23805 32318 ne
tri 23805 32310 23813 32318 sw
tri 23837 32310 23899 32372 ne
rect 23899 32364 23931 32372
tri 23931 32364 23939 32372 sw
tri 23963 32364 24025 32426 ne
rect 24025 32418 24057 32426
tri 24057 32418 24065 32426 sw
tri 24089 32418 24151 32480 ne
rect 24151 32448 24183 32480
tri 24183 32448 24215 32480 sw
tri 24215 32448 24301 32534 ne
rect 24301 32502 24309 32534
tri 24309 32502 24341 32534 sw
tri 24341 32502 24427 32588 ne
rect 24427 32581 24435 32588
tri 24435 32581 24442 32588 sw
tri 24468 32581 24529 32642 ne
rect 24529 32581 24562 32642
rect 24427 32502 24442 32581
rect 24301 32448 24341 32502
rect 24151 32418 24215 32448
rect 24025 32364 24065 32418
rect 23899 32310 23939 32364
rect 23805 32224 23813 32310
tri 23813 32224 23899 32310 sw
tri 23899 32278 23931 32310 ne
rect 23931 32278 23939 32310
tri 23939 32278 24025 32364 sw
tri 24025 32332 24057 32364 ne
rect 24057 32332 24065 32364
tri 24065 32332 24151 32418 sw
tri 24151 32386 24183 32418 ne
rect 24183 32386 24215 32418
tri 24215 32386 24277 32448 sw
tri 24301 32440 24309 32448 ne
rect 24309 32440 24341 32448
tri 24341 32440 24403 32502 sw
tri 24427 32494 24435 32502 ne
rect 24435 32494 24442 32502
tri 24442 32494 24529 32581 sw
tri 24529 32548 24562 32581 ne
tri 24562 32548 24656 32642 sw
tri 23805 32130 23899 32224 ne
tri 23899 32216 23907 32224 sw
tri 23931 32216 23993 32278 ne
rect 23993 32270 24025 32278
tri 24025 32270 24033 32278 sw
tri 24057 32270 24119 32332 ne
rect 24119 32324 24151 32332
tri 24151 32324 24159 32332 sw
tri 24183 32324 24245 32386 ne
rect 24245 32354 24277 32386
tri 24277 32354 24309 32386 sw
tri 24309 32354 24395 32440 ne
rect 24395 32408 24403 32440
tri 24403 32408 24435 32440 sw
tri 24435 32408 24521 32494 ne
rect 24521 32487 24529 32494
tri 24529 32487 24536 32494 sw
tri 24562 32487 24623 32548 ne
rect 24623 32487 24656 32548
rect 24521 32408 24536 32487
rect 24395 32354 24435 32408
rect 24245 32324 24309 32354
rect 24119 32270 24159 32324
rect 23993 32216 24033 32270
rect 23899 32130 23907 32216
tri 23907 32130 23993 32216 sw
tri 23993 32184 24025 32216 ne
rect 24025 32184 24033 32216
tri 24033 32184 24119 32270 sw
tri 24119 32238 24151 32270 ne
rect 24151 32238 24159 32270
tri 24159 32238 24245 32324 sw
tri 24245 32292 24277 32324 ne
rect 24277 32292 24309 32324
tri 24309 32292 24371 32354 sw
tri 24395 32346 24403 32354 ne
rect 24403 32346 24435 32354
tri 24435 32346 24497 32408 sw
tri 24521 32400 24529 32408 ne
rect 24529 32400 24536 32408
tri 24536 32400 24623 32487 sw
tri 24623 32454 24656 32487 ne
tri 24656 32454 24750 32548 sw
tri 23899 32036 23993 32130 ne
tri 23993 32122 24001 32130 sw
tri 24025 32122 24087 32184 ne
rect 24087 32176 24119 32184
tri 24119 32176 24127 32184 sw
tri 24151 32176 24213 32238 ne
rect 24213 32230 24245 32238
tri 24245 32230 24253 32238 sw
tri 24277 32230 24339 32292 ne
rect 24339 32260 24371 32292
tri 24371 32260 24403 32292 sw
tri 24403 32260 24489 32346 ne
rect 24489 32314 24497 32346
tri 24497 32314 24529 32346 sw
tri 24529 32314 24615 32400 ne
rect 24615 32393 24623 32400
tri 24623 32393 24630 32400 sw
tri 24656 32393 24717 32454 ne
rect 24717 32393 24750 32454
rect 24615 32314 24630 32393
rect 24489 32260 24529 32314
rect 24339 32230 24403 32260
rect 24213 32176 24253 32230
rect 24087 32122 24127 32176
rect 23993 32036 24001 32122
tri 24001 32036 24087 32122 sw
tri 24087 32090 24119 32122 ne
rect 24119 32090 24127 32122
tri 24127 32090 24213 32176 sw
tri 24213 32144 24245 32176 ne
rect 24245 32144 24253 32176
tri 24253 32144 24339 32230 sw
tri 24339 32198 24371 32230 ne
rect 24371 32198 24403 32230
tri 24403 32198 24465 32260 sw
tri 24489 32252 24497 32260 ne
rect 24497 32252 24529 32260
tri 24529 32252 24591 32314 sw
tri 24615 32306 24623 32314 ne
rect 24623 32306 24630 32314
tri 24630 32306 24717 32393 sw
tri 24717 32360 24750 32393 ne
tri 24750 32360 24844 32454 sw
tri 23993 31942 24087 32036 ne
tri 24087 32028 24095 32036 sw
tri 24119 32028 24181 32090 ne
rect 24181 32082 24213 32090
tri 24213 32082 24221 32090 sw
tri 24245 32082 24307 32144 ne
rect 24307 32136 24339 32144
tri 24339 32136 24347 32144 sw
tri 24371 32136 24433 32198 ne
rect 24433 32166 24465 32198
tri 24465 32166 24497 32198 sw
tri 24497 32166 24583 32252 ne
rect 24583 32220 24591 32252
tri 24591 32220 24623 32252 sw
tri 24623 32220 24709 32306 ne
rect 24709 32299 24717 32306
tri 24717 32299 24724 32306 sw
tri 24750 32299 24811 32360 ne
rect 24811 32299 24844 32360
rect 24709 32220 24724 32299
rect 24583 32166 24623 32220
rect 24433 32136 24497 32166
rect 24307 32082 24347 32136
rect 24181 32028 24221 32082
rect 24087 31942 24095 32028
tri 24095 31942 24181 32028 sw
tri 24181 31996 24213 32028 ne
rect 24213 31996 24221 32028
tri 24221 31996 24307 32082 sw
tri 24307 32050 24339 32082 ne
rect 24339 32050 24347 32082
tri 24347 32050 24433 32136 sw
tri 24433 32104 24465 32136 ne
rect 24465 32104 24497 32136
tri 24497 32104 24559 32166 sw
tri 24583 32158 24591 32166 ne
rect 24591 32158 24623 32166
tri 24623 32158 24685 32220 sw
tri 24709 32212 24717 32220 ne
rect 24717 32212 24724 32220
tri 24724 32212 24811 32299 sw
tri 24811 32266 24844 32299 ne
tri 24844 32266 24938 32360 sw
tri 24087 31848 24181 31942 ne
tri 24181 31934 24189 31942 sw
tri 24213 31934 24275 31996 ne
rect 24275 31988 24307 31996
tri 24307 31988 24315 31996 sw
tri 24339 31988 24401 32050 ne
rect 24401 32042 24433 32050
tri 24433 32042 24441 32050 sw
tri 24465 32042 24527 32104 ne
rect 24527 32072 24559 32104
tri 24559 32072 24591 32104 sw
tri 24591 32072 24677 32158 ne
rect 24677 32126 24685 32158
tri 24685 32126 24717 32158 sw
tri 24717 32126 24803 32212 ne
rect 24803 32205 24811 32212
tri 24811 32205 24818 32212 sw
tri 24844 32205 24905 32266 ne
rect 24905 32205 24938 32266
rect 24803 32126 24818 32205
rect 24677 32072 24717 32126
rect 24527 32042 24591 32072
rect 24401 31988 24441 32042
rect 24275 31934 24315 31988
rect 24181 31848 24189 31934
tri 24189 31848 24275 31934 sw
tri 24275 31902 24307 31934 ne
rect 24307 31902 24315 31934
tri 24315 31902 24401 31988 sw
tri 24401 31956 24433 31988 ne
rect 24433 31956 24441 31988
tri 24441 31956 24527 32042 sw
tri 24527 32010 24559 32042 ne
rect 24559 32010 24591 32042
tri 24591 32010 24653 32072 sw
tri 24677 32064 24685 32072 ne
rect 24685 32064 24717 32072
tri 24717 32064 24779 32126 sw
tri 24803 32118 24811 32126 ne
rect 24811 32118 24818 32126
tri 24818 32118 24905 32205 sw
tri 24905 32172 24938 32205 ne
tri 24938 32172 25032 32266 sw
tri 24181 31754 24275 31848 ne
tri 24275 31840 24283 31848 sw
tri 24307 31840 24369 31902 ne
rect 24369 31894 24401 31902
tri 24401 31894 24409 31902 sw
tri 24433 31894 24495 31956 ne
rect 24495 31948 24527 31956
tri 24527 31948 24535 31956 sw
tri 24559 31948 24621 32010 ne
rect 24621 31978 24653 32010
tri 24653 31978 24685 32010 sw
tri 24685 31978 24771 32064 ne
rect 24771 32032 24779 32064
tri 24779 32032 24811 32064 sw
tri 24811 32032 24897 32118 ne
rect 24897 32111 24905 32118
tri 24905 32111 24912 32118 sw
tri 24938 32111 24999 32172 ne
rect 24999 32111 25032 32172
rect 24897 32032 24912 32111
rect 24771 31978 24811 32032
rect 24621 31948 24685 31978
rect 24495 31894 24535 31948
rect 24369 31840 24409 31894
rect 24275 31754 24283 31840
tri 24283 31754 24369 31840 sw
tri 24369 31808 24401 31840 ne
rect 24401 31808 24409 31840
tri 24409 31808 24495 31894 sw
tri 24495 31862 24527 31894 ne
rect 24527 31862 24535 31894
tri 24535 31862 24621 31948 sw
tri 24621 31916 24653 31948 ne
rect 24653 31916 24685 31948
tri 24685 31916 24747 31978 sw
tri 24771 31970 24779 31978 ne
rect 24779 31970 24811 31978
tri 24811 31970 24873 32032 sw
tri 24897 32024 24905 32032 ne
rect 24905 32024 24912 32032
tri 24912 32024 24999 32111 sw
tri 24999 32078 25032 32111 ne
tri 25032 32078 25126 32172 sw
tri 24275 31660 24369 31754 ne
tri 24369 31746 24377 31754 sw
tri 24401 31746 24463 31808 ne
rect 24463 31800 24495 31808
tri 24495 31800 24503 31808 sw
tri 24527 31800 24589 31862 ne
rect 24589 31854 24621 31862
tri 24621 31854 24629 31862 sw
tri 24653 31854 24715 31916 ne
rect 24715 31884 24747 31916
tri 24747 31884 24779 31916 sw
tri 24779 31884 24865 31970 ne
rect 24865 31938 24873 31970
tri 24873 31938 24905 31970 sw
tri 24905 31938 24991 32024 ne
rect 24991 32017 24999 32024
tri 24999 32017 25006 32024 sw
tri 25032 32017 25093 32078 ne
rect 25093 32017 25126 32078
rect 24991 31938 25006 32017
rect 24865 31884 24905 31938
rect 24715 31854 24779 31884
rect 24589 31800 24629 31854
rect 24463 31746 24503 31800
rect 24369 31660 24377 31746
tri 24377 31660 24463 31746 sw
tri 24463 31714 24495 31746 ne
rect 24495 31714 24503 31746
tri 24503 31714 24589 31800 sw
tri 24589 31768 24621 31800 ne
rect 24621 31768 24629 31800
tri 24629 31768 24715 31854 sw
tri 24715 31794 24775 31854 ne
rect 24775 31822 24779 31854
tri 24779 31822 24841 31884 sw
tri 24865 31876 24873 31884 ne
rect 24873 31876 24905 31884
tri 24905 31876 24967 31938 sw
tri 24991 31930 24999 31938 ne
rect 24999 31930 25006 31938
tri 25006 31930 25093 32017 sw
tri 25093 31984 25126 32017 ne
tri 25126 31984 25220 32078 sw
tri 25126 31956 25154 31984 ne
tri 24999 31902 25027 31930 ne
tri 24873 31848 24901 31876 ne
tri 24621 31740 24649 31768 ne
tri 24495 31686 24523 31714 ne
tri 24369 31632 24397 31660 ne
rect 24397 29920 24463 31660
rect 24397 29864 24402 29920
rect 24458 29864 24463 29920
rect 24397 29840 24463 29864
rect 24397 29784 24402 29840
rect 24458 29784 24463 29840
rect 24397 29767 24463 29784
tri 5567 29493 5647 29573 sw
rect 5501 29488 5647 29493
rect 5501 29432 5506 29488
rect 5562 29432 5586 29488
rect 5642 29432 5647 29488
rect 5501 29427 5647 29432
rect 5295 29388 5441 29393
rect 5295 29332 5300 29388
rect 5356 29332 5380 29388
rect 5436 29332 5441 29388
rect 5295 29327 5441 29332
rect 21299 27345 21892 27790
rect 24523 21096 24589 31714
rect 24649 18589 24715 31768
rect 24775 20822 24841 31822
rect 24775 20766 24780 20822
rect 24836 20766 24841 20822
rect 24775 20742 24841 20766
rect 24775 20686 24780 20742
rect 24836 20686 24841 20742
rect 24775 20677 24841 20686
rect 24901 20105 24967 31876
rect 25027 21231 25093 31930
rect 25027 21175 25032 21231
rect 25088 21175 25093 21231
rect 25027 21151 25093 21175
rect 25027 21095 25032 21151
rect 25088 21095 25093 21151
rect 25027 21090 25093 21095
rect 25154 21137 25220 31984
rect 25154 21081 25159 21137
rect 25215 21081 25220 21137
rect 25154 21057 25220 21081
rect 25154 21001 25159 21057
rect 25215 21001 25220 21057
rect 25154 20996 25220 21001
rect 24901 20049 24906 20105
rect 24962 20049 24967 20105
rect 24901 20025 24967 20049
rect 24901 19969 24906 20025
rect 24962 19969 24967 20025
rect 24901 19960 24967 19969
rect 24649 18533 24654 18589
rect 24710 18533 24715 18589
rect 24649 18509 24715 18533
rect 2646 18462 2686 18491
rect 24649 18453 24654 18509
rect 24710 18453 24715 18509
rect 24649 18444 24715 18453
use sky130_fd_io__gpio_ovtv2_obpredrvr_new_i2c_fix_leak_fix  sky130_fd_io__gpio_ovtv2_obpredrvr_new_i2c_fix_leak_fix_0
timestamp 1676037725
transform 1 0 -49 0 1 28727
box 255 -19630 28132 5180
use sky130_fd_io__gpio_ovtv2_obpredrvr_old  sky130_fd_io__gpio_ovtv2_obpredrvr_old_0
timestamp 1676037725
transform 0 1 23158 -1 0 30683
box -255 631 13433 4925
<< labels >>
flabel metal3 s 2646 18462 2686 18491 0 FreeSans 200 0 0 0 NGHS_H
port 2 nsew
flabel metal3 s 21299 27345 21892 27790 3 FreeSans 520 270 0 0 VGND_IO
port 3 nsew
flabel metal3 s 21595 27567 21595 27567 3 FreeSans 520 270 0 0 VGND_IO
flabel metal1 s 11513 32365 11551 32404 3 FreeSans 520 90 0 0 OE_I_H_N
port 5 nsew
flabel metal1 s 26335 17905 26537 17947 7 FreeSans 300 270 0 0 VGND_IO
port 3 nsew
flabel metal1 s 25923 17881 26053 17923 7 FreeSans 300 270 0 0 VGND_IO
port 3 nsew
flabel metal1 s 25307 17775 25437 17817 7 FreeSans 300 270 0 0 VGND_IO
port 3 nsew
flabel metal1 s 24184 17775 24386 17817 7 FreeSans 300 270 0 0 VGND_IO
port 3 nsew
flabel metal1 s 24184 29706 24386 29748 3 FreeSans 300 270 0 0 VGND_IO
port 3 nsew
flabel metal1 s 25923 30641 26053 30683 3 FreeSans 300 270 0 0 VGND_IO
port 3 nsew
flabel metal1 s 26335 30641 26537 30683 3 FreeSans 300 270 0 0 VGND_IO
port 3 nsew
flabel metal1 s 26861 17775 27063 17817 7 FreeSans 300 270 0 0 VCC_IO
port 6 nsew
flabel metal1 s 27575 17775 27721 17812 7 FreeSans 300 270 0 0 VCC_IO
port 6 nsew
flabel metal1 s 24710 17775 24912 17817 7 FreeSans 300 270 0 0 VCC_IO
port 6 nsew
flabel metal1 s 24432 30637 24634 30679 3 FreeSans 300 270 0 0 VCC_IO
port 6 nsew
flabel metal1 s 27575 30646 27721 30683 3 FreeSans 300 270 0 0 VCC_IO
port 6 nsew
flabel metal1 s 26861 30641 27063 30683 3 FreeSans 300 270 0 0 VCC_IO
port 6 nsew
flabel metal1 s 25465 20856 25511 20902 3 FreeSans 300 270 0 0 SLOW_H
port 7 nsew
flabel metal1 s 27321 30418 27352 30562 3 FreeSans 520 270 0 0 PUEN_H[1]
port 8 nsew
flabel metal1 s 26721 23039 26752 23133 3 FreeSans 520 270 0 0 PUEN_H[0]
port 9 nsew
flabel metal1 s 27091 24740 27137 24781 3 FreeSans 300 270 0 0 PU_H_N[3]
port 10 nsew
flabel metal1 s 27091 24877 27137 24917 7 FreeSans 300 270 0 0 PU_H_N[2]
port 11 nsew
flabel metal1 s 27247 20545 27293 20585 3 FreeSans 300 270 0 0 PU_H_N[1]
port 12 nsew
flabel metal1 s 27171 22975 27217 23015 3 FreeSans 300 270 0 0 PU_H_N[0]
port 13 nsew
flabel metal1 s 27289 21535 27335 21581 3 FreeSans 300 270 0 0 PD_H[1]
port 14 nsew
flabel metal1 s 18581 32317 19176 32472 3 FreeSans 520 90 0 0 VGND_IO
port 3 nsew
flabel metal1 s 18522 33471 19108 33673 3 FreeSans 520 90 0 0 VCC_IO
port 6 nsew
flabel metal1 s 27289 22777 27335 22823 3 FreeSans 300 270 0 0 PD_H[0]
port 15 nsew
flabel metal1 s 26650 22321 26674 22407 3 FreeSans 520 270 0 0 PDEN_H_N[0]
port 16 nsew
flabel metal2 s 4839 28595 4994 28884 3 FreeSans 520 180 0 0 VGND_IO
port 3 nsew
flabel metal2 s 4916 28739 4916 28739 3 FreeSans 520 180 0 0 VGND_IO
flabel metal2 s 11274 33500 11643 33685 3 FreeSans 520 90 0 0 VCC_IO
port 6 nsew
flabel metal2 s 2028 29282 2200 29364 3 FreeSans 520 0 0 0 PD_H[3]
port 18 nsew
flabel metal2 s 2114 29323 2114 29323 3 FreeSans 520 0 0 0 PD_H[3]
flabel metal2 s 2214 29431 2333 29489 3 FreeSans 520 0 0 0 PD_H[2]
port 19 nsew
flabel metal2 s 18919 27043 19027 27411 3 FreeSans 520 180 0 0 PAD
port 20 nsew
flabel metal2 s 22701 27039 22809 27407 3 FreeSans 520 0 0 0 PAD
port 20 nsew
flabel metal2 s 22755 27223 22755 27223 3 FreeSans 520 0 0 0 PAD
flabel metal2 s 25722 23272 25873 23315 3 FreeSans 520 270 0 0 PDEN_H_N[1]
port 21 nsew
flabel metal2 s 26781 20301 26833 20359 3 FreeSans 300 270 0 0 PD_H[3]
port 18 nsew
flabel metal2 s 25098 20781 25150 20828 3 FreeSans 300 270 0 0 PD_H[2]
port 19 nsew
flabel metal2 s 26621 17940 26673 17987 7 FreeSans 300 270 0 0 DRVLO_H_N
port 22 nsew
flabel metal2 s 26693 23756 26745 23808 3 FreeSans 300 270 0 0 DRVHI_H
port 23 nsew
flabel locali s 18234 32803 18269 32838 3 FreeSans 520 90 0 0 SLOW_H_N
port 24 nsew
flabel locali s 19211 32744 19267 32788 3 FreeSans 520 90 0 0 SLEW_CTL_H_N[0]
port 25 nsew
flabel locali s 18420 32797 18456 32833 3 FreeSans 520 90 0 0 SLEW_CTL_H[1]
port 26 nsew
flabel locali s 16965 32758 16996 32798 3 FreeSans 520 90 0 0 PDEN_H_N[1]
port 21 nsew
flabel locali s 11923 32808 11954 32846 3 FreeSans 520 90 0 0 PD_DIS_H
port 27 nsew
flabel locali s 18056 32815 18086 32844 3 FreeSans 520 90 0 0 I2C_MODE_H_N
port 28 nsew
flabel locali s 16799 32751 16831 32795 3 FreeSans 520 90 0 0 DRVLO_H_N
port 22 nsew
<< properties >>
string GDS_END 33635838
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 33619980
<< end >>
