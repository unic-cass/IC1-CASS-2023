magic
tech sky130A
magscale 1 2
timestamp 1676037725
<< pwell >>
rect 15 163 1347 817
<< mvnmos >>
rect 241 189 341 791
rect 397 189 497 791
rect 553 189 653 791
rect 709 189 809 791
rect 865 189 965 791
rect 1021 189 1121 791
<< mvndiff >>
rect 181 779 241 791
rect 181 745 196 779
rect 230 745 241 779
rect 181 711 241 745
rect 181 677 196 711
rect 230 677 241 711
rect 181 643 241 677
rect 181 609 196 643
rect 230 609 241 643
rect 181 575 241 609
rect 181 541 196 575
rect 230 541 241 575
rect 181 507 241 541
rect 181 473 196 507
rect 230 473 241 507
rect 181 439 241 473
rect 181 405 196 439
rect 230 405 241 439
rect 181 371 241 405
rect 181 337 196 371
rect 230 337 241 371
rect 181 303 241 337
rect 181 269 196 303
rect 230 269 241 303
rect 181 235 241 269
rect 181 201 196 235
rect 230 201 241 235
rect 181 189 241 201
rect 341 779 397 791
rect 341 745 352 779
rect 386 745 397 779
rect 341 711 397 745
rect 341 677 352 711
rect 386 677 397 711
rect 341 643 397 677
rect 341 609 352 643
rect 386 609 397 643
rect 341 575 397 609
rect 341 541 352 575
rect 386 541 397 575
rect 341 507 397 541
rect 341 473 352 507
rect 386 473 397 507
rect 341 439 397 473
rect 341 405 352 439
rect 386 405 397 439
rect 341 371 397 405
rect 341 337 352 371
rect 386 337 397 371
rect 341 303 397 337
rect 341 269 352 303
rect 386 269 397 303
rect 341 235 397 269
rect 341 201 352 235
rect 386 201 397 235
rect 341 189 397 201
rect 497 779 553 791
rect 497 745 508 779
rect 542 745 553 779
rect 497 711 553 745
rect 497 677 508 711
rect 542 677 553 711
rect 497 643 553 677
rect 497 609 508 643
rect 542 609 553 643
rect 497 575 553 609
rect 497 541 508 575
rect 542 541 553 575
rect 497 507 553 541
rect 497 473 508 507
rect 542 473 553 507
rect 497 439 553 473
rect 497 405 508 439
rect 542 405 553 439
rect 497 371 553 405
rect 497 337 508 371
rect 542 337 553 371
rect 497 303 553 337
rect 497 269 508 303
rect 542 269 553 303
rect 497 235 553 269
rect 497 201 508 235
rect 542 201 553 235
rect 497 189 553 201
rect 653 779 709 791
rect 653 745 664 779
rect 698 745 709 779
rect 653 711 709 745
rect 653 677 664 711
rect 698 677 709 711
rect 653 643 709 677
rect 653 609 664 643
rect 698 609 709 643
rect 653 575 709 609
rect 653 541 664 575
rect 698 541 709 575
rect 653 507 709 541
rect 653 473 664 507
rect 698 473 709 507
rect 653 439 709 473
rect 653 405 664 439
rect 698 405 709 439
rect 653 371 709 405
rect 653 337 664 371
rect 698 337 709 371
rect 653 303 709 337
rect 653 269 664 303
rect 698 269 709 303
rect 653 235 709 269
rect 653 201 664 235
rect 698 201 709 235
rect 653 189 709 201
rect 809 779 865 791
rect 809 745 820 779
rect 854 745 865 779
rect 809 711 865 745
rect 809 677 820 711
rect 854 677 865 711
rect 809 643 865 677
rect 809 609 820 643
rect 854 609 865 643
rect 809 575 865 609
rect 809 541 820 575
rect 854 541 865 575
rect 809 507 865 541
rect 809 473 820 507
rect 854 473 865 507
rect 809 439 865 473
rect 809 405 820 439
rect 854 405 865 439
rect 809 371 865 405
rect 809 337 820 371
rect 854 337 865 371
rect 809 303 865 337
rect 809 269 820 303
rect 854 269 865 303
rect 809 235 865 269
rect 809 201 820 235
rect 854 201 865 235
rect 809 189 865 201
rect 965 779 1021 791
rect 965 745 976 779
rect 1010 745 1021 779
rect 965 711 1021 745
rect 965 677 976 711
rect 1010 677 1021 711
rect 965 643 1021 677
rect 965 609 976 643
rect 1010 609 1021 643
rect 965 575 1021 609
rect 965 541 976 575
rect 1010 541 1021 575
rect 965 507 1021 541
rect 965 473 976 507
rect 1010 473 1021 507
rect 965 439 1021 473
rect 965 405 976 439
rect 1010 405 1021 439
rect 965 371 1021 405
rect 965 337 976 371
rect 1010 337 1021 371
rect 965 303 1021 337
rect 965 269 976 303
rect 1010 269 1021 303
rect 965 235 1021 269
rect 965 201 976 235
rect 1010 201 1021 235
rect 965 189 1021 201
rect 1121 779 1181 791
rect 1121 745 1132 779
rect 1166 745 1181 779
rect 1121 711 1181 745
rect 1121 677 1132 711
rect 1166 677 1181 711
rect 1121 643 1181 677
rect 1121 609 1132 643
rect 1166 609 1181 643
rect 1121 575 1181 609
rect 1121 541 1132 575
rect 1166 541 1181 575
rect 1121 507 1181 541
rect 1121 473 1132 507
rect 1166 473 1181 507
rect 1121 439 1181 473
rect 1121 405 1132 439
rect 1166 405 1181 439
rect 1121 371 1181 405
rect 1121 337 1132 371
rect 1166 337 1181 371
rect 1121 303 1181 337
rect 1121 269 1132 303
rect 1166 269 1181 303
rect 1121 235 1181 269
rect 1121 201 1132 235
rect 1166 201 1181 235
rect 1121 189 1181 201
<< mvndiffc >>
rect 196 745 230 779
rect 196 677 230 711
rect 196 609 230 643
rect 196 541 230 575
rect 196 473 230 507
rect 196 405 230 439
rect 196 337 230 371
rect 196 269 230 303
rect 196 201 230 235
rect 352 745 386 779
rect 352 677 386 711
rect 352 609 386 643
rect 352 541 386 575
rect 352 473 386 507
rect 352 405 386 439
rect 352 337 386 371
rect 352 269 386 303
rect 352 201 386 235
rect 508 745 542 779
rect 508 677 542 711
rect 508 609 542 643
rect 508 541 542 575
rect 508 473 542 507
rect 508 405 542 439
rect 508 337 542 371
rect 508 269 542 303
rect 508 201 542 235
rect 664 745 698 779
rect 664 677 698 711
rect 664 609 698 643
rect 664 541 698 575
rect 664 473 698 507
rect 664 405 698 439
rect 664 337 698 371
rect 664 269 698 303
rect 664 201 698 235
rect 820 745 854 779
rect 820 677 854 711
rect 820 609 854 643
rect 820 541 854 575
rect 820 473 854 507
rect 820 405 854 439
rect 820 337 854 371
rect 820 269 854 303
rect 820 201 854 235
rect 976 745 1010 779
rect 976 677 1010 711
rect 976 609 1010 643
rect 976 541 1010 575
rect 976 473 1010 507
rect 976 405 1010 439
rect 976 337 1010 371
rect 976 269 1010 303
rect 976 201 1010 235
rect 1132 745 1166 779
rect 1132 677 1166 711
rect 1132 609 1166 643
rect 1132 541 1166 575
rect 1132 473 1166 507
rect 1132 405 1166 439
rect 1132 337 1166 371
rect 1132 269 1166 303
rect 1132 201 1166 235
<< mvpsubdiff >>
rect 41 779 181 791
rect 41 201 60 779
rect 162 201 181 779
rect 41 189 181 201
rect 1181 779 1321 791
rect 1181 201 1200 779
rect 1302 201 1321 779
rect 1181 189 1321 201
<< mvpsubdiffcont >>
rect 60 201 162 779
rect 1200 201 1302 779
<< poly >>
rect 383 959 979 980
rect 190 867 341 883
rect 190 833 206 867
rect 240 833 341 867
rect 383 857 426 959
rect 936 857 979 959
rect 383 841 979 857
rect 1021 867 1172 883
rect 190 817 341 833
rect 241 791 341 817
rect 397 791 497 841
rect 553 791 653 841
rect 709 791 809 841
rect 865 791 965 841
rect 1021 833 1122 867
rect 1156 833 1172 867
rect 1021 817 1172 833
rect 1021 791 1121 817
rect 241 163 341 189
rect 190 147 341 163
rect 190 113 206 147
rect 240 113 341 147
rect 397 139 497 189
rect 553 139 653 189
rect 709 139 809 189
rect 865 139 965 189
rect 1021 163 1121 189
rect 1021 147 1172 163
rect 190 97 341 113
rect 383 123 979 139
rect 383 21 426 123
rect 936 21 979 123
rect 1021 113 1122 147
rect 1156 113 1172 147
rect 1021 97 1172 113
rect 383 0 979 21
<< polycont >>
rect 206 833 240 867
rect 426 857 936 959
rect 1122 833 1156 867
rect 206 113 240 147
rect 426 21 936 123
rect 1122 113 1156 147
<< locali >>
rect 400 961 962 980
rect 190 867 256 883
rect 190 833 206 867
rect 240 833 256 867
rect 400 855 412 961
rect 950 855 962 961
rect 400 843 962 855
rect 1106 867 1172 883
rect 190 817 256 833
rect 1106 833 1122 867
rect 1156 833 1172 867
rect 1106 817 1172 833
rect 190 795 230 817
rect 1132 795 1172 817
rect 41 779 230 795
rect 41 201 60 779
rect 162 745 196 779
rect 162 711 230 745
rect 162 677 196 711
rect 162 643 230 677
rect 162 609 196 643
rect 162 575 230 609
rect 162 541 196 575
rect 162 507 230 541
rect 162 473 196 507
rect 162 439 230 473
rect 162 405 196 439
rect 162 371 230 405
rect 162 337 196 371
rect 162 303 230 337
rect 162 269 196 303
rect 162 235 230 269
rect 162 201 196 235
rect 41 185 230 201
rect 352 779 386 795
rect 352 711 386 725
rect 352 643 386 653
rect 352 575 386 581
rect 352 507 386 509
rect 352 471 386 473
rect 352 399 386 405
rect 352 327 386 337
rect 352 255 386 269
rect 352 185 386 201
rect 508 779 542 795
rect 508 711 542 725
rect 508 643 542 653
rect 508 575 542 581
rect 508 507 542 509
rect 508 471 542 473
rect 508 399 542 405
rect 508 327 542 337
rect 508 255 542 269
rect 508 185 542 201
rect 664 779 698 795
rect 664 711 698 725
rect 664 643 698 653
rect 664 575 698 581
rect 664 507 698 509
rect 664 471 698 473
rect 664 399 698 405
rect 664 327 698 337
rect 664 255 698 269
rect 664 185 698 201
rect 820 779 854 795
rect 820 711 854 725
rect 820 643 854 653
rect 820 575 854 581
rect 820 507 854 509
rect 820 471 854 473
rect 820 399 854 405
rect 820 327 854 337
rect 820 255 854 269
rect 820 185 854 201
rect 976 779 1010 795
rect 976 711 1010 725
rect 976 643 1010 653
rect 976 575 1010 581
rect 976 507 1010 509
rect 976 471 1010 473
rect 976 399 1010 405
rect 976 327 1010 337
rect 976 255 1010 269
rect 976 185 1010 201
rect 1132 779 1321 795
rect 1166 745 1200 779
rect 1132 711 1200 745
rect 1166 677 1200 711
rect 1132 643 1200 677
rect 1166 609 1200 643
rect 1132 575 1200 609
rect 1166 541 1200 575
rect 1132 507 1200 541
rect 1166 473 1200 507
rect 1132 439 1200 473
rect 1166 405 1200 439
rect 1132 371 1200 405
rect 1166 337 1200 371
rect 1132 303 1200 337
rect 1166 269 1200 303
rect 1132 235 1200 269
rect 1166 201 1200 235
rect 1302 201 1321 779
rect 1132 185 1321 201
rect 190 163 230 185
rect 1132 163 1172 185
rect 190 147 256 163
rect 190 113 206 147
rect 240 113 256 147
rect 1106 147 1172 163
rect 190 97 256 113
rect 400 125 962 137
rect 400 19 412 125
rect 950 19 962 125
rect 1106 113 1122 147
rect 1156 113 1172 147
rect 1106 97 1172 113
rect 400 0 962 19
<< viali >>
rect 412 959 950 961
rect 412 857 426 959
rect 426 857 936 959
rect 936 857 950 959
rect 412 855 950 857
rect 60 725 94 759
rect 60 653 94 687
rect 60 581 94 615
rect 60 509 94 543
rect 60 437 94 471
rect 60 365 94 399
rect 60 293 94 327
rect 60 221 94 255
rect 352 745 386 759
rect 352 725 386 745
rect 352 677 386 687
rect 352 653 386 677
rect 352 609 386 615
rect 352 581 386 609
rect 352 541 386 543
rect 352 509 386 541
rect 352 439 386 471
rect 352 437 386 439
rect 352 371 386 399
rect 352 365 386 371
rect 352 303 386 327
rect 352 293 386 303
rect 352 235 386 255
rect 352 221 386 235
rect 508 745 542 759
rect 508 725 542 745
rect 508 677 542 687
rect 508 653 542 677
rect 508 609 542 615
rect 508 581 542 609
rect 508 541 542 543
rect 508 509 542 541
rect 508 439 542 471
rect 508 437 542 439
rect 508 371 542 399
rect 508 365 542 371
rect 508 303 542 327
rect 508 293 542 303
rect 508 235 542 255
rect 508 221 542 235
rect 664 745 698 759
rect 664 725 698 745
rect 664 677 698 687
rect 664 653 698 677
rect 664 609 698 615
rect 664 581 698 609
rect 664 541 698 543
rect 664 509 698 541
rect 664 439 698 471
rect 664 437 698 439
rect 664 371 698 399
rect 664 365 698 371
rect 664 303 698 327
rect 664 293 698 303
rect 664 235 698 255
rect 664 221 698 235
rect 820 745 854 759
rect 820 725 854 745
rect 820 677 854 687
rect 820 653 854 677
rect 820 609 854 615
rect 820 581 854 609
rect 820 541 854 543
rect 820 509 854 541
rect 820 439 854 471
rect 820 437 854 439
rect 820 371 854 399
rect 820 365 854 371
rect 820 303 854 327
rect 820 293 854 303
rect 820 235 854 255
rect 820 221 854 235
rect 976 745 1010 759
rect 976 725 1010 745
rect 976 677 1010 687
rect 976 653 1010 677
rect 976 609 1010 615
rect 976 581 1010 609
rect 976 541 1010 543
rect 976 509 1010 541
rect 976 439 1010 471
rect 976 437 1010 439
rect 976 371 1010 399
rect 976 365 1010 371
rect 976 303 1010 327
rect 976 293 1010 303
rect 976 235 1010 255
rect 976 221 1010 235
rect 1268 725 1302 759
rect 1268 653 1302 687
rect 1268 581 1302 615
rect 1268 509 1302 543
rect 1268 437 1302 471
rect 1268 365 1302 399
rect 1268 293 1302 327
rect 1268 221 1302 255
rect 412 123 950 125
rect 412 21 426 123
rect 426 21 936 123
rect 936 21 950 123
rect 412 19 950 21
<< metal1 >>
rect 400 961 962 980
rect 400 855 412 961
rect 950 855 962 961
rect 400 843 962 855
rect 41 759 100 771
rect 41 725 60 759
rect 94 725 100 759
rect 41 687 100 725
rect 41 653 60 687
rect 94 653 100 687
rect 41 615 100 653
rect 41 581 60 615
rect 94 581 100 615
rect 41 543 100 581
rect 41 509 60 543
rect 94 509 100 543
rect 41 471 100 509
rect 41 437 60 471
rect 94 437 100 471
rect 41 399 100 437
rect 41 365 60 399
rect 94 365 100 399
rect 41 327 100 365
rect 41 293 60 327
rect 94 293 100 327
rect 41 255 100 293
rect 41 221 60 255
rect 94 221 100 255
rect 41 209 100 221
rect 343 759 395 771
rect 343 725 352 759
rect 386 725 395 759
rect 343 687 395 725
rect 343 653 352 687
rect 386 653 395 687
rect 343 615 395 653
rect 343 581 352 615
rect 386 581 395 615
rect 343 543 395 581
rect 343 509 352 543
rect 386 509 395 543
rect 343 471 395 509
rect 343 459 352 471
rect 386 459 395 471
rect 343 399 395 407
rect 343 395 352 399
rect 386 395 395 399
rect 343 331 395 343
rect 343 267 395 279
rect 343 209 395 215
rect 499 765 551 771
rect 499 701 551 713
rect 499 637 551 649
rect 499 581 508 585
rect 542 581 551 585
rect 499 573 551 581
rect 499 509 508 521
rect 542 509 551 521
rect 499 471 551 509
rect 499 437 508 471
rect 542 437 551 471
rect 499 399 551 437
rect 499 365 508 399
rect 542 365 551 399
rect 499 327 551 365
rect 499 293 508 327
rect 542 293 551 327
rect 499 255 551 293
rect 499 221 508 255
rect 542 221 551 255
rect 499 209 551 221
rect 655 759 707 771
rect 655 725 664 759
rect 698 725 707 759
rect 655 687 707 725
rect 655 653 664 687
rect 698 653 707 687
rect 655 615 707 653
rect 655 581 664 615
rect 698 581 707 615
rect 655 543 707 581
rect 655 509 664 543
rect 698 509 707 543
rect 655 471 707 509
rect 655 459 664 471
rect 698 459 707 471
rect 655 399 707 407
rect 655 395 664 399
rect 698 395 707 399
rect 655 331 707 343
rect 655 267 707 279
rect 655 209 707 215
rect 811 765 863 771
rect 811 701 863 713
rect 811 637 863 649
rect 811 581 820 585
rect 854 581 863 585
rect 811 573 863 581
rect 811 509 820 521
rect 854 509 863 521
rect 811 471 863 509
rect 811 437 820 471
rect 854 437 863 471
rect 811 399 863 437
rect 811 365 820 399
rect 854 365 863 399
rect 811 327 863 365
rect 811 293 820 327
rect 854 293 863 327
rect 811 255 863 293
rect 811 221 820 255
rect 854 221 863 255
rect 811 209 863 221
rect 967 759 1019 771
rect 967 725 976 759
rect 1010 725 1019 759
rect 967 687 1019 725
rect 967 653 976 687
rect 1010 653 1019 687
rect 967 615 1019 653
rect 967 581 976 615
rect 1010 581 1019 615
rect 967 543 1019 581
rect 967 509 976 543
rect 1010 509 1019 543
rect 967 471 1019 509
rect 967 459 976 471
rect 1010 459 1019 471
rect 967 399 1019 407
rect 967 395 976 399
rect 1010 395 1019 399
rect 967 331 1019 343
rect 967 267 1019 279
rect 967 209 1019 215
rect 1262 759 1321 771
rect 1262 725 1268 759
rect 1302 725 1321 759
rect 1262 687 1321 725
rect 1262 653 1268 687
rect 1302 653 1321 687
rect 1262 615 1321 653
rect 1262 581 1268 615
rect 1302 581 1321 615
rect 1262 543 1321 581
rect 1262 509 1268 543
rect 1302 509 1321 543
rect 1262 471 1321 509
rect 1262 437 1268 471
rect 1302 437 1321 471
rect 1262 399 1321 437
rect 1262 365 1268 399
rect 1302 365 1321 399
rect 1262 327 1321 365
rect 1262 293 1268 327
rect 1302 293 1321 327
rect 1262 255 1321 293
rect 1262 221 1268 255
rect 1302 221 1321 255
rect 1262 209 1321 221
rect 400 125 962 137
rect 400 19 412 125
rect 950 19 962 125
rect 400 0 962 19
<< via1 >>
rect 343 437 352 459
rect 352 437 386 459
rect 386 437 395 459
rect 343 407 395 437
rect 343 365 352 395
rect 352 365 386 395
rect 386 365 395 395
rect 343 343 395 365
rect 343 327 395 331
rect 343 293 352 327
rect 352 293 386 327
rect 386 293 395 327
rect 343 279 395 293
rect 343 255 395 267
rect 343 221 352 255
rect 352 221 386 255
rect 386 221 395 255
rect 343 215 395 221
rect 499 759 551 765
rect 499 725 508 759
rect 508 725 542 759
rect 542 725 551 759
rect 499 713 551 725
rect 499 687 551 701
rect 499 653 508 687
rect 508 653 542 687
rect 542 653 551 687
rect 499 649 551 653
rect 499 615 551 637
rect 499 585 508 615
rect 508 585 542 615
rect 542 585 551 615
rect 499 543 551 573
rect 499 521 508 543
rect 508 521 542 543
rect 542 521 551 543
rect 655 437 664 459
rect 664 437 698 459
rect 698 437 707 459
rect 655 407 707 437
rect 655 365 664 395
rect 664 365 698 395
rect 698 365 707 395
rect 655 343 707 365
rect 655 327 707 331
rect 655 293 664 327
rect 664 293 698 327
rect 698 293 707 327
rect 655 279 707 293
rect 655 255 707 267
rect 655 221 664 255
rect 664 221 698 255
rect 698 221 707 255
rect 655 215 707 221
rect 811 759 863 765
rect 811 725 820 759
rect 820 725 854 759
rect 854 725 863 759
rect 811 713 863 725
rect 811 687 863 701
rect 811 653 820 687
rect 820 653 854 687
rect 854 653 863 687
rect 811 649 863 653
rect 811 615 863 637
rect 811 585 820 615
rect 820 585 854 615
rect 854 585 863 615
rect 811 543 863 573
rect 811 521 820 543
rect 820 521 854 543
rect 854 521 863 543
rect 967 437 976 459
rect 976 437 1010 459
rect 1010 437 1019 459
rect 967 407 1019 437
rect 967 365 976 395
rect 976 365 1010 395
rect 1010 365 1019 395
rect 967 343 1019 365
rect 967 327 1019 331
rect 967 293 976 327
rect 976 293 1010 327
rect 1010 293 1019 327
rect 967 279 1019 293
rect 967 255 1019 267
rect 967 221 976 255
rect 976 221 1010 255
rect 1010 221 1019 255
rect 967 215 1019 221
<< metal2 >>
rect 14 765 1348 771
rect 14 713 499 765
rect 551 713 811 765
rect 863 713 1348 765
rect 14 701 1348 713
rect 14 649 499 701
rect 551 649 811 701
rect 863 649 1348 701
rect 14 637 1348 649
rect 14 585 499 637
rect 551 585 811 637
rect 863 585 1348 637
rect 14 573 1348 585
rect 14 521 499 573
rect 551 521 811 573
rect 863 521 1348 573
rect 14 515 1348 521
rect 14 459 1348 465
rect 14 407 343 459
rect 395 407 655 459
rect 707 407 967 459
rect 1019 407 1348 459
rect 14 395 1348 407
rect 14 343 343 395
rect 395 343 655 395
rect 707 343 967 395
rect 1019 343 1348 395
rect 14 331 1348 343
rect 14 279 343 331
rect 395 279 655 331
rect 707 279 967 331
rect 1019 279 1348 331
rect 14 267 1348 279
rect 14 215 343 267
rect 395 215 655 267
rect 707 215 967 267
rect 1019 215 1348 267
rect 14 209 1348 215
<< labels >>
flabel metal1 s 628 853 729 893 0 FreeSans 400 0 0 0 GATE
port 2 nsew
flabel metal1 s 628 17 729 57 0 FreeSans 200 0 0 0 GATE
port 2 nsew
flabel metal2 s 35 602 70 699 0 FreeSans 400 270 0 0 DRAIN
port 1 nsew
flabel metal2 s 36 313 66 417 0 FreeSans 400 90 0 0 SOURCE
port 3 nsew
flabel comment s 993 490 993 490 0 FreeSans 300 0 0 0 S
flabel comment s 837 490 837 490 0 FreeSans 300 0 0 0 D
flabel comment s 681 490 681 490 0 FreeSans 300 0 0 0 S
flabel comment s 525 490 525 490 0 FreeSans 300 0 0 0 D
flabel comment s 369 490 369 490 0 FreeSans 300 0 0 0 S
flabel comment s 837 490 837 490 0 FreeSans 300 0 0 0 S
flabel comment s 681 490 681 490 0 FreeSans 300 0 0 0 S
flabel comment s 525 490 525 490 0 FreeSans 300 0 0 0 S
flabel comment s 369 490 369 490 0 FreeSans 300 0 0 0 S
flabel comment s 281 514 281 514 0 FreeSans 400 90 0 0 dummy_poly
flabel comment s 1069 516 1069 516 0 FreeSans 400 90 0 0 dummy_poly
flabel metal1 s 41 466 100 496 0 FreeSans 200 90 0 0 SUBSTRATE
port 4 nsew
flabel metal1 s 1262 469 1321 499 0 FreeSans 200 90 0 0 SUBSTRATE
port 4 nsew
<< properties >>
string GDS_END 8485672
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 8463118
string device primitive
<< end >>
