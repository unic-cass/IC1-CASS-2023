magic
tech sky130A
magscale 1 2
timestamp 1676037725
<< metal1 >>
rect 91 2168 97 2220
rect 149 2168 155 2220
rect 196 1130 230 2256
rect 272 1142 300 2256
rect 1339 2168 1345 2220
rect 1397 2168 1403 2220
rect 425 2068 477 2074
rect 425 2010 477 2016
rect 343 1294 395 1300
rect 343 1236 395 1242
rect 1444 1130 1478 2256
rect 1520 1142 1548 2256
rect 2587 2168 2593 2220
rect 2645 2168 2651 2220
rect 1673 2068 1725 2074
rect 1673 2010 1725 2016
rect 1591 1294 1643 1300
rect 1591 1236 1643 1242
rect 2692 1130 2726 2256
rect 2768 1142 2796 2256
rect 3835 2168 3841 2220
rect 3893 2168 3899 2220
rect 2921 2068 2973 2074
rect 2921 2010 2973 2016
rect 2839 1294 2891 1300
rect 2839 1236 2891 1242
rect 3940 1130 3974 2256
rect 4016 1142 4044 2256
rect 5083 2168 5089 2220
rect 5141 2168 5147 2220
rect 4169 2068 4221 2074
rect 4169 2010 4221 2016
rect 4087 1294 4139 1300
rect 4087 1236 4139 1242
rect 5188 1130 5222 2256
rect 5264 1142 5292 2256
rect 6331 2168 6337 2220
rect 6389 2168 6395 2220
rect 5417 2068 5469 2074
rect 5417 2010 5469 2016
rect 5335 1294 5387 1300
rect 5335 1236 5387 1242
rect 6436 1130 6470 2256
rect 6512 1142 6540 2256
rect 7579 2168 7585 2220
rect 7637 2168 7643 2220
rect 6665 2068 6717 2074
rect 6665 2010 6717 2016
rect 6583 1294 6635 1300
rect 6583 1236 6635 1242
rect 7684 1130 7718 2256
rect 7760 1142 7788 2256
rect 8827 2168 8833 2220
rect 8885 2168 8891 2220
rect 7913 2068 7965 2074
rect 7913 2010 7965 2016
rect 7831 1294 7883 1300
rect 7831 1236 7883 1242
rect 8932 1130 8966 2256
rect 9008 1142 9036 2256
rect 10075 2168 10081 2220
rect 10133 2168 10139 2220
rect 9161 2068 9213 2074
rect 9161 2010 9213 2016
rect 9079 1294 9131 1300
rect 9079 1236 9131 1242
rect 10180 1130 10214 2256
rect 10256 1142 10284 2256
rect 11323 2168 11329 2220
rect 11381 2168 11387 2220
rect 10409 2068 10461 2074
rect 10409 2010 10461 2016
rect 10327 1294 10379 1300
rect 10327 1236 10379 1242
rect 11428 1130 11462 2256
rect 11504 1142 11532 2256
rect 12571 2168 12577 2220
rect 12629 2168 12635 2220
rect 11657 2068 11709 2074
rect 11657 2010 11709 2016
rect 11575 1294 11627 1300
rect 11575 1236 11627 1242
rect 12676 1130 12710 2256
rect 12752 1142 12780 2256
rect 13819 2168 13825 2220
rect 13877 2168 13883 2220
rect 12905 2068 12957 2074
rect 12905 2010 12957 2016
rect 12823 1294 12875 1300
rect 12823 1236 12875 1242
rect 13924 1130 13958 2256
rect 14000 1142 14028 2256
rect 15067 2168 15073 2220
rect 15125 2168 15131 2220
rect 14153 2068 14205 2074
rect 14153 2010 14205 2016
rect 14071 1294 14123 1300
rect 14071 1236 14123 1242
rect 15172 1130 15206 2256
rect 15248 1142 15276 2256
rect 16315 2168 16321 2220
rect 16373 2168 16379 2220
rect 15401 2068 15453 2074
rect 15401 2010 15453 2016
rect 15319 1294 15371 1300
rect 15319 1236 15371 1242
rect 16420 1130 16454 2256
rect 16496 1142 16524 2256
rect 17563 2168 17569 2220
rect 17621 2168 17627 2220
rect 16649 2068 16701 2074
rect 16649 2010 16701 2016
rect 16567 1294 16619 1300
rect 16567 1236 16619 1242
rect 17668 1130 17702 2256
rect 17744 1142 17772 2256
rect 18811 2168 18817 2220
rect 18869 2168 18875 2220
rect 17897 2068 17949 2074
rect 17897 2010 17949 2016
rect 17815 1294 17867 1300
rect 17815 1236 17867 1242
rect 18916 1130 18950 2256
rect 18992 1142 19020 2256
rect 20059 2168 20065 2220
rect 20117 2168 20123 2220
rect 19145 2068 19197 2074
rect 19145 2010 19197 2016
rect 19063 1294 19115 1300
rect 19063 1236 19115 1242
rect 20164 1130 20198 2256
rect 20240 1142 20268 2256
rect 21307 2168 21313 2220
rect 21365 2168 21371 2220
rect 20393 2068 20445 2074
rect 20393 2010 20445 2016
rect 20311 1294 20363 1300
rect 20311 1236 20363 1242
rect 21412 1130 21446 2256
rect 21488 1142 21516 2256
rect 22555 2168 22561 2220
rect 22613 2168 22619 2220
rect 21641 2068 21693 2074
rect 21641 2010 21693 2016
rect 21559 1294 21611 1300
rect 21559 1236 21611 1242
rect 22660 1130 22694 2256
rect 22736 1142 22764 2256
rect 23803 2168 23809 2220
rect 23861 2168 23867 2220
rect 22889 2068 22941 2074
rect 22889 2010 22941 2016
rect 22807 1294 22859 1300
rect 22807 1236 22859 1242
rect 23908 1130 23942 2256
rect 23984 1142 24012 2256
rect 25051 2168 25057 2220
rect 25109 2168 25115 2220
rect 24137 2068 24189 2074
rect 24137 2010 24189 2016
rect 24055 1294 24107 1300
rect 24055 1236 24107 1242
rect 25156 1130 25190 2256
rect 25232 1142 25260 2256
rect 26299 2168 26305 2220
rect 26357 2168 26363 2220
rect 25385 2068 25437 2074
rect 25385 2010 25437 2016
rect 25303 1294 25355 1300
rect 25303 1236 25355 1242
rect 26404 1130 26438 2256
rect 26480 1142 26508 2256
rect 27547 2168 27553 2220
rect 27605 2168 27611 2220
rect 26633 2068 26685 2074
rect 26633 2010 26685 2016
rect 26551 1294 26603 1300
rect 26551 1236 26603 1242
rect 27652 1130 27686 2256
rect 27728 1142 27756 2256
rect 28795 2168 28801 2220
rect 28853 2168 28859 2220
rect 27881 2068 27933 2074
rect 27881 2010 27933 2016
rect 27799 1294 27851 1300
rect 27799 1236 27851 1242
rect 28900 1130 28934 2256
rect 28976 1142 29004 2256
rect 30043 2168 30049 2220
rect 30101 2168 30107 2220
rect 29129 2068 29181 2074
rect 29129 2010 29181 2016
rect 29047 1294 29099 1300
rect 29047 1236 29099 1242
rect 30148 1130 30182 2256
rect 30224 1142 30252 2256
rect 31291 2168 31297 2220
rect 31349 2168 31355 2220
rect 30377 2068 30429 2074
rect 30377 2010 30429 2016
rect 30295 1294 30347 1300
rect 30295 1236 30347 1242
rect 31396 1130 31430 2256
rect 31472 1142 31500 2256
rect 32539 2168 32545 2220
rect 32597 2168 32603 2220
rect 31625 2068 31677 2074
rect 31625 2010 31677 2016
rect 31543 1294 31595 1300
rect 31543 1236 31595 1242
rect 32644 1130 32678 2256
rect 32720 1142 32748 2256
rect 33787 2168 33793 2220
rect 33845 2168 33851 2220
rect 32873 2068 32925 2074
rect 32873 2010 32925 2016
rect 32791 1294 32843 1300
rect 32791 1236 32843 1242
rect 33892 1130 33926 2256
rect 33968 1142 33996 2256
rect 35035 2168 35041 2220
rect 35093 2168 35099 2220
rect 34121 2068 34173 2074
rect 34121 2010 34173 2016
rect 34039 1294 34091 1300
rect 34039 1236 34091 1242
rect 35140 1130 35174 2256
rect 35216 1142 35244 2256
rect 36283 2168 36289 2220
rect 36341 2168 36347 2220
rect 35369 2068 35421 2074
rect 35369 2010 35421 2016
rect 35287 1294 35339 1300
rect 35287 1236 35339 1242
rect 36388 1130 36422 2256
rect 36464 1142 36492 2256
rect 37531 2168 37537 2220
rect 37589 2168 37595 2220
rect 36617 2068 36669 2074
rect 36617 2010 36669 2016
rect 36535 1294 36587 1300
rect 36535 1236 36587 1242
rect 37636 1130 37670 2256
rect 37712 1142 37740 2256
rect 38779 2168 38785 2220
rect 38837 2168 38843 2220
rect 37865 2068 37917 2074
rect 37865 2010 37917 2016
rect 37783 1294 37835 1300
rect 37783 1236 37835 1242
rect 38884 1130 38918 2256
rect 38960 1142 38988 2256
rect 39113 2068 39165 2074
rect 39113 2010 39165 2016
rect 39031 1294 39083 1300
rect 39031 1236 39083 1242
rect 355 456 407 462
rect 355 398 407 404
rect 1603 456 1655 462
rect 1603 398 1655 404
rect 2851 456 2903 462
rect 2851 398 2903 404
rect 4099 456 4151 462
rect 4099 398 4151 404
rect 5347 456 5399 462
rect 5347 398 5399 404
rect 6595 456 6647 462
rect 6595 398 6647 404
rect 7843 456 7895 462
rect 7843 398 7895 404
rect 9091 456 9143 462
rect 9091 398 9143 404
rect 10339 456 10391 462
rect 10339 398 10391 404
rect 11587 456 11639 462
rect 11587 398 11639 404
rect 12835 456 12887 462
rect 12835 398 12887 404
rect 14083 456 14135 462
rect 14083 398 14135 404
rect 15331 456 15383 462
rect 15331 398 15383 404
rect 16579 456 16631 462
rect 16579 398 16631 404
rect 17827 456 17879 462
rect 17827 398 17879 404
rect 19075 456 19127 462
rect 19075 398 19127 404
rect 20323 456 20375 462
rect 20323 398 20375 404
rect 21571 456 21623 462
rect 21571 398 21623 404
rect 22819 456 22871 462
rect 22819 398 22871 404
rect 24067 456 24119 462
rect 24067 398 24119 404
rect 25315 456 25367 462
rect 25315 398 25367 404
rect 26563 456 26615 462
rect 26563 398 26615 404
rect 27811 456 27863 462
rect 27811 398 27863 404
rect 29059 456 29111 462
rect 29059 398 29111 404
rect 30307 456 30359 462
rect 30307 398 30359 404
rect 31555 456 31607 462
rect 31555 398 31607 404
rect 32803 456 32855 462
rect 32803 398 32855 404
rect 34051 456 34103 462
rect 34051 398 34103 404
rect 35299 456 35351 462
rect 35299 398 35351 404
rect 36547 456 36599 462
rect 36547 398 36599 404
rect 37795 456 37847 462
rect 37795 398 37847 404
rect 39043 456 39095 462
rect 39043 398 39095 404
rect 104 0 150 254
rect 355 134 407 140
rect 355 76 407 82
rect 1352 0 1398 254
rect 1603 134 1655 140
rect 1603 76 1655 82
rect 2600 0 2646 254
rect 2851 134 2903 140
rect 2851 76 2903 82
rect 3848 0 3894 254
rect 4099 134 4151 140
rect 4099 76 4151 82
rect 5096 0 5142 254
rect 5347 134 5399 140
rect 5347 76 5399 82
rect 6344 0 6390 254
rect 6595 134 6647 140
rect 6595 76 6647 82
rect 7592 0 7638 254
rect 7843 134 7895 140
rect 7843 76 7895 82
rect 8840 0 8886 254
rect 9091 134 9143 140
rect 9091 76 9143 82
rect 10088 0 10134 254
rect 10339 134 10391 140
rect 10339 76 10391 82
rect 11336 0 11382 254
rect 11587 134 11639 140
rect 11587 76 11639 82
rect 12584 0 12630 254
rect 12835 134 12887 140
rect 12835 76 12887 82
rect 13832 0 13878 254
rect 14083 134 14135 140
rect 14083 76 14135 82
rect 15080 0 15126 254
rect 15331 134 15383 140
rect 15331 76 15383 82
rect 16328 0 16374 254
rect 16579 134 16631 140
rect 16579 76 16631 82
rect 17576 0 17622 254
rect 17827 134 17879 140
rect 17827 76 17879 82
rect 18824 0 18870 254
rect 19075 134 19127 140
rect 19075 76 19127 82
rect 20072 0 20118 254
rect 20323 134 20375 140
rect 20323 76 20375 82
rect 21320 0 21366 254
rect 21571 134 21623 140
rect 21571 76 21623 82
rect 22568 0 22614 254
rect 22819 134 22871 140
rect 22819 76 22871 82
rect 23816 0 23862 254
rect 24067 134 24119 140
rect 24067 76 24119 82
rect 25064 0 25110 254
rect 25315 134 25367 140
rect 25315 76 25367 82
rect 26312 0 26358 254
rect 26563 134 26615 140
rect 26563 76 26615 82
rect 27560 0 27606 254
rect 27811 134 27863 140
rect 27811 76 27863 82
rect 28808 0 28854 254
rect 29059 134 29111 140
rect 29059 76 29111 82
rect 30056 0 30102 254
rect 30307 134 30359 140
rect 30307 76 30359 82
rect 31304 0 31350 254
rect 31555 134 31607 140
rect 31555 76 31607 82
rect 32552 0 32598 254
rect 32803 134 32855 140
rect 32803 76 32855 82
rect 33800 0 33846 254
rect 34051 134 34103 140
rect 34051 76 34103 82
rect 35048 0 35094 254
rect 35299 134 35351 140
rect 35299 76 35351 82
rect 36296 0 36342 254
rect 36547 134 36599 140
rect 36547 76 36599 82
rect 37544 0 37590 254
rect 37795 134 37847 140
rect 37795 76 37847 82
rect 38792 0 38838 254
rect 39043 134 39095 140
rect 39043 76 39095 82
<< via1 >>
rect 97 2168 149 2220
rect 1345 2168 1397 2220
rect 425 2016 477 2068
rect 343 1242 395 1294
rect 2593 2168 2645 2220
rect 1673 2016 1725 2068
rect 1591 1242 1643 1294
rect 3841 2168 3893 2220
rect 2921 2016 2973 2068
rect 2839 1242 2891 1294
rect 5089 2168 5141 2220
rect 4169 2016 4221 2068
rect 4087 1242 4139 1294
rect 6337 2168 6389 2220
rect 5417 2016 5469 2068
rect 5335 1242 5387 1294
rect 7585 2168 7637 2220
rect 6665 2016 6717 2068
rect 6583 1242 6635 1294
rect 8833 2168 8885 2220
rect 7913 2016 7965 2068
rect 7831 1242 7883 1294
rect 10081 2168 10133 2220
rect 9161 2016 9213 2068
rect 9079 1242 9131 1294
rect 11329 2168 11381 2220
rect 10409 2016 10461 2068
rect 10327 1242 10379 1294
rect 12577 2168 12629 2220
rect 11657 2016 11709 2068
rect 11575 1242 11627 1294
rect 13825 2168 13877 2220
rect 12905 2016 12957 2068
rect 12823 1242 12875 1294
rect 15073 2168 15125 2220
rect 14153 2016 14205 2068
rect 14071 1242 14123 1294
rect 16321 2168 16373 2220
rect 15401 2016 15453 2068
rect 15319 1242 15371 1294
rect 17569 2168 17621 2220
rect 16649 2016 16701 2068
rect 16567 1242 16619 1294
rect 18817 2168 18869 2220
rect 17897 2016 17949 2068
rect 17815 1242 17867 1294
rect 20065 2168 20117 2220
rect 19145 2016 19197 2068
rect 19063 1242 19115 1294
rect 21313 2168 21365 2220
rect 20393 2016 20445 2068
rect 20311 1242 20363 1294
rect 22561 2168 22613 2220
rect 21641 2016 21693 2068
rect 21559 1242 21611 1294
rect 23809 2168 23861 2220
rect 22889 2016 22941 2068
rect 22807 1242 22859 1294
rect 25057 2168 25109 2220
rect 24137 2016 24189 2068
rect 24055 1242 24107 1294
rect 26305 2168 26357 2220
rect 25385 2016 25437 2068
rect 25303 1242 25355 1294
rect 27553 2168 27605 2220
rect 26633 2016 26685 2068
rect 26551 1242 26603 1294
rect 28801 2168 28853 2220
rect 27881 2016 27933 2068
rect 27799 1242 27851 1294
rect 30049 2168 30101 2220
rect 29129 2016 29181 2068
rect 29047 1242 29099 1294
rect 31297 2168 31349 2220
rect 30377 2016 30429 2068
rect 30295 1242 30347 1294
rect 32545 2168 32597 2220
rect 31625 2016 31677 2068
rect 31543 1242 31595 1294
rect 33793 2168 33845 2220
rect 32873 2016 32925 2068
rect 32791 1242 32843 1294
rect 35041 2168 35093 2220
rect 34121 2016 34173 2068
rect 34039 1242 34091 1294
rect 36289 2168 36341 2220
rect 35369 2016 35421 2068
rect 35287 1242 35339 1294
rect 37537 2168 37589 2220
rect 36617 2016 36669 2068
rect 36535 1242 36587 1294
rect 38785 2168 38837 2220
rect 37865 2016 37917 2068
rect 37783 1242 37835 1294
rect 39113 2016 39165 2068
rect 39031 1242 39083 1294
rect 355 404 407 456
rect 1603 404 1655 456
rect 2851 404 2903 456
rect 4099 404 4151 456
rect 5347 404 5399 456
rect 6595 404 6647 456
rect 7843 404 7895 456
rect 9091 404 9143 456
rect 10339 404 10391 456
rect 11587 404 11639 456
rect 12835 404 12887 456
rect 14083 404 14135 456
rect 15331 404 15383 456
rect 16579 404 16631 456
rect 17827 404 17879 456
rect 19075 404 19127 456
rect 20323 404 20375 456
rect 21571 404 21623 456
rect 22819 404 22871 456
rect 24067 404 24119 456
rect 25315 404 25367 456
rect 26563 404 26615 456
rect 27811 404 27863 456
rect 29059 404 29111 456
rect 30307 404 30359 456
rect 31555 404 31607 456
rect 32803 404 32855 456
rect 34051 404 34103 456
rect 35299 404 35351 456
rect 36547 404 36599 456
rect 37795 404 37847 456
rect 39043 404 39095 456
rect 355 82 407 134
rect 1603 82 1655 134
rect 2851 82 2903 134
rect 4099 82 4151 134
rect 5347 82 5399 134
rect 6595 82 6647 134
rect 7843 82 7895 134
rect 9091 82 9143 134
rect 10339 82 10391 134
rect 11587 82 11639 134
rect 12835 82 12887 134
rect 14083 82 14135 134
rect 15331 82 15383 134
rect 16579 82 16631 134
rect 17827 82 17879 134
rect 19075 82 19127 134
rect 20323 82 20375 134
rect 21571 82 21623 134
rect 22819 82 22871 134
rect 24067 82 24119 134
rect 25315 82 25367 134
rect 26563 82 26615 134
rect 27811 82 27863 134
rect 29059 82 29111 134
rect 30307 82 30359 134
rect 31555 82 31607 134
rect 32803 82 32855 134
rect 34051 82 34103 134
rect 35299 82 35351 134
rect 36547 82 36599 134
rect 37795 82 37847 134
rect 39043 82 39095 134
<< metal2 >>
rect 95 2222 151 2231
rect 95 2157 151 2166
rect 1343 2222 1399 2231
rect 1343 2157 1399 2166
rect 2591 2222 2647 2231
rect 2591 2157 2647 2166
rect 3839 2222 3895 2231
rect 3839 2157 3895 2166
rect 5087 2222 5143 2231
rect 5087 2157 5143 2166
rect 6335 2222 6391 2231
rect 6335 2157 6391 2166
rect 7583 2222 7639 2231
rect 7583 2157 7639 2166
rect 8831 2222 8887 2231
rect 8831 2157 8887 2166
rect 10079 2222 10135 2231
rect 10079 2157 10135 2166
rect 11327 2222 11383 2231
rect 11327 2157 11383 2166
rect 12575 2222 12631 2231
rect 12575 2157 12631 2166
rect 13823 2222 13879 2231
rect 13823 2157 13879 2166
rect 15071 2222 15127 2231
rect 15071 2157 15127 2166
rect 16319 2222 16375 2231
rect 16319 2157 16375 2166
rect 17567 2222 17623 2231
rect 17567 2157 17623 2166
rect 18815 2222 18871 2231
rect 18815 2157 18871 2166
rect 20063 2222 20119 2231
rect 20063 2157 20119 2166
rect 21311 2222 21367 2231
rect 21311 2157 21367 2166
rect 22559 2222 22615 2231
rect 22559 2157 22615 2166
rect 23807 2222 23863 2231
rect 23807 2157 23863 2166
rect 25055 2222 25111 2231
rect 25055 2157 25111 2166
rect 26303 2222 26359 2231
rect 26303 2157 26359 2166
rect 27551 2222 27607 2231
rect 27551 2157 27607 2166
rect 28799 2222 28855 2231
rect 28799 2157 28855 2166
rect 30047 2222 30103 2231
rect 30047 2157 30103 2166
rect 31295 2222 31351 2231
rect 31295 2157 31351 2166
rect 32543 2222 32599 2231
rect 32543 2157 32599 2166
rect 33791 2222 33847 2231
rect 33791 2157 33847 2166
rect 35039 2222 35095 2231
rect 35039 2157 35095 2166
rect 36287 2222 36343 2231
rect 36287 2157 36343 2166
rect 37535 2222 37591 2231
rect 37535 2157 37591 2166
rect 38783 2222 38839 2231
rect 38783 2157 38839 2166
rect 423 2070 479 2079
rect 423 2005 479 2014
rect 1671 2070 1727 2079
rect 1671 2005 1727 2014
rect 2919 2070 2975 2079
rect 2919 2005 2975 2014
rect 4167 2070 4223 2079
rect 4167 2005 4223 2014
rect 5415 2070 5471 2079
rect 5415 2005 5471 2014
rect 6663 2070 6719 2079
rect 6663 2005 6719 2014
rect 7911 2070 7967 2079
rect 7911 2005 7967 2014
rect 9159 2070 9215 2079
rect 9159 2005 9215 2014
rect 10407 2070 10463 2079
rect 10407 2005 10463 2014
rect 11655 2070 11711 2079
rect 11655 2005 11711 2014
rect 12903 2070 12959 2079
rect 12903 2005 12959 2014
rect 14151 2070 14207 2079
rect 14151 2005 14207 2014
rect 15399 2070 15455 2079
rect 15399 2005 15455 2014
rect 16647 2070 16703 2079
rect 16647 2005 16703 2014
rect 17895 2070 17951 2079
rect 17895 2005 17951 2014
rect 19143 2070 19199 2079
rect 19143 2005 19199 2014
rect 20391 2070 20447 2079
rect 20391 2005 20447 2014
rect 21639 2070 21695 2079
rect 21639 2005 21695 2014
rect 22887 2070 22943 2079
rect 22887 2005 22943 2014
rect 24135 2070 24191 2079
rect 24135 2005 24191 2014
rect 25383 2070 25439 2079
rect 25383 2005 25439 2014
rect 26631 2070 26687 2079
rect 26631 2005 26687 2014
rect 27879 2070 27935 2079
rect 27879 2005 27935 2014
rect 29127 2070 29183 2079
rect 29127 2005 29183 2014
rect 30375 2070 30431 2079
rect 30375 2005 30431 2014
rect 31623 2070 31679 2079
rect 31623 2005 31679 2014
rect 32871 2070 32927 2079
rect 32871 2005 32927 2014
rect 34119 2070 34175 2079
rect 34119 2005 34175 2014
rect 35367 2070 35423 2079
rect 35367 2005 35423 2014
rect 36615 2070 36671 2079
rect 36615 2005 36671 2014
rect 37863 2070 37919 2079
rect 37863 2005 37919 2014
rect 39111 2070 39167 2079
rect 39111 2005 39167 2014
rect 341 1296 397 1305
rect 341 1231 397 1240
rect 1589 1296 1645 1305
rect 1589 1231 1645 1240
rect 2837 1296 2893 1305
rect 2837 1231 2893 1240
rect 4085 1296 4141 1305
rect 4085 1231 4141 1240
rect 5333 1296 5389 1305
rect 5333 1231 5389 1240
rect 6581 1296 6637 1305
rect 6581 1231 6637 1240
rect 7829 1296 7885 1305
rect 7829 1231 7885 1240
rect 9077 1296 9133 1305
rect 9077 1231 9133 1240
rect 10325 1296 10381 1305
rect 10325 1231 10381 1240
rect 11573 1296 11629 1305
rect 11573 1231 11629 1240
rect 12821 1296 12877 1305
rect 12821 1231 12877 1240
rect 14069 1296 14125 1305
rect 14069 1231 14125 1240
rect 15317 1296 15373 1305
rect 15317 1231 15373 1240
rect 16565 1296 16621 1305
rect 16565 1231 16621 1240
rect 17813 1296 17869 1305
rect 17813 1231 17869 1240
rect 19061 1296 19117 1305
rect 19061 1231 19117 1240
rect 20309 1296 20365 1305
rect 20309 1231 20365 1240
rect 21557 1296 21613 1305
rect 21557 1231 21613 1240
rect 22805 1296 22861 1305
rect 22805 1231 22861 1240
rect 24053 1296 24109 1305
rect 24053 1231 24109 1240
rect 25301 1296 25357 1305
rect 25301 1231 25357 1240
rect 26549 1296 26605 1305
rect 26549 1231 26605 1240
rect 27797 1296 27853 1305
rect 27797 1231 27853 1240
rect 29045 1296 29101 1305
rect 29045 1231 29101 1240
rect 30293 1296 30349 1305
rect 30293 1231 30349 1240
rect 31541 1296 31597 1305
rect 31541 1231 31597 1240
rect 32789 1296 32845 1305
rect 32789 1231 32845 1240
rect 34037 1296 34093 1305
rect 34037 1231 34093 1240
rect 35285 1296 35341 1305
rect 35285 1231 35341 1240
rect 36533 1296 36589 1305
rect 36533 1231 36589 1240
rect 37781 1296 37837 1305
rect 37781 1231 37837 1240
rect 39029 1296 39085 1305
rect 39029 1231 39085 1240
rect 353 458 409 467
rect 353 393 409 402
rect 1601 458 1657 467
rect 1601 393 1657 402
rect 2849 458 2905 467
rect 2849 393 2905 402
rect 4097 458 4153 467
rect 4097 393 4153 402
rect 5345 458 5401 467
rect 5345 393 5401 402
rect 6593 458 6649 467
rect 6593 393 6649 402
rect 7841 458 7897 467
rect 7841 393 7897 402
rect 9089 458 9145 467
rect 9089 393 9145 402
rect 10337 458 10393 467
rect 10337 393 10393 402
rect 11585 458 11641 467
rect 11585 393 11641 402
rect 12833 458 12889 467
rect 12833 393 12889 402
rect 14081 458 14137 467
rect 14081 393 14137 402
rect 15329 458 15385 467
rect 15329 393 15385 402
rect 16577 458 16633 467
rect 16577 393 16633 402
rect 17825 458 17881 467
rect 17825 393 17881 402
rect 19073 458 19129 467
rect 19073 393 19129 402
rect 20321 458 20377 467
rect 20321 393 20377 402
rect 21569 458 21625 467
rect 21569 393 21625 402
rect 22817 458 22873 467
rect 22817 393 22873 402
rect 24065 458 24121 467
rect 24065 393 24121 402
rect 25313 458 25369 467
rect 25313 393 25369 402
rect 26561 458 26617 467
rect 26561 393 26617 402
rect 27809 458 27865 467
rect 27809 393 27865 402
rect 29057 458 29113 467
rect 29057 393 29113 402
rect 30305 458 30361 467
rect 30305 393 30361 402
rect 31553 458 31609 467
rect 31553 393 31609 402
rect 32801 458 32857 467
rect 32801 393 32857 402
rect 34049 458 34105 467
rect 34049 393 34105 402
rect 35297 458 35353 467
rect 35297 393 35353 402
rect 36545 458 36601 467
rect 36545 393 36601 402
rect 37793 458 37849 467
rect 37793 393 37849 402
rect 39041 458 39097 467
rect 39041 393 39097 402
rect 353 136 409 145
rect 353 71 409 80
rect 1601 136 1657 145
rect 1601 71 1657 80
rect 2849 136 2905 145
rect 2849 71 2905 80
rect 4097 136 4153 145
rect 4097 71 4153 80
rect 5345 136 5401 145
rect 5345 71 5401 80
rect 6593 136 6649 145
rect 6593 71 6649 80
rect 7841 136 7897 145
rect 7841 71 7897 80
rect 9089 136 9145 145
rect 9089 71 9145 80
rect 10337 136 10393 145
rect 10337 71 10393 80
rect 11585 136 11641 145
rect 11585 71 11641 80
rect 12833 136 12889 145
rect 12833 71 12889 80
rect 14081 136 14137 145
rect 14081 71 14137 80
rect 15329 136 15385 145
rect 15329 71 15385 80
rect 16577 136 16633 145
rect 16577 71 16633 80
rect 17825 136 17881 145
rect 17825 71 17881 80
rect 19073 136 19129 145
rect 19073 71 19129 80
rect 20321 136 20377 145
rect 20321 71 20377 80
rect 21569 136 21625 145
rect 21569 71 21625 80
rect 22817 136 22873 145
rect 22817 71 22873 80
rect 24065 136 24121 145
rect 24065 71 24121 80
rect 25313 136 25369 145
rect 25313 71 25369 80
rect 26561 136 26617 145
rect 26561 71 26617 80
rect 27809 136 27865 145
rect 27809 71 27865 80
rect 29057 136 29113 145
rect 29057 71 29113 80
rect 30305 136 30361 145
rect 30305 71 30361 80
rect 31553 136 31609 145
rect 31553 71 31609 80
rect 32801 136 32857 145
rect 32801 71 32857 80
rect 34049 136 34105 145
rect 34049 71 34105 80
rect 35297 136 35353 145
rect 35297 71 35353 80
rect 36545 136 36601 145
rect 36545 71 36601 80
rect 37793 136 37849 145
rect 37793 71 37849 80
rect 39041 136 39097 145
rect 39041 71 39097 80
<< via2 >>
rect 95 2220 151 2222
rect 95 2168 97 2220
rect 97 2168 149 2220
rect 149 2168 151 2220
rect 95 2166 151 2168
rect 1343 2220 1399 2222
rect 1343 2168 1345 2220
rect 1345 2168 1397 2220
rect 1397 2168 1399 2220
rect 1343 2166 1399 2168
rect 2591 2220 2647 2222
rect 2591 2168 2593 2220
rect 2593 2168 2645 2220
rect 2645 2168 2647 2220
rect 2591 2166 2647 2168
rect 3839 2220 3895 2222
rect 3839 2168 3841 2220
rect 3841 2168 3893 2220
rect 3893 2168 3895 2220
rect 3839 2166 3895 2168
rect 5087 2220 5143 2222
rect 5087 2168 5089 2220
rect 5089 2168 5141 2220
rect 5141 2168 5143 2220
rect 5087 2166 5143 2168
rect 6335 2220 6391 2222
rect 6335 2168 6337 2220
rect 6337 2168 6389 2220
rect 6389 2168 6391 2220
rect 6335 2166 6391 2168
rect 7583 2220 7639 2222
rect 7583 2168 7585 2220
rect 7585 2168 7637 2220
rect 7637 2168 7639 2220
rect 7583 2166 7639 2168
rect 8831 2220 8887 2222
rect 8831 2168 8833 2220
rect 8833 2168 8885 2220
rect 8885 2168 8887 2220
rect 8831 2166 8887 2168
rect 10079 2220 10135 2222
rect 10079 2168 10081 2220
rect 10081 2168 10133 2220
rect 10133 2168 10135 2220
rect 10079 2166 10135 2168
rect 11327 2220 11383 2222
rect 11327 2168 11329 2220
rect 11329 2168 11381 2220
rect 11381 2168 11383 2220
rect 11327 2166 11383 2168
rect 12575 2220 12631 2222
rect 12575 2168 12577 2220
rect 12577 2168 12629 2220
rect 12629 2168 12631 2220
rect 12575 2166 12631 2168
rect 13823 2220 13879 2222
rect 13823 2168 13825 2220
rect 13825 2168 13877 2220
rect 13877 2168 13879 2220
rect 13823 2166 13879 2168
rect 15071 2220 15127 2222
rect 15071 2168 15073 2220
rect 15073 2168 15125 2220
rect 15125 2168 15127 2220
rect 15071 2166 15127 2168
rect 16319 2220 16375 2222
rect 16319 2168 16321 2220
rect 16321 2168 16373 2220
rect 16373 2168 16375 2220
rect 16319 2166 16375 2168
rect 17567 2220 17623 2222
rect 17567 2168 17569 2220
rect 17569 2168 17621 2220
rect 17621 2168 17623 2220
rect 17567 2166 17623 2168
rect 18815 2220 18871 2222
rect 18815 2168 18817 2220
rect 18817 2168 18869 2220
rect 18869 2168 18871 2220
rect 18815 2166 18871 2168
rect 20063 2220 20119 2222
rect 20063 2168 20065 2220
rect 20065 2168 20117 2220
rect 20117 2168 20119 2220
rect 20063 2166 20119 2168
rect 21311 2220 21367 2222
rect 21311 2168 21313 2220
rect 21313 2168 21365 2220
rect 21365 2168 21367 2220
rect 21311 2166 21367 2168
rect 22559 2220 22615 2222
rect 22559 2168 22561 2220
rect 22561 2168 22613 2220
rect 22613 2168 22615 2220
rect 22559 2166 22615 2168
rect 23807 2220 23863 2222
rect 23807 2168 23809 2220
rect 23809 2168 23861 2220
rect 23861 2168 23863 2220
rect 23807 2166 23863 2168
rect 25055 2220 25111 2222
rect 25055 2168 25057 2220
rect 25057 2168 25109 2220
rect 25109 2168 25111 2220
rect 25055 2166 25111 2168
rect 26303 2220 26359 2222
rect 26303 2168 26305 2220
rect 26305 2168 26357 2220
rect 26357 2168 26359 2220
rect 26303 2166 26359 2168
rect 27551 2220 27607 2222
rect 27551 2168 27553 2220
rect 27553 2168 27605 2220
rect 27605 2168 27607 2220
rect 27551 2166 27607 2168
rect 28799 2220 28855 2222
rect 28799 2168 28801 2220
rect 28801 2168 28853 2220
rect 28853 2168 28855 2220
rect 28799 2166 28855 2168
rect 30047 2220 30103 2222
rect 30047 2168 30049 2220
rect 30049 2168 30101 2220
rect 30101 2168 30103 2220
rect 30047 2166 30103 2168
rect 31295 2220 31351 2222
rect 31295 2168 31297 2220
rect 31297 2168 31349 2220
rect 31349 2168 31351 2220
rect 31295 2166 31351 2168
rect 32543 2220 32599 2222
rect 32543 2168 32545 2220
rect 32545 2168 32597 2220
rect 32597 2168 32599 2220
rect 32543 2166 32599 2168
rect 33791 2220 33847 2222
rect 33791 2168 33793 2220
rect 33793 2168 33845 2220
rect 33845 2168 33847 2220
rect 33791 2166 33847 2168
rect 35039 2220 35095 2222
rect 35039 2168 35041 2220
rect 35041 2168 35093 2220
rect 35093 2168 35095 2220
rect 35039 2166 35095 2168
rect 36287 2220 36343 2222
rect 36287 2168 36289 2220
rect 36289 2168 36341 2220
rect 36341 2168 36343 2220
rect 36287 2166 36343 2168
rect 37535 2220 37591 2222
rect 37535 2168 37537 2220
rect 37537 2168 37589 2220
rect 37589 2168 37591 2220
rect 37535 2166 37591 2168
rect 38783 2220 38839 2222
rect 38783 2168 38785 2220
rect 38785 2168 38837 2220
rect 38837 2168 38839 2220
rect 38783 2166 38839 2168
rect 423 2068 479 2070
rect 423 2016 425 2068
rect 425 2016 477 2068
rect 477 2016 479 2068
rect 423 2014 479 2016
rect 1671 2068 1727 2070
rect 1671 2016 1673 2068
rect 1673 2016 1725 2068
rect 1725 2016 1727 2068
rect 1671 2014 1727 2016
rect 2919 2068 2975 2070
rect 2919 2016 2921 2068
rect 2921 2016 2973 2068
rect 2973 2016 2975 2068
rect 2919 2014 2975 2016
rect 4167 2068 4223 2070
rect 4167 2016 4169 2068
rect 4169 2016 4221 2068
rect 4221 2016 4223 2068
rect 4167 2014 4223 2016
rect 5415 2068 5471 2070
rect 5415 2016 5417 2068
rect 5417 2016 5469 2068
rect 5469 2016 5471 2068
rect 5415 2014 5471 2016
rect 6663 2068 6719 2070
rect 6663 2016 6665 2068
rect 6665 2016 6717 2068
rect 6717 2016 6719 2068
rect 6663 2014 6719 2016
rect 7911 2068 7967 2070
rect 7911 2016 7913 2068
rect 7913 2016 7965 2068
rect 7965 2016 7967 2068
rect 7911 2014 7967 2016
rect 9159 2068 9215 2070
rect 9159 2016 9161 2068
rect 9161 2016 9213 2068
rect 9213 2016 9215 2068
rect 9159 2014 9215 2016
rect 10407 2068 10463 2070
rect 10407 2016 10409 2068
rect 10409 2016 10461 2068
rect 10461 2016 10463 2068
rect 10407 2014 10463 2016
rect 11655 2068 11711 2070
rect 11655 2016 11657 2068
rect 11657 2016 11709 2068
rect 11709 2016 11711 2068
rect 11655 2014 11711 2016
rect 12903 2068 12959 2070
rect 12903 2016 12905 2068
rect 12905 2016 12957 2068
rect 12957 2016 12959 2068
rect 12903 2014 12959 2016
rect 14151 2068 14207 2070
rect 14151 2016 14153 2068
rect 14153 2016 14205 2068
rect 14205 2016 14207 2068
rect 14151 2014 14207 2016
rect 15399 2068 15455 2070
rect 15399 2016 15401 2068
rect 15401 2016 15453 2068
rect 15453 2016 15455 2068
rect 15399 2014 15455 2016
rect 16647 2068 16703 2070
rect 16647 2016 16649 2068
rect 16649 2016 16701 2068
rect 16701 2016 16703 2068
rect 16647 2014 16703 2016
rect 17895 2068 17951 2070
rect 17895 2016 17897 2068
rect 17897 2016 17949 2068
rect 17949 2016 17951 2068
rect 17895 2014 17951 2016
rect 19143 2068 19199 2070
rect 19143 2016 19145 2068
rect 19145 2016 19197 2068
rect 19197 2016 19199 2068
rect 19143 2014 19199 2016
rect 20391 2068 20447 2070
rect 20391 2016 20393 2068
rect 20393 2016 20445 2068
rect 20445 2016 20447 2068
rect 20391 2014 20447 2016
rect 21639 2068 21695 2070
rect 21639 2016 21641 2068
rect 21641 2016 21693 2068
rect 21693 2016 21695 2068
rect 21639 2014 21695 2016
rect 22887 2068 22943 2070
rect 22887 2016 22889 2068
rect 22889 2016 22941 2068
rect 22941 2016 22943 2068
rect 22887 2014 22943 2016
rect 24135 2068 24191 2070
rect 24135 2016 24137 2068
rect 24137 2016 24189 2068
rect 24189 2016 24191 2068
rect 24135 2014 24191 2016
rect 25383 2068 25439 2070
rect 25383 2016 25385 2068
rect 25385 2016 25437 2068
rect 25437 2016 25439 2068
rect 25383 2014 25439 2016
rect 26631 2068 26687 2070
rect 26631 2016 26633 2068
rect 26633 2016 26685 2068
rect 26685 2016 26687 2068
rect 26631 2014 26687 2016
rect 27879 2068 27935 2070
rect 27879 2016 27881 2068
rect 27881 2016 27933 2068
rect 27933 2016 27935 2068
rect 27879 2014 27935 2016
rect 29127 2068 29183 2070
rect 29127 2016 29129 2068
rect 29129 2016 29181 2068
rect 29181 2016 29183 2068
rect 29127 2014 29183 2016
rect 30375 2068 30431 2070
rect 30375 2016 30377 2068
rect 30377 2016 30429 2068
rect 30429 2016 30431 2068
rect 30375 2014 30431 2016
rect 31623 2068 31679 2070
rect 31623 2016 31625 2068
rect 31625 2016 31677 2068
rect 31677 2016 31679 2068
rect 31623 2014 31679 2016
rect 32871 2068 32927 2070
rect 32871 2016 32873 2068
rect 32873 2016 32925 2068
rect 32925 2016 32927 2068
rect 32871 2014 32927 2016
rect 34119 2068 34175 2070
rect 34119 2016 34121 2068
rect 34121 2016 34173 2068
rect 34173 2016 34175 2068
rect 34119 2014 34175 2016
rect 35367 2068 35423 2070
rect 35367 2016 35369 2068
rect 35369 2016 35421 2068
rect 35421 2016 35423 2068
rect 35367 2014 35423 2016
rect 36615 2068 36671 2070
rect 36615 2016 36617 2068
rect 36617 2016 36669 2068
rect 36669 2016 36671 2068
rect 36615 2014 36671 2016
rect 37863 2068 37919 2070
rect 37863 2016 37865 2068
rect 37865 2016 37917 2068
rect 37917 2016 37919 2068
rect 37863 2014 37919 2016
rect 39111 2068 39167 2070
rect 39111 2016 39113 2068
rect 39113 2016 39165 2068
rect 39165 2016 39167 2068
rect 39111 2014 39167 2016
rect 341 1294 397 1296
rect 341 1242 343 1294
rect 343 1242 395 1294
rect 395 1242 397 1294
rect 341 1240 397 1242
rect 1589 1294 1645 1296
rect 1589 1242 1591 1294
rect 1591 1242 1643 1294
rect 1643 1242 1645 1294
rect 1589 1240 1645 1242
rect 2837 1294 2893 1296
rect 2837 1242 2839 1294
rect 2839 1242 2891 1294
rect 2891 1242 2893 1294
rect 2837 1240 2893 1242
rect 4085 1294 4141 1296
rect 4085 1242 4087 1294
rect 4087 1242 4139 1294
rect 4139 1242 4141 1294
rect 4085 1240 4141 1242
rect 5333 1294 5389 1296
rect 5333 1242 5335 1294
rect 5335 1242 5387 1294
rect 5387 1242 5389 1294
rect 5333 1240 5389 1242
rect 6581 1294 6637 1296
rect 6581 1242 6583 1294
rect 6583 1242 6635 1294
rect 6635 1242 6637 1294
rect 6581 1240 6637 1242
rect 7829 1294 7885 1296
rect 7829 1242 7831 1294
rect 7831 1242 7883 1294
rect 7883 1242 7885 1294
rect 7829 1240 7885 1242
rect 9077 1294 9133 1296
rect 9077 1242 9079 1294
rect 9079 1242 9131 1294
rect 9131 1242 9133 1294
rect 9077 1240 9133 1242
rect 10325 1294 10381 1296
rect 10325 1242 10327 1294
rect 10327 1242 10379 1294
rect 10379 1242 10381 1294
rect 10325 1240 10381 1242
rect 11573 1294 11629 1296
rect 11573 1242 11575 1294
rect 11575 1242 11627 1294
rect 11627 1242 11629 1294
rect 11573 1240 11629 1242
rect 12821 1294 12877 1296
rect 12821 1242 12823 1294
rect 12823 1242 12875 1294
rect 12875 1242 12877 1294
rect 12821 1240 12877 1242
rect 14069 1294 14125 1296
rect 14069 1242 14071 1294
rect 14071 1242 14123 1294
rect 14123 1242 14125 1294
rect 14069 1240 14125 1242
rect 15317 1294 15373 1296
rect 15317 1242 15319 1294
rect 15319 1242 15371 1294
rect 15371 1242 15373 1294
rect 15317 1240 15373 1242
rect 16565 1294 16621 1296
rect 16565 1242 16567 1294
rect 16567 1242 16619 1294
rect 16619 1242 16621 1294
rect 16565 1240 16621 1242
rect 17813 1294 17869 1296
rect 17813 1242 17815 1294
rect 17815 1242 17867 1294
rect 17867 1242 17869 1294
rect 17813 1240 17869 1242
rect 19061 1294 19117 1296
rect 19061 1242 19063 1294
rect 19063 1242 19115 1294
rect 19115 1242 19117 1294
rect 19061 1240 19117 1242
rect 20309 1294 20365 1296
rect 20309 1242 20311 1294
rect 20311 1242 20363 1294
rect 20363 1242 20365 1294
rect 20309 1240 20365 1242
rect 21557 1294 21613 1296
rect 21557 1242 21559 1294
rect 21559 1242 21611 1294
rect 21611 1242 21613 1294
rect 21557 1240 21613 1242
rect 22805 1294 22861 1296
rect 22805 1242 22807 1294
rect 22807 1242 22859 1294
rect 22859 1242 22861 1294
rect 22805 1240 22861 1242
rect 24053 1294 24109 1296
rect 24053 1242 24055 1294
rect 24055 1242 24107 1294
rect 24107 1242 24109 1294
rect 24053 1240 24109 1242
rect 25301 1294 25357 1296
rect 25301 1242 25303 1294
rect 25303 1242 25355 1294
rect 25355 1242 25357 1294
rect 25301 1240 25357 1242
rect 26549 1294 26605 1296
rect 26549 1242 26551 1294
rect 26551 1242 26603 1294
rect 26603 1242 26605 1294
rect 26549 1240 26605 1242
rect 27797 1294 27853 1296
rect 27797 1242 27799 1294
rect 27799 1242 27851 1294
rect 27851 1242 27853 1294
rect 27797 1240 27853 1242
rect 29045 1294 29101 1296
rect 29045 1242 29047 1294
rect 29047 1242 29099 1294
rect 29099 1242 29101 1294
rect 29045 1240 29101 1242
rect 30293 1294 30349 1296
rect 30293 1242 30295 1294
rect 30295 1242 30347 1294
rect 30347 1242 30349 1294
rect 30293 1240 30349 1242
rect 31541 1294 31597 1296
rect 31541 1242 31543 1294
rect 31543 1242 31595 1294
rect 31595 1242 31597 1294
rect 31541 1240 31597 1242
rect 32789 1294 32845 1296
rect 32789 1242 32791 1294
rect 32791 1242 32843 1294
rect 32843 1242 32845 1294
rect 32789 1240 32845 1242
rect 34037 1294 34093 1296
rect 34037 1242 34039 1294
rect 34039 1242 34091 1294
rect 34091 1242 34093 1294
rect 34037 1240 34093 1242
rect 35285 1294 35341 1296
rect 35285 1242 35287 1294
rect 35287 1242 35339 1294
rect 35339 1242 35341 1294
rect 35285 1240 35341 1242
rect 36533 1294 36589 1296
rect 36533 1242 36535 1294
rect 36535 1242 36587 1294
rect 36587 1242 36589 1294
rect 36533 1240 36589 1242
rect 37781 1294 37837 1296
rect 37781 1242 37783 1294
rect 37783 1242 37835 1294
rect 37835 1242 37837 1294
rect 37781 1240 37837 1242
rect 39029 1294 39085 1296
rect 39029 1242 39031 1294
rect 39031 1242 39083 1294
rect 39083 1242 39085 1294
rect 39029 1240 39085 1242
rect 353 456 409 458
rect 353 404 355 456
rect 355 404 407 456
rect 407 404 409 456
rect 353 402 409 404
rect 1601 456 1657 458
rect 1601 404 1603 456
rect 1603 404 1655 456
rect 1655 404 1657 456
rect 1601 402 1657 404
rect 2849 456 2905 458
rect 2849 404 2851 456
rect 2851 404 2903 456
rect 2903 404 2905 456
rect 2849 402 2905 404
rect 4097 456 4153 458
rect 4097 404 4099 456
rect 4099 404 4151 456
rect 4151 404 4153 456
rect 4097 402 4153 404
rect 5345 456 5401 458
rect 5345 404 5347 456
rect 5347 404 5399 456
rect 5399 404 5401 456
rect 5345 402 5401 404
rect 6593 456 6649 458
rect 6593 404 6595 456
rect 6595 404 6647 456
rect 6647 404 6649 456
rect 6593 402 6649 404
rect 7841 456 7897 458
rect 7841 404 7843 456
rect 7843 404 7895 456
rect 7895 404 7897 456
rect 7841 402 7897 404
rect 9089 456 9145 458
rect 9089 404 9091 456
rect 9091 404 9143 456
rect 9143 404 9145 456
rect 9089 402 9145 404
rect 10337 456 10393 458
rect 10337 404 10339 456
rect 10339 404 10391 456
rect 10391 404 10393 456
rect 10337 402 10393 404
rect 11585 456 11641 458
rect 11585 404 11587 456
rect 11587 404 11639 456
rect 11639 404 11641 456
rect 11585 402 11641 404
rect 12833 456 12889 458
rect 12833 404 12835 456
rect 12835 404 12887 456
rect 12887 404 12889 456
rect 12833 402 12889 404
rect 14081 456 14137 458
rect 14081 404 14083 456
rect 14083 404 14135 456
rect 14135 404 14137 456
rect 14081 402 14137 404
rect 15329 456 15385 458
rect 15329 404 15331 456
rect 15331 404 15383 456
rect 15383 404 15385 456
rect 15329 402 15385 404
rect 16577 456 16633 458
rect 16577 404 16579 456
rect 16579 404 16631 456
rect 16631 404 16633 456
rect 16577 402 16633 404
rect 17825 456 17881 458
rect 17825 404 17827 456
rect 17827 404 17879 456
rect 17879 404 17881 456
rect 17825 402 17881 404
rect 19073 456 19129 458
rect 19073 404 19075 456
rect 19075 404 19127 456
rect 19127 404 19129 456
rect 19073 402 19129 404
rect 20321 456 20377 458
rect 20321 404 20323 456
rect 20323 404 20375 456
rect 20375 404 20377 456
rect 20321 402 20377 404
rect 21569 456 21625 458
rect 21569 404 21571 456
rect 21571 404 21623 456
rect 21623 404 21625 456
rect 21569 402 21625 404
rect 22817 456 22873 458
rect 22817 404 22819 456
rect 22819 404 22871 456
rect 22871 404 22873 456
rect 22817 402 22873 404
rect 24065 456 24121 458
rect 24065 404 24067 456
rect 24067 404 24119 456
rect 24119 404 24121 456
rect 24065 402 24121 404
rect 25313 456 25369 458
rect 25313 404 25315 456
rect 25315 404 25367 456
rect 25367 404 25369 456
rect 25313 402 25369 404
rect 26561 456 26617 458
rect 26561 404 26563 456
rect 26563 404 26615 456
rect 26615 404 26617 456
rect 26561 402 26617 404
rect 27809 456 27865 458
rect 27809 404 27811 456
rect 27811 404 27863 456
rect 27863 404 27865 456
rect 27809 402 27865 404
rect 29057 456 29113 458
rect 29057 404 29059 456
rect 29059 404 29111 456
rect 29111 404 29113 456
rect 29057 402 29113 404
rect 30305 456 30361 458
rect 30305 404 30307 456
rect 30307 404 30359 456
rect 30359 404 30361 456
rect 30305 402 30361 404
rect 31553 456 31609 458
rect 31553 404 31555 456
rect 31555 404 31607 456
rect 31607 404 31609 456
rect 31553 402 31609 404
rect 32801 456 32857 458
rect 32801 404 32803 456
rect 32803 404 32855 456
rect 32855 404 32857 456
rect 32801 402 32857 404
rect 34049 456 34105 458
rect 34049 404 34051 456
rect 34051 404 34103 456
rect 34103 404 34105 456
rect 34049 402 34105 404
rect 35297 456 35353 458
rect 35297 404 35299 456
rect 35299 404 35351 456
rect 35351 404 35353 456
rect 35297 402 35353 404
rect 36545 456 36601 458
rect 36545 404 36547 456
rect 36547 404 36599 456
rect 36599 404 36601 456
rect 36545 402 36601 404
rect 37793 456 37849 458
rect 37793 404 37795 456
rect 37795 404 37847 456
rect 37847 404 37849 456
rect 37793 402 37849 404
rect 39041 456 39097 458
rect 39041 404 39043 456
rect 39043 404 39095 456
rect 39095 404 39097 456
rect 39041 402 39097 404
rect 353 134 409 136
rect 353 82 355 134
rect 355 82 407 134
rect 407 82 409 134
rect 353 80 409 82
rect 1601 134 1657 136
rect 1601 82 1603 134
rect 1603 82 1655 134
rect 1655 82 1657 134
rect 1601 80 1657 82
rect 2849 134 2905 136
rect 2849 82 2851 134
rect 2851 82 2903 134
rect 2903 82 2905 134
rect 2849 80 2905 82
rect 4097 134 4153 136
rect 4097 82 4099 134
rect 4099 82 4151 134
rect 4151 82 4153 134
rect 4097 80 4153 82
rect 5345 134 5401 136
rect 5345 82 5347 134
rect 5347 82 5399 134
rect 5399 82 5401 134
rect 5345 80 5401 82
rect 6593 134 6649 136
rect 6593 82 6595 134
rect 6595 82 6647 134
rect 6647 82 6649 134
rect 6593 80 6649 82
rect 7841 134 7897 136
rect 7841 82 7843 134
rect 7843 82 7895 134
rect 7895 82 7897 134
rect 7841 80 7897 82
rect 9089 134 9145 136
rect 9089 82 9091 134
rect 9091 82 9143 134
rect 9143 82 9145 134
rect 9089 80 9145 82
rect 10337 134 10393 136
rect 10337 82 10339 134
rect 10339 82 10391 134
rect 10391 82 10393 134
rect 10337 80 10393 82
rect 11585 134 11641 136
rect 11585 82 11587 134
rect 11587 82 11639 134
rect 11639 82 11641 134
rect 11585 80 11641 82
rect 12833 134 12889 136
rect 12833 82 12835 134
rect 12835 82 12887 134
rect 12887 82 12889 134
rect 12833 80 12889 82
rect 14081 134 14137 136
rect 14081 82 14083 134
rect 14083 82 14135 134
rect 14135 82 14137 134
rect 14081 80 14137 82
rect 15329 134 15385 136
rect 15329 82 15331 134
rect 15331 82 15383 134
rect 15383 82 15385 134
rect 15329 80 15385 82
rect 16577 134 16633 136
rect 16577 82 16579 134
rect 16579 82 16631 134
rect 16631 82 16633 134
rect 16577 80 16633 82
rect 17825 134 17881 136
rect 17825 82 17827 134
rect 17827 82 17879 134
rect 17879 82 17881 134
rect 17825 80 17881 82
rect 19073 134 19129 136
rect 19073 82 19075 134
rect 19075 82 19127 134
rect 19127 82 19129 134
rect 19073 80 19129 82
rect 20321 134 20377 136
rect 20321 82 20323 134
rect 20323 82 20375 134
rect 20375 82 20377 134
rect 20321 80 20377 82
rect 21569 134 21625 136
rect 21569 82 21571 134
rect 21571 82 21623 134
rect 21623 82 21625 134
rect 21569 80 21625 82
rect 22817 134 22873 136
rect 22817 82 22819 134
rect 22819 82 22871 134
rect 22871 82 22873 134
rect 22817 80 22873 82
rect 24065 134 24121 136
rect 24065 82 24067 134
rect 24067 82 24119 134
rect 24119 82 24121 134
rect 24065 80 24121 82
rect 25313 134 25369 136
rect 25313 82 25315 134
rect 25315 82 25367 134
rect 25367 82 25369 134
rect 25313 80 25369 82
rect 26561 134 26617 136
rect 26561 82 26563 134
rect 26563 82 26615 134
rect 26615 82 26617 134
rect 26561 80 26617 82
rect 27809 134 27865 136
rect 27809 82 27811 134
rect 27811 82 27863 134
rect 27863 82 27865 134
rect 27809 80 27865 82
rect 29057 134 29113 136
rect 29057 82 29059 134
rect 29059 82 29111 134
rect 29111 82 29113 134
rect 29057 80 29113 82
rect 30305 134 30361 136
rect 30305 82 30307 134
rect 30307 82 30359 134
rect 30359 82 30361 134
rect 30305 80 30361 82
rect 31553 134 31609 136
rect 31553 82 31555 134
rect 31555 82 31607 134
rect 31607 82 31609 134
rect 31553 80 31609 82
rect 32801 134 32857 136
rect 32801 82 32803 134
rect 32803 82 32855 134
rect 32855 82 32857 134
rect 32801 80 32857 82
rect 34049 134 34105 136
rect 34049 82 34051 134
rect 34051 82 34103 134
rect 34103 82 34105 134
rect 34049 80 34105 82
rect 35297 134 35353 136
rect 35297 82 35299 134
rect 35299 82 35351 134
rect 35351 82 35353 134
rect 35297 80 35353 82
rect 36545 134 36601 136
rect 36545 82 36547 134
rect 36547 82 36599 134
rect 36599 82 36601 134
rect 36545 80 36601 82
rect 37793 134 37849 136
rect 37793 82 37795 134
rect 37795 82 37847 134
rect 37847 82 37849 134
rect 37793 80 37849 82
rect 39041 134 39097 136
rect 39041 82 39043 134
rect 39043 82 39095 134
rect 39095 82 39097 134
rect 39041 80 39097 82
<< metal3 >>
rect 90 2224 156 2227
rect 1338 2224 1404 2227
rect 2586 2224 2652 2227
rect 3834 2224 3900 2227
rect 5082 2224 5148 2227
rect 6330 2224 6396 2227
rect 7578 2224 7644 2227
rect 8826 2224 8892 2227
rect 10074 2224 10140 2227
rect 11322 2224 11388 2227
rect 12570 2224 12636 2227
rect 13818 2224 13884 2227
rect 15066 2224 15132 2227
rect 16314 2224 16380 2227
rect 17562 2224 17628 2227
rect 18810 2224 18876 2227
rect 20058 2224 20124 2227
rect 21306 2224 21372 2227
rect 22554 2224 22620 2227
rect 23802 2224 23868 2227
rect 25050 2224 25116 2227
rect 26298 2224 26364 2227
rect 27546 2224 27612 2227
rect 28794 2224 28860 2227
rect 30042 2224 30108 2227
rect 31290 2224 31356 2227
rect 32538 2224 32604 2227
rect 33786 2224 33852 2227
rect 35034 2224 35100 2227
rect 36282 2224 36348 2227
rect 37530 2224 37596 2227
rect 38778 2224 38844 2227
rect 0 2222 39936 2224
rect 0 2166 95 2222
rect 151 2166 1343 2222
rect 1399 2166 2591 2222
rect 2647 2166 3839 2222
rect 3895 2166 5087 2222
rect 5143 2166 6335 2222
rect 6391 2166 7583 2222
rect 7639 2166 8831 2222
rect 8887 2166 10079 2222
rect 10135 2166 11327 2222
rect 11383 2166 12575 2222
rect 12631 2166 13823 2222
rect 13879 2166 15071 2222
rect 15127 2166 16319 2222
rect 16375 2166 17567 2222
rect 17623 2166 18815 2222
rect 18871 2166 20063 2222
rect 20119 2166 21311 2222
rect 21367 2166 22559 2222
rect 22615 2166 23807 2222
rect 23863 2166 25055 2222
rect 25111 2166 26303 2222
rect 26359 2166 27551 2222
rect 27607 2166 28799 2222
rect 28855 2166 30047 2222
rect 30103 2166 31295 2222
rect 31351 2166 32543 2222
rect 32599 2166 33791 2222
rect 33847 2166 35039 2222
rect 35095 2166 36287 2222
rect 36343 2166 37535 2222
rect 37591 2166 38783 2222
rect 38839 2166 39936 2222
rect 0 2164 39936 2166
rect 90 2161 156 2164
rect 1338 2161 1404 2164
rect 2586 2161 2652 2164
rect 3834 2161 3900 2164
rect 5082 2161 5148 2164
rect 6330 2161 6396 2164
rect 7578 2161 7644 2164
rect 8826 2161 8892 2164
rect 10074 2161 10140 2164
rect 11322 2161 11388 2164
rect 12570 2161 12636 2164
rect 13818 2161 13884 2164
rect 15066 2161 15132 2164
rect 16314 2161 16380 2164
rect 17562 2161 17628 2164
rect 18810 2161 18876 2164
rect 20058 2161 20124 2164
rect 21306 2161 21372 2164
rect 22554 2161 22620 2164
rect 23802 2161 23868 2164
rect 25050 2161 25116 2164
rect 26298 2161 26364 2164
rect 27546 2161 27612 2164
rect 28794 2161 28860 2164
rect 30042 2161 30108 2164
rect 31290 2161 31356 2164
rect 32538 2161 32604 2164
rect 33786 2161 33852 2164
rect 35034 2161 35100 2164
rect 36282 2161 36348 2164
rect 37530 2161 37596 2164
rect 38778 2161 38844 2164
rect 402 2070 500 2091
rect 402 2014 423 2070
rect 479 2014 500 2070
rect 402 1993 500 2014
rect 1650 2070 1748 2091
rect 1650 2014 1671 2070
rect 1727 2014 1748 2070
rect 1650 1993 1748 2014
rect 2898 2070 2996 2091
rect 2898 2014 2919 2070
rect 2975 2014 2996 2070
rect 2898 1993 2996 2014
rect 4146 2070 4244 2091
rect 4146 2014 4167 2070
rect 4223 2014 4244 2070
rect 4146 1993 4244 2014
rect 5394 2070 5492 2091
rect 5394 2014 5415 2070
rect 5471 2014 5492 2070
rect 5394 1993 5492 2014
rect 6642 2070 6740 2091
rect 6642 2014 6663 2070
rect 6719 2014 6740 2070
rect 6642 1993 6740 2014
rect 7890 2070 7988 2091
rect 7890 2014 7911 2070
rect 7967 2014 7988 2070
rect 7890 1993 7988 2014
rect 9138 2070 9236 2091
rect 9138 2014 9159 2070
rect 9215 2014 9236 2070
rect 9138 1993 9236 2014
rect 10386 2070 10484 2091
rect 10386 2014 10407 2070
rect 10463 2014 10484 2070
rect 10386 1993 10484 2014
rect 11634 2070 11732 2091
rect 11634 2014 11655 2070
rect 11711 2014 11732 2070
rect 11634 1993 11732 2014
rect 12882 2070 12980 2091
rect 12882 2014 12903 2070
rect 12959 2014 12980 2070
rect 12882 1993 12980 2014
rect 14130 2070 14228 2091
rect 14130 2014 14151 2070
rect 14207 2014 14228 2070
rect 14130 1993 14228 2014
rect 15378 2070 15476 2091
rect 15378 2014 15399 2070
rect 15455 2014 15476 2070
rect 15378 1993 15476 2014
rect 16626 2070 16724 2091
rect 16626 2014 16647 2070
rect 16703 2014 16724 2070
rect 16626 1993 16724 2014
rect 17874 2070 17972 2091
rect 17874 2014 17895 2070
rect 17951 2014 17972 2070
rect 17874 1993 17972 2014
rect 19122 2070 19220 2091
rect 19122 2014 19143 2070
rect 19199 2014 19220 2070
rect 19122 1993 19220 2014
rect 20370 2070 20468 2091
rect 20370 2014 20391 2070
rect 20447 2014 20468 2070
rect 20370 1993 20468 2014
rect 21618 2070 21716 2091
rect 21618 2014 21639 2070
rect 21695 2014 21716 2070
rect 21618 1993 21716 2014
rect 22866 2070 22964 2091
rect 22866 2014 22887 2070
rect 22943 2014 22964 2070
rect 22866 1993 22964 2014
rect 24114 2070 24212 2091
rect 24114 2014 24135 2070
rect 24191 2014 24212 2070
rect 24114 1993 24212 2014
rect 25362 2070 25460 2091
rect 25362 2014 25383 2070
rect 25439 2014 25460 2070
rect 25362 1993 25460 2014
rect 26610 2070 26708 2091
rect 26610 2014 26631 2070
rect 26687 2014 26708 2070
rect 26610 1993 26708 2014
rect 27858 2070 27956 2091
rect 27858 2014 27879 2070
rect 27935 2014 27956 2070
rect 27858 1993 27956 2014
rect 29106 2070 29204 2091
rect 29106 2014 29127 2070
rect 29183 2014 29204 2070
rect 29106 1993 29204 2014
rect 30354 2070 30452 2091
rect 30354 2014 30375 2070
rect 30431 2014 30452 2070
rect 30354 1993 30452 2014
rect 31602 2070 31700 2091
rect 31602 2014 31623 2070
rect 31679 2014 31700 2070
rect 31602 1993 31700 2014
rect 32850 2070 32948 2091
rect 32850 2014 32871 2070
rect 32927 2014 32948 2070
rect 32850 1993 32948 2014
rect 34098 2070 34196 2091
rect 34098 2014 34119 2070
rect 34175 2014 34196 2070
rect 34098 1993 34196 2014
rect 35346 2070 35444 2091
rect 35346 2014 35367 2070
rect 35423 2014 35444 2070
rect 35346 1993 35444 2014
rect 36594 2070 36692 2091
rect 36594 2014 36615 2070
rect 36671 2014 36692 2070
rect 36594 1993 36692 2014
rect 37842 2070 37940 2091
rect 37842 2014 37863 2070
rect 37919 2014 37940 2070
rect 37842 1993 37940 2014
rect 39090 2070 39188 2091
rect 39090 2014 39111 2070
rect 39167 2014 39188 2070
rect 39090 1993 39188 2014
rect 320 1296 418 1317
rect 320 1240 341 1296
rect 397 1240 418 1296
rect 320 1219 418 1240
rect 1568 1296 1666 1317
rect 1568 1240 1589 1296
rect 1645 1240 1666 1296
rect 1568 1219 1666 1240
rect 2816 1296 2914 1317
rect 2816 1240 2837 1296
rect 2893 1240 2914 1296
rect 2816 1219 2914 1240
rect 4064 1296 4162 1317
rect 4064 1240 4085 1296
rect 4141 1240 4162 1296
rect 4064 1219 4162 1240
rect 5312 1296 5410 1317
rect 5312 1240 5333 1296
rect 5389 1240 5410 1296
rect 5312 1219 5410 1240
rect 6560 1296 6658 1317
rect 6560 1240 6581 1296
rect 6637 1240 6658 1296
rect 6560 1219 6658 1240
rect 7808 1296 7906 1317
rect 7808 1240 7829 1296
rect 7885 1240 7906 1296
rect 7808 1219 7906 1240
rect 9056 1296 9154 1317
rect 9056 1240 9077 1296
rect 9133 1240 9154 1296
rect 9056 1219 9154 1240
rect 10304 1296 10402 1317
rect 10304 1240 10325 1296
rect 10381 1240 10402 1296
rect 10304 1219 10402 1240
rect 11552 1296 11650 1317
rect 11552 1240 11573 1296
rect 11629 1240 11650 1296
rect 11552 1219 11650 1240
rect 12800 1296 12898 1317
rect 12800 1240 12821 1296
rect 12877 1240 12898 1296
rect 12800 1219 12898 1240
rect 14048 1296 14146 1317
rect 14048 1240 14069 1296
rect 14125 1240 14146 1296
rect 14048 1219 14146 1240
rect 15296 1296 15394 1317
rect 15296 1240 15317 1296
rect 15373 1240 15394 1296
rect 15296 1219 15394 1240
rect 16544 1296 16642 1317
rect 16544 1240 16565 1296
rect 16621 1240 16642 1296
rect 16544 1219 16642 1240
rect 17792 1296 17890 1317
rect 17792 1240 17813 1296
rect 17869 1240 17890 1296
rect 17792 1219 17890 1240
rect 19040 1296 19138 1317
rect 19040 1240 19061 1296
rect 19117 1240 19138 1296
rect 19040 1219 19138 1240
rect 20288 1296 20386 1317
rect 20288 1240 20309 1296
rect 20365 1240 20386 1296
rect 20288 1219 20386 1240
rect 21536 1296 21634 1317
rect 21536 1240 21557 1296
rect 21613 1240 21634 1296
rect 21536 1219 21634 1240
rect 22784 1296 22882 1317
rect 22784 1240 22805 1296
rect 22861 1240 22882 1296
rect 22784 1219 22882 1240
rect 24032 1296 24130 1317
rect 24032 1240 24053 1296
rect 24109 1240 24130 1296
rect 24032 1219 24130 1240
rect 25280 1296 25378 1317
rect 25280 1240 25301 1296
rect 25357 1240 25378 1296
rect 25280 1219 25378 1240
rect 26528 1296 26626 1317
rect 26528 1240 26549 1296
rect 26605 1240 26626 1296
rect 26528 1219 26626 1240
rect 27776 1296 27874 1317
rect 27776 1240 27797 1296
rect 27853 1240 27874 1296
rect 27776 1219 27874 1240
rect 29024 1296 29122 1317
rect 29024 1240 29045 1296
rect 29101 1240 29122 1296
rect 29024 1219 29122 1240
rect 30272 1296 30370 1317
rect 30272 1240 30293 1296
rect 30349 1240 30370 1296
rect 30272 1219 30370 1240
rect 31520 1296 31618 1317
rect 31520 1240 31541 1296
rect 31597 1240 31618 1296
rect 31520 1219 31618 1240
rect 32768 1296 32866 1317
rect 32768 1240 32789 1296
rect 32845 1240 32866 1296
rect 32768 1219 32866 1240
rect 34016 1296 34114 1317
rect 34016 1240 34037 1296
rect 34093 1240 34114 1296
rect 34016 1219 34114 1240
rect 35264 1296 35362 1317
rect 35264 1240 35285 1296
rect 35341 1240 35362 1296
rect 35264 1219 35362 1240
rect 36512 1296 36610 1317
rect 36512 1240 36533 1296
rect 36589 1240 36610 1296
rect 36512 1219 36610 1240
rect 37760 1296 37858 1317
rect 37760 1240 37781 1296
rect 37837 1240 37858 1296
rect 37760 1219 37858 1240
rect 39008 1296 39106 1317
rect 39008 1240 39029 1296
rect 39085 1240 39106 1296
rect 39008 1219 39106 1240
rect 332 458 430 479
rect 332 402 353 458
rect 409 402 430 458
rect 332 381 430 402
rect 1580 458 1678 479
rect 1580 402 1601 458
rect 1657 402 1678 458
rect 1580 381 1678 402
rect 2828 458 2926 479
rect 2828 402 2849 458
rect 2905 402 2926 458
rect 2828 381 2926 402
rect 4076 458 4174 479
rect 4076 402 4097 458
rect 4153 402 4174 458
rect 4076 381 4174 402
rect 5324 458 5422 479
rect 5324 402 5345 458
rect 5401 402 5422 458
rect 5324 381 5422 402
rect 6572 458 6670 479
rect 6572 402 6593 458
rect 6649 402 6670 458
rect 6572 381 6670 402
rect 7820 458 7918 479
rect 7820 402 7841 458
rect 7897 402 7918 458
rect 7820 381 7918 402
rect 9068 458 9166 479
rect 9068 402 9089 458
rect 9145 402 9166 458
rect 9068 381 9166 402
rect 10316 458 10414 479
rect 10316 402 10337 458
rect 10393 402 10414 458
rect 10316 381 10414 402
rect 11564 458 11662 479
rect 11564 402 11585 458
rect 11641 402 11662 458
rect 11564 381 11662 402
rect 12812 458 12910 479
rect 12812 402 12833 458
rect 12889 402 12910 458
rect 12812 381 12910 402
rect 14060 458 14158 479
rect 14060 402 14081 458
rect 14137 402 14158 458
rect 14060 381 14158 402
rect 15308 458 15406 479
rect 15308 402 15329 458
rect 15385 402 15406 458
rect 15308 381 15406 402
rect 16556 458 16654 479
rect 16556 402 16577 458
rect 16633 402 16654 458
rect 16556 381 16654 402
rect 17804 458 17902 479
rect 17804 402 17825 458
rect 17881 402 17902 458
rect 17804 381 17902 402
rect 19052 458 19150 479
rect 19052 402 19073 458
rect 19129 402 19150 458
rect 19052 381 19150 402
rect 20300 458 20398 479
rect 20300 402 20321 458
rect 20377 402 20398 458
rect 20300 381 20398 402
rect 21548 458 21646 479
rect 21548 402 21569 458
rect 21625 402 21646 458
rect 21548 381 21646 402
rect 22796 458 22894 479
rect 22796 402 22817 458
rect 22873 402 22894 458
rect 22796 381 22894 402
rect 24044 458 24142 479
rect 24044 402 24065 458
rect 24121 402 24142 458
rect 24044 381 24142 402
rect 25292 458 25390 479
rect 25292 402 25313 458
rect 25369 402 25390 458
rect 25292 381 25390 402
rect 26540 458 26638 479
rect 26540 402 26561 458
rect 26617 402 26638 458
rect 26540 381 26638 402
rect 27788 458 27886 479
rect 27788 402 27809 458
rect 27865 402 27886 458
rect 27788 381 27886 402
rect 29036 458 29134 479
rect 29036 402 29057 458
rect 29113 402 29134 458
rect 29036 381 29134 402
rect 30284 458 30382 479
rect 30284 402 30305 458
rect 30361 402 30382 458
rect 30284 381 30382 402
rect 31532 458 31630 479
rect 31532 402 31553 458
rect 31609 402 31630 458
rect 31532 381 31630 402
rect 32780 458 32878 479
rect 32780 402 32801 458
rect 32857 402 32878 458
rect 32780 381 32878 402
rect 34028 458 34126 479
rect 34028 402 34049 458
rect 34105 402 34126 458
rect 34028 381 34126 402
rect 35276 458 35374 479
rect 35276 402 35297 458
rect 35353 402 35374 458
rect 35276 381 35374 402
rect 36524 458 36622 479
rect 36524 402 36545 458
rect 36601 402 36622 458
rect 36524 381 36622 402
rect 37772 458 37870 479
rect 37772 402 37793 458
rect 37849 402 37870 458
rect 37772 381 37870 402
rect 39020 458 39118 479
rect 39020 402 39041 458
rect 39097 402 39118 458
rect 39020 381 39118 402
rect 332 136 430 157
rect 332 80 353 136
rect 409 80 430 136
rect 332 59 430 80
rect 1580 136 1678 157
rect 1580 80 1601 136
rect 1657 80 1678 136
rect 1580 59 1678 80
rect 2828 136 2926 157
rect 2828 80 2849 136
rect 2905 80 2926 136
rect 2828 59 2926 80
rect 4076 136 4174 157
rect 4076 80 4097 136
rect 4153 80 4174 136
rect 4076 59 4174 80
rect 5324 136 5422 157
rect 5324 80 5345 136
rect 5401 80 5422 136
rect 5324 59 5422 80
rect 6572 136 6670 157
rect 6572 80 6593 136
rect 6649 80 6670 136
rect 6572 59 6670 80
rect 7820 136 7918 157
rect 7820 80 7841 136
rect 7897 80 7918 136
rect 7820 59 7918 80
rect 9068 136 9166 157
rect 9068 80 9089 136
rect 9145 80 9166 136
rect 9068 59 9166 80
rect 10316 136 10414 157
rect 10316 80 10337 136
rect 10393 80 10414 136
rect 10316 59 10414 80
rect 11564 136 11662 157
rect 11564 80 11585 136
rect 11641 80 11662 136
rect 11564 59 11662 80
rect 12812 136 12910 157
rect 12812 80 12833 136
rect 12889 80 12910 136
rect 12812 59 12910 80
rect 14060 136 14158 157
rect 14060 80 14081 136
rect 14137 80 14158 136
rect 14060 59 14158 80
rect 15308 136 15406 157
rect 15308 80 15329 136
rect 15385 80 15406 136
rect 15308 59 15406 80
rect 16556 136 16654 157
rect 16556 80 16577 136
rect 16633 80 16654 136
rect 16556 59 16654 80
rect 17804 136 17902 157
rect 17804 80 17825 136
rect 17881 80 17902 136
rect 17804 59 17902 80
rect 19052 136 19150 157
rect 19052 80 19073 136
rect 19129 80 19150 136
rect 19052 59 19150 80
rect 20300 136 20398 157
rect 20300 80 20321 136
rect 20377 80 20398 136
rect 20300 59 20398 80
rect 21548 136 21646 157
rect 21548 80 21569 136
rect 21625 80 21646 136
rect 21548 59 21646 80
rect 22796 136 22894 157
rect 22796 80 22817 136
rect 22873 80 22894 136
rect 22796 59 22894 80
rect 24044 136 24142 157
rect 24044 80 24065 136
rect 24121 80 24142 136
rect 24044 59 24142 80
rect 25292 136 25390 157
rect 25292 80 25313 136
rect 25369 80 25390 136
rect 25292 59 25390 80
rect 26540 136 26638 157
rect 26540 80 26561 136
rect 26617 80 26638 136
rect 26540 59 26638 80
rect 27788 136 27886 157
rect 27788 80 27809 136
rect 27865 80 27886 136
rect 27788 59 27886 80
rect 29036 136 29134 157
rect 29036 80 29057 136
rect 29113 80 29134 136
rect 29036 59 29134 80
rect 30284 136 30382 157
rect 30284 80 30305 136
rect 30361 80 30382 136
rect 30284 59 30382 80
rect 31532 136 31630 157
rect 31532 80 31553 136
rect 31609 80 31630 136
rect 31532 59 31630 80
rect 32780 136 32878 157
rect 32780 80 32801 136
rect 32857 80 32878 136
rect 32780 59 32878 80
rect 34028 136 34126 157
rect 34028 80 34049 136
rect 34105 80 34126 136
rect 34028 59 34126 80
rect 35276 136 35374 157
rect 35276 80 35297 136
rect 35353 80 35374 136
rect 35276 59 35374 80
rect 36524 136 36622 157
rect 36524 80 36545 136
rect 36601 80 36622 136
rect 36524 59 36622 80
rect 37772 136 37870 157
rect 37772 80 37793 136
rect 37849 80 37870 136
rect 37772 59 37870 80
rect 39020 136 39118 157
rect 39020 80 39041 136
rect 39097 80 39118 136
rect 39020 59 39118 80
use contact_8  contact_8_0
timestamp 1676037725
transform 1 0 8827 0 1 2162
box 0 0 1 1
use contact_8  contact_8_1
timestamp 1676037725
transform 1 0 7579 0 1 2162
box 0 0 1 1
use contact_8  contact_8_2
timestamp 1676037725
transform 1 0 6331 0 1 2162
box 0 0 1 1
use contact_8  contact_8_3
timestamp 1676037725
transform 1 0 5083 0 1 2162
box 0 0 1 1
use contact_8  contact_8_4
timestamp 1676037725
transform 1 0 3835 0 1 2162
box 0 0 1 1
use contact_8  contact_8_5
timestamp 1676037725
transform 1 0 2587 0 1 2162
box 0 0 1 1
use contact_8  contact_8_6
timestamp 1676037725
transform 1 0 1339 0 1 2162
box 0 0 1 1
use contact_8  contact_8_7
timestamp 1676037725
transform 1 0 91 0 1 2162
box 0 0 1 1
use contact_8  contact_8_8
timestamp 1676037725
transform 1 0 18811 0 1 2162
box 0 0 1 1
use contact_8  contact_8_9
timestamp 1676037725
transform 1 0 17563 0 1 2162
box 0 0 1 1
use contact_8  contact_8_10
timestamp 1676037725
transform 1 0 16315 0 1 2162
box 0 0 1 1
use contact_8  contact_8_11
timestamp 1676037725
transform 1 0 15067 0 1 2162
box 0 0 1 1
use contact_8  contact_8_12
timestamp 1676037725
transform 1 0 13819 0 1 2162
box 0 0 1 1
use contact_8  contact_8_13
timestamp 1676037725
transform 1 0 12571 0 1 2162
box 0 0 1 1
use contact_8  contact_8_14
timestamp 1676037725
transform 1 0 11323 0 1 2162
box 0 0 1 1
use contact_8  contact_8_15
timestamp 1676037725
transform 1 0 10075 0 1 2162
box 0 0 1 1
use contact_8  contact_8_16
timestamp 1676037725
transform 1 0 23803 0 1 2162
box 0 0 1 1
use contact_8  contact_8_17
timestamp 1676037725
transform 1 0 22555 0 1 2162
box 0 0 1 1
use contact_8  contact_8_18
timestamp 1676037725
transform 1 0 21307 0 1 2162
box 0 0 1 1
use contact_8  contact_8_19
timestamp 1676037725
transform 1 0 20059 0 1 2162
box 0 0 1 1
use contact_8  contact_8_20
timestamp 1676037725
transform 1 0 28795 0 1 2162
box 0 0 1 1
use contact_8  contact_8_21
timestamp 1676037725
transform 1 0 27547 0 1 2162
box 0 0 1 1
use contact_8  contact_8_22
timestamp 1676037725
transform 1 0 26299 0 1 2162
box 0 0 1 1
use contact_8  contact_8_23
timestamp 1676037725
transform 1 0 25051 0 1 2162
box 0 0 1 1
use contact_8  contact_8_24
timestamp 1676037725
transform 1 0 38779 0 1 2162
box 0 0 1 1
use contact_8  contact_8_25
timestamp 1676037725
transform 1 0 37531 0 1 2162
box 0 0 1 1
use contact_8  contact_8_26
timestamp 1676037725
transform 1 0 36283 0 1 2162
box 0 0 1 1
use contact_8  contact_8_27
timestamp 1676037725
transform 1 0 35035 0 1 2162
box 0 0 1 1
use contact_8  contact_8_28
timestamp 1676037725
transform 1 0 33787 0 1 2162
box 0 0 1 1
use contact_8  contact_8_29
timestamp 1676037725
transform 1 0 32539 0 1 2162
box 0 0 1 1
use contact_8  contact_8_30
timestamp 1676037725
transform 1 0 31291 0 1 2162
box 0 0 1 1
use contact_8  contact_8_31
timestamp 1676037725
transform 1 0 30043 0 1 2162
box 0 0 1 1
use contact_9  contact_9_0
timestamp 1676037725
transform 1 0 8826 0 1 2157
box 0 0 1 1
use contact_9  contact_9_1
timestamp 1676037725
transform 1 0 7578 0 1 2157
box 0 0 1 1
use contact_9  contact_9_2
timestamp 1676037725
transform 1 0 6330 0 1 2157
box 0 0 1 1
use contact_9  contact_9_3
timestamp 1676037725
transform 1 0 5082 0 1 2157
box 0 0 1 1
use contact_9  contact_9_4
timestamp 1676037725
transform 1 0 3834 0 1 2157
box 0 0 1 1
use contact_9  contact_9_5
timestamp 1676037725
transform 1 0 2586 0 1 2157
box 0 0 1 1
use contact_9  contact_9_6
timestamp 1676037725
transform 1 0 1338 0 1 2157
box 0 0 1 1
use contact_9  contact_9_7
timestamp 1676037725
transform 1 0 90 0 1 2157
box 0 0 1 1
use contact_9  contact_9_8
timestamp 1676037725
transform 1 0 18810 0 1 2157
box 0 0 1 1
use contact_9  contact_9_9
timestamp 1676037725
transform 1 0 17562 0 1 2157
box 0 0 1 1
use contact_9  contact_9_10
timestamp 1676037725
transform 1 0 16314 0 1 2157
box 0 0 1 1
use contact_9  contact_9_11
timestamp 1676037725
transform 1 0 15066 0 1 2157
box 0 0 1 1
use contact_9  contact_9_12
timestamp 1676037725
transform 1 0 13818 0 1 2157
box 0 0 1 1
use contact_9  contact_9_13
timestamp 1676037725
transform 1 0 12570 0 1 2157
box 0 0 1 1
use contact_9  contact_9_14
timestamp 1676037725
transform 1 0 11322 0 1 2157
box 0 0 1 1
use contact_9  contact_9_15
timestamp 1676037725
transform 1 0 10074 0 1 2157
box 0 0 1 1
use contact_9  contact_9_16
timestamp 1676037725
transform 1 0 23802 0 1 2157
box 0 0 1 1
use contact_9  contact_9_17
timestamp 1676037725
transform 1 0 22554 0 1 2157
box 0 0 1 1
use contact_9  contact_9_18
timestamp 1676037725
transform 1 0 21306 0 1 2157
box 0 0 1 1
use contact_9  contact_9_19
timestamp 1676037725
transform 1 0 20058 0 1 2157
box 0 0 1 1
use contact_9  contact_9_20
timestamp 1676037725
transform 1 0 28794 0 1 2157
box 0 0 1 1
use contact_9  contact_9_21
timestamp 1676037725
transform 1 0 27546 0 1 2157
box 0 0 1 1
use contact_9  contact_9_22
timestamp 1676037725
transform 1 0 26298 0 1 2157
box 0 0 1 1
use contact_9  contact_9_23
timestamp 1676037725
transform 1 0 25050 0 1 2157
box 0 0 1 1
use contact_9  contact_9_24
timestamp 1676037725
transform 1 0 38778 0 1 2157
box 0 0 1 1
use contact_9  contact_9_25
timestamp 1676037725
transform 1 0 37530 0 1 2157
box 0 0 1 1
use contact_9  contact_9_26
timestamp 1676037725
transform 1 0 36282 0 1 2157
box 0 0 1 1
use contact_9  contact_9_27
timestamp 1676037725
transform 1 0 35034 0 1 2157
box 0 0 1 1
use contact_9  contact_9_28
timestamp 1676037725
transform 1 0 33786 0 1 2157
box 0 0 1 1
use contact_9  contact_9_29
timestamp 1676037725
transform 1 0 32538 0 1 2157
box 0 0 1 1
use contact_9  contact_9_30
timestamp 1676037725
transform 1 0 31290 0 1 2157
box 0 0 1 1
use contact_9  contact_9_31
timestamp 1676037725
transform 1 0 30042 0 1 2157
box 0 0 1 1
use contact_14  contact_14_0
timestamp 1676037725
transform 1 0 5335 0 1 1236
box 0 0 1 1
use contact_14  contact_14_1
timestamp 1676037725
transform 1 0 7843 0 1 76
box 0 0 1 1
use contact_14  contact_14_2
timestamp 1676037725
transform 1 0 5417 0 1 2010
box 0 0 1 1
use contact_14  contact_14_3
timestamp 1676037725
transform 1 0 355 0 1 398
box 0 0 1 1
use contact_14  contact_14_4
timestamp 1676037725
transform 1 0 4087 0 1 1236
box 0 0 1 1
use contact_14  contact_14_5
timestamp 1676037725
transform 1 0 6595 0 1 398
box 0 0 1 1
use contact_14  contact_14_6
timestamp 1676037725
transform 1 0 4169 0 1 2010
box 0 0 1 1
use contact_14  contact_14_7
timestamp 1676037725
transform 1 0 2851 0 1 398
box 0 0 1 1
use contact_14  contact_14_8
timestamp 1676037725
transform 1 0 2839 0 1 1236
box 0 0 1 1
use contact_14  contact_14_9
timestamp 1676037725
transform 1 0 6595 0 1 76
box 0 0 1 1
use contact_14  contact_14_10
timestamp 1676037725
transform 1 0 2921 0 1 2010
box 0 0 1 1
use contact_14  contact_14_11
timestamp 1676037725
transform 1 0 1603 0 1 76
box 0 0 1 1
use contact_14  contact_14_12
timestamp 1676037725
transform 1 0 1591 0 1 1236
box 0 0 1 1
use contact_14  contact_14_13
timestamp 1676037725
transform 1 0 5347 0 1 398
box 0 0 1 1
use contact_14  contact_14_14
timestamp 1676037725
transform 1 0 1673 0 1 2010
box 0 0 1 1
use contact_14  contact_14_15
timestamp 1676037725
transform 1 0 2851 0 1 76
box 0 0 1 1
use contact_14  contact_14_16
timestamp 1676037725
transform 1 0 343 0 1 1236
box 0 0 1 1
use contact_14  contact_14_17
timestamp 1676037725
transform 1 0 5347 0 1 76
box 0 0 1 1
use contact_14  contact_14_18
timestamp 1676037725
transform 1 0 425 0 1 2010
box 0 0 1 1
use contact_14  contact_14_19
timestamp 1676037725
transform 1 0 355 0 1 76
box 0 0 1 1
use contact_14  contact_14_20
timestamp 1676037725
transform 1 0 9079 0 1 1236
box 0 0 1 1
use contact_14  contact_14_21
timestamp 1676037725
transform 1 0 9091 0 1 398
box 0 0 1 1
use contact_14  contact_14_22
timestamp 1676037725
transform 1 0 9161 0 1 2010
box 0 0 1 1
use contact_14  contact_14_23
timestamp 1676037725
transform 1 0 4099 0 1 398
box 0 0 1 1
use contact_14  contact_14_24
timestamp 1676037725
transform 1 0 7831 0 1 1236
box 0 0 1 1
use contact_14  contact_14_25
timestamp 1676037725
transform 1 0 9091 0 1 76
box 0 0 1 1
use contact_14  contact_14_26
timestamp 1676037725
transform 1 0 7913 0 1 2010
box 0 0 1 1
use contact_14  contact_14_27
timestamp 1676037725
transform 1 0 1603 0 1 398
box 0 0 1 1
use contact_14  contact_14_28
timestamp 1676037725
transform 1 0 6583 0 1 1236
box 0 0 1 1
use contact_14  contact_14_29
timestamp 1676037725
transform 1 0 7843 0 1 398
box 0 0 1 1
use contact_14  contact_14_30
timestamp 1676037725
transform 1 0 6665 0 1 2010
box 0 0 1 1
use contact_14  contact_14_31
timestamp 1676037725
transform 1 0 4099 0 1 76
box 0 0 1 1
use contact_14  contact_14_32
timestamp 1676037725
transform 1 0 19063 0 1 1236
box 0 0 1 1
use contact_14  contact_14_33
timestamp 1676037725
transform 1 0 19145 0 1 2010
box 0 0 1 1
use contact_14  contact_14_34
timestamp 1676037725
transform 1 0 17815 0 1 1236
box 0 0 1 1
use contact_14  contact_14_35
timestamp 1676037725
transform 1 0 17897 0 1 2010
box 0 0 1 1
use contact_14  contact_14_36
timestamp 1676037725
transform 1 0 16567 0 1 1236
box 0 0 1 1
use contact_14  contact_14_37
timestamp 1676037725
transform 1 0 16649 0 1 2010
box 0 0 1 1
use contact_14  contact_14_38
timestamp 1676037725
transform 1 0 15319 0 1 1236
box 0 0 1 1
use contact_14  contact_14_39
timestamp 1676037725
transform 1 0 15401 0 1 2010
box 0 0 1 1
use contact_14  contact_14_40
timestamp 1676037725
transform 1 0 14071 0 1 1236
box 0 0 1 1
use contact_14  contact_14_41
timestamp 1676037725
transform 1 0 14153 0 1 2010
box 0 0 1 1
use contact_14  contact_14_42
timestamp 1676037725
transform 1 0 12823 0 1 1236
box 0 0 1 1
use contact_14  contact_14_43
timestamp 1676037725
transform 1 0 12905 0 1 2010
box 0 0 1 1
use contact_14  contact_14_44
timestamp 1676037725
transform 1 0 11575 0 1 1236
box 0 0 1 1
use contact_14  contact_14_45
timestamp 1676037725
transform 1 0 11657 0 1 2010
box 0 0 1 1
use contact_14  contact_14_46
timestamp 1676037725
transform 1 0 10327 0 1 1236
box 0 0 1 1
use contact_14  contact_14_47
timestamp 1676037725
transform 1 0 10409 0 1 2010
box 0 0 1 1
use contact_14  contact_14_48
timestamp 1676037725
transform 1 0 19075 0 1 398
box 0 0 1 1
use contact_14  contact_14_49
timestamp 1676037725
transform 1 0 19075 0 1 76
box 0 0 1 1
use contact_14  contact_14_50
timestamp 1676037725
transform 1 0 17827 0 1 398
box 0 0 1 1
use contact_14  contact_14_51
timestamp 1676037725
transform 1 0 17827 0 1 76
box 0 0 1 1
use contact_14  contact_14_52
timestamp 1676037725
transform 1 0 16579 0 1 398
box 0 0 1 1
use contact_14  contact_14_53
timestamp 1676037725
transform 1 0 16579 0 1 76
box 0 0 1 1
use contact_14  contact_14_54
timestamp 1676037725
transform 1 0 15331 0 1 398
box 0 0 1 1
use contact_14  contact_14_55
timestamp 1676037725
transform 1 0 15331 0 1 76
box 0 0 1 1
use contact_14  contact_14_56
timestamp 1676037725
transform 1 0 14083 0 1 398
box 0 0 1 1
use contact_14  contact_14_57
timestamp 1676037725
transform 1 0 14083 0 1 76
box 0 0 1 1
use contact_14  contact_14_58
timestamp 1676037725
transform 1 0 12835 0 1 398
box 0 0 1 1
use contact_14  contact_14_59
timestamp 1676037725
transform 1 0 12835 0 1 76
box 0 0 1 1
use contact_14  contact_14_60
timestamp 1676037725
transform 1 0 11587 0 1 398
box 0 0 1 1
use contact_14  contact_14_61
timestamp 1676037725
transform 1 0 11587 0 1 76
box 0 0 1 1
use contact_14  contact_14_62
timestamp 1676037725
transform 1 0 10339 0 1 398
box 0 0 1 1
use contact_14  contact_14_63
timestamp 1676037725
transform 1 0 10339 0 1 76
box 0 0 1 1
use contact_14  contact_14_64
timestamp 1676037725
transform 1 0 29059 0 1 398
box 0 0 1 1
use contact_14  contact_14_65
timestamp 1676037725
transform 1 0 24067 0 1 398
box 0 0 1 1
use contact_14  contact_14_66
timestamp 1676037725
transform 1 0 29059 0 1 76
box 0 0 1 1
use contact_14  contact_14_67
timestamp 1676037725
transform 1 0 21571 0 1 398
box 0 0 1 1
use contact_14  contact_14_68
timestamp 1676037725
transform 1 0 26551 0 1 1236
box 0 0 1 1
use contact_14  contact_14_69
timestamp 1676037725
transform 1 0 27811 0 1 398
box 0 0 1 1
use contact_14  contact_14_70
timestamp 1676037725
transform 1 0 26633 0 1 2010
box 0 0 1 1
use contact_14  contact_14_71
timestamp 1676037725
transform 1 0 24067 0 1 76
box 0 0 1 1
use contact_14  contact_14_72
timestamp 1676037725
transform 1 0 25303 0 1 1236
box 0 0 1 1
use contact_14  contact_14_73
timestamp 1676037725
transform 1 0 27811 0 1 76
box 0 0 1 1
use contact_14  contact_14_74
timestamp 1676037725
transform 1 0 25385 0 1 2010
box 0 0 1 1
use contact_14  contact_14_75
timestamp 1676037725
transform 1 0 20323 0 1 398
box 0 0 1 1
use contact_14  contact_14_76
timestamp 1676037725
transform 1 0 24055 0 1 1236
box 0 0 1 1
use contact_14  contact_14_77
timestamp 1676037725
transform 1 0 26563 0 1 398
box 0 0 1 1
use contact_14  contact_14_78
timestamp 1676037725
transform 1 0 24137 0 1 2010
box 0 0 1 1
use contact_14  contact_14_79
timestamp 1676037725
transform 1 0 22819 0 1 398
box 0 0 1 1
use contact_14  contact_14_80
timestamp 1676037725
transform 1 0 22807 0 1 1236
box 0 0 1 1
use contact_14  contact_14_81
timestamp 1676037725
transform 1 0 26563 0 1 76
box 0 0 1 1
use contact_14  contact_14_82
timestamp 1676037725
transform 1 0 22889 0 1 2010
box 0 0 1 1
use contact_14  contact_14_83
timestamp 1676037725
transform 1 0 21571 0 1 76
box 0 0 1 1
use contact_14  contact_14_84
timestamp 1676037725
transform 1 0 21559 0 1 1236
box 0 0 1 1
use contact_14  contact_14_85
timestamp 1676037725
transform 1 0 25315 0 1 398
box 0 0 1 1
use contact_14  contact_14_86
timestamp 1676037725
transform 1 0 21641 0 1 2010
box 0 0 1 1
use contact_14  contact_14_87
timestamp 1676037725
transform 1 0 22819 0 1 76
box 0 0 1 1
use contact_14  contact_14_88
timestamp 1676037725
transform 1 0 20311 0 1 1236
box 0 0 1 1
use contact_14  contact_14_89
timestamp 1676037725
transform 1 0 25315 0 1 76
box 0 0 1 1
use contact_14  contact_14_90
timestamp 1676037725
transform 1 0 20393 0 1 2010
box 0 0 1 1
use contact_14  contact_14_91
timestamp 1676037725
transform 1 0 20323 0 1 76
box 0 0 1 1
use contact_14  contact_14_92
timestamp 1676037725
transform 1 0 29047 0 1 1236
box 0 0 1 1
use contact_14  contact_14_93
timestamp 1676037725
transform 1 0 29129 0 1 2010
box 0 0 1 1
use contact_14  contact_14_94
timestamp 1676037725
transform 1 0 27799 0 1 1236
box 0 0 1 1
use contact_14  contact_14_95
timestamp 1676037725
transform 1 0 27881 0 1 2010
box 0 0 1 1
use contact_14  contact_14_96
timestamp 1676037725
transform 1 0 39043 0 1 398
box 0 0 1 1
use contact_14  contact_14_97
timestamp 1676037725
transform 1 0 39043 0 1 76
box 0 0 1 1
use contact_14  contact_14_98
timestamp 1676037725
transform 1 0 37795 0 1 398
box 0 0 1 1
use contact_14  contact_14_99
timestamp 1676037725
transform 1 0 37795 0 1 76
box 0 0 1 1
use contact_14  contact_14_100
timestamp 1676037725
transform 1 0 36547 0 1 398
box 0 0 1 1
use contact_14  contact_14_101
timestamp 1676037725
transform 1 0 36547 0 1 76
box 0 0 1 1
use contact_14  contact_14_102
timestamp 1676037725
transform 1 0 35299 0 1 398
box 0 0 1 1
use contact_14  contact_14_103
timestamp 1676037725
transform 1 0 35299 0 1 76
box 0 0 1 1
use contact_14  contact_14_104
timestamp 1676037725
transform 1 0 34051 0 1 398
box 0 0 1 1
use contact_14  contact_14_105
timestamp 1676037725
transform 1 0 34051 0 1 76
box 0 0 1 1
use contact_14  contact_14_106
timestamp 1676037725
transform 1 0 32803 0 1 398
box 0 0 1 1
use contact_14  contact_14_107
timestamp 1676037725
transform 1 0 32803 0 1 76
box 0 0 1 1
use contact_14  contact_14_108
timestamp 1676037725
transform 1 0 31555 0 1 398
box 0 0 1 1
use contact_14  contact_14_109
timestamp 1676037725
transform 1 0 31555 0 1 76
box 0 0 1 1
use contact_14  contact_14_110
timestamp 1676037725
transform 1 0 30307 0 1 398
box 0 0 1 1
use contact_14  contact_14_111
timestamp 1676037725
transform 1 0 30307 0 1 76
box 0 0 1 1
use contact_14  contact_14_112
timestamp 1676037725
transform 1 0 39031 0 1 1236
box 0 0 1 1
use contact_14  contact_14_113
timestamp 1676037725
transform 1 0 39113 0 1 2010
box 0 0 1 1
use contact_14  contact_14_114
timestamp 1676037725
transform 1 0 37783 0 1 1236
box 0 0 1 1
use contact_14  contact_14_115
timestamp 1676037725
transform 1 0 37865 0 1 2010
box 0 0 1 1
use contact_14  contact_14_116
timestamp 1676037725
transform 1 0 36535 0 1 1236
box 0 0 1 1
use contact_14  contact_14_117
timestamp 1676037725
transform 1 0 36617 0 1 2010
box 0 0 1 1
use contact_14  contact_14_118
timestamp 1676037725
transform 1 0 35287 0 1 1236
box 0 0 1 1
use contact_14  contact_14_119
timestamp 1676037725
transform 1 0 35369 0 1 2010
box 0 0 1 1
use contact_14  contact_14_120
timestamp 1676037725
transform 1 0 34039 0 1 1236
box 0 0 1 1
use contact_14  contact_14_121
timestamp 1676037725
transform 1 0 34121 0 1 2010
box 0 0 1 1
use contact_14  contact_14_122
timestamp 1676037725
transform 1 0 32791 0 1 1236
box 0 0 1 1
use contact_14  contact_14_123
timestamp 1676037725
transform 1 0 32873 0 1 2010
box 0 0 1 1
use contact_14  contact_14_124
timestamp 1676037725
transform 1 0 31543 0 1 1236
box 0 0 1 1
use contact_14  contact_14_125
timestamp 1676037725
transform 1 0 31625 0 1 2010
box 0 0 1 1
use contact_14  contact_14_126
timestamp 1676037725
transform 1 0 30295 0 1 1236
box 0 0 1 1
use contact_14  contact_14_127
timestamp 1676037725
transform 1 0 30377 0 1 2010
box 0 0 1 1
use contact_15  contact_15_0
timestamp 1676037725
transform 1 0 5328 0 1 1231
box 0 0 1 1
use contact_15  contact_15_1
timestamp 1676037725
transform 1 0 7836 0 1 71
box 0 0 1 1
use contact_15  contact_15_2
timestamp 1676037725
transform 1 0 5410 0 1 2005
box 0 0 1 1
use contact_15  contact_15_3
timestamp 1676037725
transform 1 0 348 0 1 393
box 0 0 1 1
use contact_15  contact_15_4
timestamp 1676037725
transform 1 0 4080 0 1 1231
box 0 0 1 1
use contact_15  contact_15_5
timestamp 1676037725
transform 1 0 6588 0 1 393
box 0 0 1 1
use contact_15  contact_15_6
timestamp 1676037725
transform 1 0 4162 0 1 2005
box 0 0 1 1
use contact_15  contact_15_7
timestamp 1676037725
transform 1 0 2844 0 1 393
box 0 0 1 1
use contact_15  contact_15_8
timestamp 1676037725
transform 1 0 2832 0 1 1231
box 0 0 1 1
use contact_15  contact_15_9
timestamp 1676037725
transform 1 0 6588 0 1 71
box 0 0 1 1
use contact_15  contact_15_10
timestamp 1676037725
transform 1 0 2914 0 1 2005
box 0 0 1 1
use contact_15  contact_15_11
timestamp 1676037725
transform 1 0 1596 0 1 71
box 0 0 1 1
use contact_15  contact_15_12
timestamp 1676037725
transform 1 0 1584 0 1 1231
box 0 0 1 1
use contact_15  contact_15_13
timestamp 1676037725
transform 1 0 5340 0 1 393
box 0 0 1 1
use contact_15  contact_15_14
timestamp 1676037725
transform 1 0 1666 0 1 2005
box 0 0 1 1
use contact_15  contact_15_15
timestamp 1676037725
transform 1 0 2844 0 1 71
box 0 0 1 1
use contact_15  contact_15_16
timestamp 1676037725
transform 1 0 336 0 1 1231
box 0 0 1 1
use contact_15  contact_15_17
timestamp 1676037725
transform 1 0 5340 0 1 71
box 0 0 1 1
use contact_15  contact_15_18
timestamp 1676037725
transform 1 0 418 0 1 2005
box 0 0 1 1
use contact_15  contact_15_19
timestamp 1676037725
transform 1 0 348 0 1 71
box 0 0 1 1
use contact_15  contact_15_20
timestamp 1676037725
transform 1 0 9072 0 1 1231
box 0 0 1 1
use contact_15  contact_15_21
timestamp 1676037725
transform 1 0 9084 0 1 393
box 0 0 1 1
use contact_15  contact_15_22
timestamp 1676037725
transform 1 0 9154 0 1 2005
box 0 0 1 1
use contact_15  contact_15_23
timestamp 1676037725
transform 1 0 4092 0 1 393
box 0 0 1 1
use contact_15  contact_15_24
timestamp 1676037725
transform 1 0 7824 0 1 1231
box 0 0 1 1
use contact_15  contact_15_25
timestamp 1676037725
transform 1 0 9084 0 1 71
box 0 0 1 1
use contact_15  contact_15_26
timestamp 1676037725
transform 1 0 7906 0 1 2005
box 0 0 1 1
use contact_15  contact_15_27
timestamp 1676037725
transform 1 0 1596 0 1 393
box 0 0 1 1
use contact_15  contact_15_28
timestamp 1676037725
transform 1 0 6576 0 1 1231
box 0 0 1 1
use contact_15  contact_15_29
timestamp 1676037725
transform 1 0 7836 0 1 393
box 0 0 1 1
use contact_15  contact_15_30
timestamp 1676037725
transform 1 0 6658 0 1 2005
box 0 0 1 1
use contact_15  contact_15_31
timestamp 1676037725
transform 1 0 4092 0 1 71
box 0 0 1 1
use contact_15  contact_15_32
timestamp 1676037725
transform 1 0 19056 0 1 1231
box 0 0 1 1
use contact_15  contact_15_33
timestamp 1676037725
transform 1 0 19138 0 1 2005
box 0 0 1 1
use contact_15  contact_15_34
timestamp 1676037725
transform 1 0 17808 0 1 1231
box 0 0 1 1
use contact_15  contact_15_35
timestamp 1676037725
transform 1 0 17890 0 1 2005
box 0 0 1 1
use contact_15  contact_15_36
timestamp 1676037725
transform 1 0 16560 0 1 1231
box 0 0 1 1
use contact_15  contact_15_37
timestamp 1676037725
transform 1 0 16642 0 1 2005
box 0 0 1 1
use contact_15  contact_15_38
timestamp 1676037725
transform 1 0 15312 0 1 1231
box 0 0 1 1
use contact_15  contact_15_39
timestamp 1676037725
transform 1 0 15394 0 1 2005
box 0 0 1 1
use contact_15  contact_15_40
timestamp 1676037725
transform 1 0 14064 0 1 1231
box 0 0 1 1
use contact_15  contact_15_41
timestamp 1676037725
transform 1 0 14146 0 1 2005
box 0 0 1 1
use contact_15  contact_15_42
timestamp 1676037725
transform 1 0 12816 0 1 1231
box 0 0 1 1
use contact_15  contact_15_43
timestamp 1676037725
transform 1 0 12898 0 1 2005
box 0 0 1 1
use contact_15  contact_15_44
timestamp 1676037725
transform 1 0 11568 0 1 1231
box 0 0 1 1
use contact_15  contact_15_45
timestamp 1676037725
transform 1 0 11650 0 1 2005
box 0 0 1 1
use contact_15  contact_15_46
timestamp 1676037725
transform 1 0 10320 0 1 1231
box 0 0 1 1
use contact_15  contact_15_47
timestamp 1676037725
transform 1 0 10402 0 1 2005
box 0 0 1 1
use contact_15  contact_15_48
timestamp 1676037725
transform 1 0 19068 0 1 393
box 0 0 1 1
use contact_15  contact_15_49
timestamp 1676037725
transform 1 0 19068 0 1 71
box 0 0 1 1
use contact_15  contact_15_50
timestamp 1676037725
transform 1 0 17820 0 1 393
box 0 0 1 1
use contact_15  contact_15_51
timestamp 1676037725
transform 1 0 17820 0 1 71
box 0 0 1 1
use contact_15  contact_15_52
timestamp 1676037725
transform 1 0 16572 0 1 393
box 0 0 1 1
use contact_15  contact_15_53
timestamp 1676037725
transform 1 0 16572 0 1 71
box 0 0 1 1
use contact_15  contact_15_54
timestamp 1676037725
transform 1 0 15324 0 1 393
box 0 0 1 1
use contact_15  contact_15_55
timestamp 1676037725
transform 1 0 15324 0 1 71
box 0 0 1 1
use contact_15  contact_15_56
timestamp 1676037725
transform 1 0 14076 0 1 393
box 0 0 1 1
use contact_15  contact_15_57
timestamp 1676037725
transform 1 0 14076 0 1 71
box 0 0 1 1
use contact_15  contact_15_58
timestamp 1676037725
transform 1 0 12828 0 1 393
box 0 0 1 1
use contact_15  contact_15_59
timestamp 1676037725
transform 1 0 12828 0 1 71
box 0 0 1 1
use contact_15  contact_15_60
timestamp 1676037725
transform 1 0 11580 0 1 393
box 0 0 1 1
use contact_15  contact_15_61
timestamp 1676037725
transform 1 0 11580 0 1 71
box 0 0 1 1
use contact_15  contact_15_62
timestamp 1676037725
transform 1 0 10332 0 1 393
box 0 0 1 1
use contact_15  contact_15_63
timestamp 1676037725
transform 1 0 10332 0 1 71
box 0 0 1 1
use contact_15  contact_15_64
timestamp 1676037725
transform 1 0 29052 0 1 393
box 0 0 1 1
use contact_15  contact_15_65
timestamp 1676037725
transform 1 0 24060 0 1 393
box 0 0 1 1
use contact_15  contact_15_66
timestamp 1676037725
transform 1 0 29052 0 1 71
box 0 0 1 1
use contact_15  contact_15_67
timestamp 1676037725
transform 1 0 21564 0 1 393
box 0 0 1 1
use contact_15  contact_15_68
timestamp 1676037725
transform 1 0 26544 0 1 1231
box 0 0 1 1
use contact_15  contact_15_69
timestamp 1676037725
transform 1 0 27804 0 1 393
box 0 0 1 1
use contact_15  contact_15_70
timestamp 1676037725
transform 1 0 26626 0 1 2005
box 0 0 1 1
use contact_15  contact_15_71
timestamp 1676037725
transform 1 0 24060 0 1 71
box 0 0 1 1
use contact_15  contact_15_72
timestamp 1676037725
transform 1 0 25296 0 1 1231
box 0 0 1 1
use contact_15  contact_15_73
timestamp 1676037725
transform 1 0 27804 0 1 71
box 0 0 1 1
use contact_15  contact_15_74
timestamp 1676037725
transform 1 0 25378 0 1 2005
box 0 0 1 1
use contact_15  contact_15_75
timestamp 1676037725
transform 1 0 20316 0 1 393
box 0 0 1 1
use contact_15  contact_15_76
timestamp 1676037725
transform 1 0 24048 0 1 1231
box 0 0 1 1
use contact_15  contact_15_77
timestamp 1676037725
transform 1 0 26556 0 1 393
box 0 0 1 1
use contact_15  contact_15_78
timestamp 1676037725
transform 1 0 24130 0 1 2005
box 0 0 1 1
use contact_15  contact_15_79
timestamp 1676037725
transform 1 0 22812 0 1 393
box 0 0 1 1
use contact_15  contact_15_80
timestamp 1676037725
transform 1 0 22800 0 1 1231
box 0 0 1 1
use contact_15  contact_15_81
timestamp 1676037725
transform 1 0 26556 0 1 71
box 0 0 1 1
use contact_15  contact_15_82
timestamp 1676037725
transform 1 0 22882 0 1 2005
box 0 0 1 1
use contact_15  contact_15_83
timestamp 1676037725
transform 1 0 21564 0 1 71
box 0 0 1 1
use contact_15  contact_15_84
timestamp 1676037725
transform 1 0 21552 0 1 1231
box 0 0 1 1
use contact_15  contact_15_85
timestamp 1676037725
transform 1 0 25308 0 1 393
box 0 0 1 1
use contact_15  contact_15_86
timestamp 1676037725
transform 1 0 21634 0 1 2005
box 0 0 1 1
use contact_15  contact_15_87
timestamp 1676037725
transform 1 0 22812 0 1 71
box 0 0 1 1
use contact_15  contact_15_88
timestamp 1676037725
transform 1 0 20304 0 1 1231
box 0 0 1 1
use contact_15  contact_15_89
timestamp 1676037725
transform 1 0 25308 0 1 71
box 0 0 1 1
use contact_15  contact_15_90
timestamp 1676037725
transform 1 0 20386 0 1 2005
box 0 0 1 1
use contact_15  contact_15_91
timestamp 1676037725
transform 1 0 20316 0 1 71
box 0 0 1 1
use contact_15  contact_15_92
timestamp 1676037725
transform 1 0 29040 0 1 1231
box 0 0 1 1
use contact_15  contact_15_93
timestamp 1676037725
transform 1 0 29122 0 1 2005
box 0 0 1 1
use contact_15  contact_15_94
timestamp 1676037725
transform 1 0 27792 0 1 1231
box 0 0 1 1
use contact_15  contact_15_95
timestamp 1676037725
transform 1 0 27874 0 1 2005
box 0 0 1 1
use contact_15  contact_15_96
timestamp 1676037725
transform 1 0 39036 0 1 393
box 0 0 1 1
use contact_15  contact_15_97
timestamp 1676037725
transform 1 0 39036 0 1 71
box 0 0 1 1
use contact_15  contact_15_98
timestamp 1676037725
transform 1 0 37788 0 1 393
box 0 0 1 1
use contact_15  contact_15_99
timestamp 1676037725
transform 1 0 37788 0 1 71
box 0 0 1 1
use contact_15  contact_15_100
timestamp 1676037725
transform 1 0 36540 0 1 393
box 0 0 1 1
use contact_15  contact_15_101
timestamp 1676037725
transform 1 0 36540 0 1 71
box 0 0 1 1
use contact_15  contact_15_102
timestamp 1676037725
transform 1 0 35292 0 1 393
box 0 0 1 1
use contact_15  contact_15_103
timestamp 1676037725
transform 1 0 35292 0 1 71
box 0 0 1 1
use contact_15  contact_15_104
timestamp 1676037725
transform 1 0 34044 0 1 393
box 0 0 1 1
use contact_15  contact_15_105
timestamp 1676037725
transform 1 0 34044 0 1 71
box 0 0 1 1
use contact_15  contact_15_106
timestamp 1676037725
transform 1 0 32796 0 1 393
box 0 0 1 1
use contact_15  contact_15_107
timestamp 1676037725
transform 1 0 32796 0 1 71
box 0 0 1 1
use contact_15  contact_15_108
timestamp 1676037725
transform 1 0 31548 0 1 393
box 0 0 1 1
use contact_15  contact_15_109
timestamp 1676037725
transform 1 0 31548 0 1 71
box 0 0 1 1
use contact_15  contact_15_110
timestamp 1676037725
transform 1 0 30300 0 1 393
box 0 0 1 1
use contact_15  contact_15_111
timestamp 1676037725
transform 1 0 30300 0 1 71
box 0 0 1 1
use contact_15  contact_15_112
timestamp 1676037725
transform 1 0 39024 0 1 1231
box 0 0 1 1
use contact_15  contact_15_113
timestamp 1676037725
transform 1 0 39106 0 1 2005
box 0 0 1 1
use contact_15  contact_15_114
timestamp 1676037725
transform 1 0 37776 0 1 1231
box 0 0 1 1
use contact_15  contact_15_115
timestamp 1676037725
transform 1 0 37858 0 1 2005
box 0 0 1 1
use contact_15  contact_15_116
timestamp 1676037725
transform 1 0 36528 0 1 1231
box 0 0 1 1
use contact_15  contact_15_117
timestamp 1676037725
transform 1 0 36610 0 1 2005
box 0 0 1 1
use contact_15  contact_15_118
timestamp 1676037725
transform 1 0 35280 0 1 1231
box 0 0 1 1
use contact_15  contact_15_119
timestamp 1676037725
transform 1 0 35362 0 1 2005
box 0 0 1 1
use contact_15  contact_15_120
timestamp 1676037725
transform 1 0 34032 0 1 1231
box 0 0 1 1
use contact_15  contact_15_121
timestamp 1676037725
transform 1 0 34114 0 1 2005
box 0 0 1 1
use contact_15  contact_15_122
timestamp 1676037725
transform 1 0 32784 0 1 1231
box 0 0 1 1
use contact_15  contact_15_123
timestamp 1676037725
transform 1 0 32866 0 1 2005
box 0 0 1 1
use contact_15  contact_15_124
timestamp 1676037725
transform 1 0 31536 0 1 1231
box 0 0 1 1
use contact_15  contact_15_125
timestamp 1676037725
transform 1 0 31618 0 1 2005
box 0 0 1 1
use contact_15  contact_15_126
timestamp 1676037725
transform 1 0 30288 0 1 1231
box 0 0 1 1
use contact_15  contact_15_127
timestamp 1676037725
transform 1 0 30370 0 1 2005
box 0 0 1 1
use sense_amp  sense_amp_0
timestamp 1676037725
transform 1 0 8736 0 1 0
box -160 0 684 2256
use sense_amp  sense_amp_1
timestamp 1676037725
transform 1 0 7488 0 1 0
box -160 0 684 2256
use sense_amp  sense_amp_2
timestamp 1676037725
transform 1 0 6240 0 1 0
box -160 0 684 2256
use sense_amp  sense_amp_3
timestamp 1676037725
transform 1 0 4992 0 1 0
box -160 0 684 2256
use sense_amp  sense_amp_4
timestamp 1676037725
transform 1 0 3744 0 1 0
box -160 0 684 2256
use sense_amp  sense_amp_5
timestamp 1676037725
transform 1 0 2496 0 1 0
box -160 0 684 2256
use sense_amp  sense_amp_6
timestamp 1676037725
transform 1 0 1248 0 1 0
box -160 0 684 2256
use sense_amp  sense_amp_7
timestamp 1676037725
transform 1 0 0 0 1 0
box -160 0 684 2256
use sense_amp  sense_amp_8
timestamp 1676037725
transform 1 0 18720 0 1 0
box -160 0 684 2256
use sense_amp  sense_amp_9
timestamp 1676037725
transform 1 0 17472 0 1 0
box -160 0 684 2256
use sense_amp  sense_amp_10
timestamp 1676037725
transform 1 0 16224 0 1 0
box -160 0 684 2256
use sense_amp  sense_amp_11
timestamp 1676037725
transform 1 0 14976 0 1 0
box -160 0 684 2256
use sense_amp  sense_amp_12
timestamp 1676037725
transform 1 0 13728 0 1 0
box -160 0 684 2256
use sense_amp  sense_amp_13
timestamp 1676037725
transform 1 0 12480 0 1 0
box -160 0 684 2256
use sense_amp  sense_amp_14
timestamp 1676037725
transform 1 0 11232 0 1 0
box -160 0 684 2256
use sense_amp  sense_amp_15
timestamp 1676037725
transform 1 0 9984 0 1 0
box -160 0 684 2256
use sense_amp  sense_amp_16
timestamp 1676037725
transform 1 0 28704 0 1 0
box -160 0 684 2256
use sense_amp  sense_amp_17
timestamp 1676037725
transform 1 0 27456 0 1 0
box -160 0 684 2256
use sense_amp  sense_amp_18
timestamp 1676037725
transform 1 0 26208 0 1 0
box -160 0 684 2256
use sense_amp  sense_amp_19
timestamp 1676037725
transform 1 0 24960 0 1 0
box -160 0 684 2256
use sense_amp  sense_amp_20
timestamp 1676037725
transform 1 0 23712 0 1 0
box -160 0 684 2256
use sense_amp  sense_amp_21
timestamp 1676037725
transform 1 0 22464 0 1 0
box -160 0 684 2256
use sense_amp  sense_amp_22
timestamp 1676037725
transform 1 0 21216 0 1 0
box -160 0 684 2256
use sense_amp  sense_amp_23
timestamp 1676037725
transform 1 0 19968 0 1 0
box -160 0 684 2256
use sense_amp  sense_amp_24
timestamp 1676037725
transform 1 0 38688 0 1 0
box -160 0 684 2256
use sense_amp  sense_amp_25
timestamp 1676037725
transform 1 0 37440 0 1 0
box -160 0 684 2256
use sense_amp  sense_amp_26
timestamp 1676037725
transform 1 0 36192 0 1 0
box -160 0 684 2256
use sense_amp  sense_amp_27
timestamp 1676037725
transform 1 0 34944 0 1 0
box -160 0 684 2256
use sense_amp  sense_amp_28
timestamp 1676037725
transform 1 0 33696 0 1 0
box -160 0 684 2256
use sense_amp  sense_amp_29
timestamp 1676037725
transform 1 0 32448 0 1 0
box -160 0 684 2256
use sense_amp  sense_amp_30
timestamp 1676037725
transform 1 0 31200 0 1 0
box -160 0 684 2256
use sense_amp  sense_amp_31
timestamp 1676037725
transform 1 0 29952 0 1 0
box -160 0 684 2256
<< labels >>
rlabel metal1 s 28917 1693 28917 1693 4 bl_23
port 71 nsew
rlabel metal1 s 14014 1699 14014 1699 4 br_11
port 36 nsew
rlabel metal1 s 1534 1699 1534 1699 4 br_1
port 6 nsew
rlabel metal1 s 2709 1693 2709 1693 4 bl_2
port 8 nsew
rlabel metal1 s 15262 1699 15262 1699 4 br_12
port 39 nsew
rlabel metal1 s 21343 127 21343 127 4 data_17
port 52 nsew
rlabel metal1 s 213 1693 213 1693 4 bl_0
port 2 nsew
rlabel metal1 s 28990 1699 28990 1699 4 br_23
port 72 nsew
rlabel metal1 s 17599 127 17599 127 4 data_14
port 43 nsew
rlabel metal1 s 18847 127 18847 127 4 data_15
port 46 nsew
rlabel metal1 s 35230 1699 35230 1699 4 br_28
port 87 nsew
rlabel metal1 s 32661 1693 32661 1693 4 bl_26
port 80 nsew
rlabel metal1 s 22591 127 22591 127 4 data_18
port 55 nsew
rlabel metal1 s 5278 1699 5278 1699 4 br_4
port 15 nsew
rlabel metal1 s 36319 127 36319 127 4 data_29
port 88 nsew
rlabel metal1 s 17685 1693 17685 1693 4 bl_14
port 44 nsew
rlabel metal1 s 12693 1693 12693 1693 4 bl_10
port 32 nsew
rlabel metal1 s 20181 1693 20181 1693 4 bl_16
port 50 nsew
rlabel metal1 s 31327 127 31327 127 4 data_25
port 76 nsew
rlabel metal1 s 38901 1693 38901 1693 4 bl_31
port 95 nsew
rlabel metal1 s 37653 1693 37653 1693 4 bl_30
port 92 nsew
rlabel metal1 s 6367 127 6367 127 4 data_5
port 16 nsew
rlabel metal1 s 32575 127 32575 127 4 data_26
port 79 nsew
rlabel metal1 s 3957 1693 3957 1693 4 bl_3
port 11 nsew
rlabel metal1 s 286 1699 286 1699 4 br_0
port 3 nsew
rlabel metal1 s 22677 1693 22677 1693 4 bl_18
port 56 nsew
rlabel metal1 s 15189 1693 15189 1693 4 bl_12
port 38 nsew
rlabel metal1 s 16510 1699 16510 1699 4 br_13
port 42 nsew
rlabel metal1 s 35071 127 35071 127 4 data_28
port 85 nsew
rlabel metal1 s 27742 1699 27742 1699 4 br_22
port 69 nsew
rlabel metal1 s 33909 1693 33909 1693 4 bl_27
port 83 nsew
rlabel metal1 s 1375 127 1375 127 4 data_1
port 4 nsew
rlabel metal1 s 20254 1699 20254 1699 4 br_16
port 51 nsew
rlabel metal1 s 4030 1699 4030 1699 4 br_3
port 12 nsew
rlabel metal1 s 23925 1693 23925 1693 4 bl_19
port 59 nsew
rlabel metal1 s 8863 127 8863 127 4 data_7
port 22 nsew
rlabel metal1 s 27583 127 27583 127 4 data_22
port 67 nsew
rlabel metal1 s 27669 1693 27669 1693 4 bl_22
port 68 nsew
rlabel metal1 s 21429 1693 21429 1693 4 bl_17
port 53 nsew
rlabel metal1 s 7701 1693 7701 1693 4 bl_6
port 20 nsew
rlabel metal1 s 38974 1699 38974 1699 4 br_31
port 96 nsew
rlabel metal1 s 26421 1693 26421 1693 4 bl_21
port 65 nsew
rlabel metal1 s 127 127 127 127 4 data_0
port 1 nsew
rlabel metal1 s 16351 127 16351 127 4 data_13
port 40 nsew
rlabel metal1 s 12766 1699 12766 1699 4 br_10
port 33 nsew
rlabel metal1 s 15103 127 15103 127 4 data_12
port 37 nsew
rlabel metal1 s 32734 1699 32734 1699 4 br_26
port 81 nsew
rlabel metal1 s 22750 1699 22750 1699 4 br_18
port 57 nsew
rlabel metal1 s 1461 1693 1461 1693 4 bl_1
port 5 nsew
rlabel metal1 s 36478 1699 36478 1699 4 br_29
port 90 nsew
rlabel metal1 s 28831 127 28831 127 4 data_23
port 70 nsew
rlabel metal1 s 36405 1693 36405 1693 4 bl_29
port 89 nsew
rlabel metal1 s 30165 1693 30165 1693 4 bl_24
port 74 nsew
rlabel metal1 s 12607 127 12607 127 4 data_10
port 31 nsew
rlabel metal1 s 37726 1699 37726 1699 4 br_30
port 93 nsew
rlabel metal1 s 6453 1693 6453 1693 4 bl_5
port 17 nsew
rlabel metal1 s 21502 1699 21502 1699 4 br_17
port 54 nsew
rlabel metal1 s 25173 1693 25173 1693 4 bl_20
port 62 nsew
rlabel metal1 s 8949 1693 8949 1693 4 bl_7
port 23 nsew
rlabel metal1 s 11518 1699 11518 1699 4 br_9
port 30 nsew
rlabel metal1 s 26494 1699 26494 1699 4 br_21
port 66 nsew
rlabel metal1 s 7615 127 7615 127 4 data_6
port 19 nsew
rlabel metal1 s 20095 127 20095 127 4 data_16
port 49 nsew
rlabel metal1 s 11359 127 11359 127 4 data_9
port 28 nsew
rlabel metal1 s 7774 1699 7774 1699 4 br_6
port 21 nsew
rlabel metal1 s 31413 1693 31413 1693 4 bl_25
port 77 nsew
rlabel metal1 s 13941 1693 13941 1693 4 bl_11
port 35 nsew
rlabel metal1 s 25246 1699 25246 1699 4 br_20
port 63 nsew
rlabel metal1 s 5119 127 5119 127 4 data_4
port 13 nsew
rlabel metal1 s 31486 1699 31486 1699 4 br_25
port 78 nsew
rlabel metal1 s 2623 127 2623 127 4 data_2
port 7 nsew
rlabel metal1 s 25087 127 25087 127 4 data_20
port 61 nsew
rlabel metal1 s 38815 127 38815 127 4 data_31
port 94 nsew
rlabel metal1 s 19006 1699 19006 1699 4 br_15
port 48 nsew
rlabel metal1 s 6526 1699 6526 1699 4 br_5
port 18 nsew
rlabel metal1 s 23998 1699 23998 1699 4 br_19
port 60 nsew
rlabel metal1 s 18933 1693 18933 1693 4 bl_15
port 47 nsew
rlabel metal1 s 16437 1693 16437 1693 4 bl_13
port 41 nsew
rlabel metal1 s 33982 1699 33982 1699 4 br_27
port 84 nsew
rlabel metal1 s 10197 1693 10197 1693 4 bl_8
port 26 nsew
rlabel metal1 s 10111 127 10111 127 4 data_8
port 25 nsew
rlabel metal1 s 23839 127 23839 127 4 data_19
port 58 nsew
rlabel metal1 s 2782 1699 2782 1699 4 br_2
port 9 nsew
rlabel metal1 s 9022 1699 9022 1699 4 br_7
port 24 nsew
rlabel metal1 s 10270 1699 10270 1699 4 br_8
port 27 nsew
rlabel metal1 s 30238 1699 30238 1699 4 br_24
port 75 nsew
rlabel metal1 s 11445 1693 11445 1693 4 bl_9
port 29 nsew
rlabel metal1 s 3871 127 3871 127 4 data_3
port 10 nsew
rlabel metal1 s 33823 127 33823 127 4 data_27
port 82 nsew
rlabel metal1 s 35157 1693 35157 1693 4 bl_28
port 86 nsew
rlabel metal1 s 13855 127 13855 127 4 data_11
port 34 nsew
rlabel metal1 s 26335 127 26335 127 4 data_21
port 64 nsew
rlabel metal1 s 37567 127 37567 127 4 data_30
port 91 nsew
rlabel metal1 s 17758 1699 17758 1699 4 br_14
port 45 nsew
rlabel metal1 s 5205 1693 5205 1693 4 bl_4
port 14 nsew
rlabel metal1 s 30079 127 30079 127 4 data_24
port 73 nsew
rlabel metal3 s 21585 1268 21585 1268 4 vdd
port 98 nsew
rlabel metal3 s 26577 1268 26577 1268 4 vdd
port 98 nsew
rlabel metal3 s 30321 1268 30321 1268 4 vdd
port 98 nsew
rlabel metal3 s 31569 1268 31569 1268 4 vdd
port 98 nsew
rlabel metal3 s 32817 1268 32817 1268 4 vdd
port 98 nsew
rlabel metal3 s 27825 1268 27825 1268 4 vdd
port 98 nsew
rlabel metal3 s 24081 1268 24081 1268 4 vdd
port 98 nsew
rlabel metal3 s 29073 1268 29073 1268 4 vdd
port 98 nsew
rlabel metal3 s 20337 1268 20337 1268 4 vdd
port 98 nsew
rlabel metal3 s 35313 1268 35313 1268 4 vdd
port 98 nsew
rlabel metal3 s 37809 1268 37809 1268 4 vdd
port 98 nsew
rlabel metal3 s 39057 1268 39057 1268 4 vdd
port 98 nsew
rlabel metal3 s 36561 1268 36561 1268 4 vdd
port 98 nsew
rlabel metal3 s 25329 1268 25329 1268 4 vdd
port 98 nsew
rlabel metal3 s 34065 1268 34065 1268 4 vdd
port 98 nsew
rlabel metal3 s 22833 1268 22833 1268 4 vdd
port 98 nsew
rlabel metal3 s 19968 2194 19968 2194 4 en
port 97 nsew
rlabel metal3 s 22915 2042 22915 2042 4 gnd
port 99 nsew
rlabel metal3 s 35395 2042 35395 2042 4 gnd
port 99 nsew
rlabel metal3 s 39139 2042 39139 2042 4 gnd
port 99 nsew
rlabel metal3 s 37891 2042 37891 2042 4 gnd
port 99 nsew
rlabel metal3 s 27907 2042 27907 2042 4 gnd
port 99 nsew
rlabel metal3 s 30403 2042 30403 2042 4 gnd
port 99 nsew
rlabel metal3 s 31651 2042 31651 2042 4 gnd
port 99 nsew
rlabel metal3 s 24163 2042 24163 2042 4 gnd
port 99 nsew
rlabel metal3 s 34147 2042 34147 2042 4 gnd
port 99 nsew
rlabel metal3 s 32899 2042 32899 2042 4 gnd
port 99 nsew
rlabel metal3 s 29155 2042 29155 2042 4 gnd
port 99 nsew
rlabel metal3 s 36643 2042 36643 2042 4 gnd
port 99 nsew
rlabel metal3 s 21667 2042 21667 2042 4 gnd
port 99 nsew
rlabel metal3 s 25411 2042 25411 2042 4 gnd
port 99 nsew
rlabel metal3 s 20419 2042 20419 2042 4 gnd
port 99 nsew
rlabel metal3 s 26659 2042 26659 2042 4 gnd
port 99 nsew
rlabel metal3 s 29085 430 29085 430 4 vdd
port 98 nsew
rlabel metal3 s 22845 430 22845 430 4 vdd
port 98 nsew
rlabel metal3 s 27837 430 27837 430 4 vdd
port 98 nsew
rlabel metal3 s 30333 430 30333 430 4 vdd
port 98 nsew
rlabel metal3 s 31581 430 31581 430 4 vdd
port 98 nsew
rlabel metal3 s 34077 430 34077 430 4 vdd
port 98 nsew
rlabel metal3 s 35325 430 35325 430 4 vdd
port 98 nsew
rlabel metal3 s 26589 430 26589 430 4 vdd
port 98 nsew
rlabel metal3 s 39069 430 39069 430 4 vdd
port 98 nsew
rlabel metal3 s 25341 430 25341 430 4 vdd
port 98 nsew
rlabel metal3 s 24093 430 24093 430 4 vdd
port 98 nsew
rlabel metal3 s 32829 430 32829 430 4 vdd
port 98 nsew
rlabel metal3 s 36573 430 36573 430 4 vdd
port 98 nsew
rlabel metal3 s 21597 430 21597 430 4 vdd
port 98 nsew
rlabel metal3 s 37821 430 37821 430 4 vdd
port 98 nsew
rlabel metal3 s 20349 430 20349 430 4 vdd
port 98 nsew
rlabel metal3 s 5361 1268 5361 1268 4 vdd
port 98 nsew
rlabel metal3 s 17841 1268 17841 1268 4 vdd
port 98 nsew
rlabel metal3 s 10353 1268 10353 1268 4 vdd
port 98 nsew
rlabel metal3 s 7939 2042 7939 2042 4 gnd
port 99 nsew
rlabel metal3 s 15345 1268 15345 1268 4 vdd
port 98 nsew
rlabel metal3 s 9187 2042 9187 2042 4 gnd
port 99 nsew
rlabel metal3 s 11601 1268 11601 1268 4 vdd
port 98 nsew
rlabel metal3 s 10435 2042 10435 2042 4 gnd
port 99 nsew
rlabel metal3 s 19171 2042 19171 2042 4 gnd
port 99 nsew
rlabel metal3 s 4195 2042 4195 2042 4 gnd
port 99 nsew
rlabel metal3 s 7857 1268 7857 1268 4 vdd
port 98 nsew
rlabel metal3 s 12849 1268 12849 1268 4 vdd
port 98 nsew
rlabel metal3 s 5443 2042 5443 2042 4 gnd
port 99 nsew
rlabel metal3 s 4113 1268 4113 1268 4 vdd
port 98 nsew
rlabel metal3 s 12931 2042 12931 2042 4 gnd
port 99 nsew
rlabel metal3 s 14179 2042 14179 2042 4 gnd
port 99 nsew
rlabel metal3 s 19101 430 19101 430 4 vdd
port 98 nsew
rlabel metal3 s 12861 430 12861 430 4 vdd
port 98 nsew
rlabel metal3 s 17853 430 17853 430 4 vdd
port 98 nsew
rlabel metal3 s 10365 430 10365 430 4 vdd
port 98 nsew
rlabel metal3 s 5373 430 5373 430 4 vdd
port 98 nsew
rlabel metal3 s 9117 430 9117 430 4 vdd
port 98 nsew
rlabel metal3 s 15357 430 15357 430 4 vdd
port 98 nsew
rlabel metal3 s 11613 430 11613 430 4 vdd
port 98 nsew
rlabel metal3 s 2877 430 2877 430 4 vdd
port 98 nsew
rlabel metal3 s 7869 430 7869 430 4 vdd
port 98 nsew
rlabel metal3 s 1629 430 1629 430 4 vdd
port 98 nsew
rlabel metal3 s 6621 430 6621 430 4 vdd
port 98 nsew
rlabel metal3 s 14109 430 14109 430 4 vdd
port 98 nsew
rlabel metal3 s 16605 430 16605 430 4 vdd
port 98 nsew
rlabel metal3 s 381 430 381 430 4 vdd
port 98 nsew
rlabel metal3 s 4125 430 4125 430 4 vdd
port 98 nsew
rlabel metal3 s 15427 2042 15427 2042 4 gnd
port 99 nsew
rlabel metal3 s 11683 2042 11683 2042 4 gnd
port 99 nsew
rlabel metal3 s 1617 1268 1617 1268 4 vdd
port 98 nsew
rlabel metal3 s 9105 1268 9105 1268 4 vdd
port 98 nsew
rlabel metal3 s 6691 2042 6691 2042 4 gnd
port 99 nsew
rlabel metal3 s 1699 2042 1699 2042 4 gnd
port 99 nsew
rlabel metal3 s 369 1268 369 1268 4 vdd
port 98 nsew
rlabel metal3 s 14097 1268 14097 1268 4 vdd
port 98 nsew
rlabel metal3 s 6609 1268 6609 1268 4 vdd
port 98 nsew
rlabel metal3 s 19089 1268 19089 1268 4 vdd
port 98 nsew
rlabel metal3 s 451 2042 451 2042 4 gnd
port 99 nsew
rlabel metal3 s 17923 2042 17923 2042 4 gnd
port 99 nsew
rlabel metal3 s 2947 2042 2947 2042 4 gnd
port 99 nsew
rlabel metal3 s 16593 1268 16593 1268 4 vdd
port 98 nsew
rlabel metal3 s 16675 2042 16675 2042 4 gnd
port 99 nsew
rlabel metal3 s 2865 1268 2865 1268 4 vdd
port 98 nsew
rlabel metal3 s 1629 108 1629 108 4 gnd
port 99 nsew
rlabel metal3 s 4125 108 4125 108 4 gnd
port 99 nsew
rlabel metal3 s 381 108 381 108 4 gnd
port 99 nsew
rlabel metal3 s 5373 108 5373 108 4 gnd
port 99 nsew
rlabel metal3 s 14109 108 14109 108 4 gnd
port 99 nsew
rlabel metal3 s 12861 108 12861 108 4 gnd
port 99 nsew
rlabel metal3 s 15357 108 15357 108 4 gnd
port 99 nsew
rlabel metal3 s 16605 108 16605 108 4 gnd
port 99 nsew
rlabel metal3 s 19101 108 19101 108 4 gnd
port 99 nsew
rlabel metal3 s 2877 108 2877 108 4 gnd
port 99 nsew
rlabel metal3 s 17853 108 17853 108 4 gnd
port 99 nsew
rlabel metal3 s 9117 108 9117 108 4 gnd
port 99 nsew
rlabel metal3 s 10365 108 10365 108 4 gnd
port 99 nsew
rlabel metal3 s 6621 108 6621 108 4 gnd
port 99 nsew
rlabel metal3 s 11613 108 11613 108 4 gnd
port 99 nsew
rlabel metal3 s 7869 108 7869 108 4 gnd
port 99 nsew
rlabel metal3 s 21597 108 21597 108 4 gnd
port 99 nsew
rlabel metal3 s 27837 108 27837 108 4 gnd
port 99 nsew
rlabel metal3 s 37821 108 37821 108 4 gnd
port 99 nsew
rlabel metal3 s 31581 108 31581 108 4 gnd
port 99 nsew
rlabel metal3 s 35325 108 35325 108 4 gnd
port 99 nsew
rlabel metal3 s 29085 108 29085 108 4 gnd
port 99 nsew
rlabel metal3 s 39069 108 39069 108 4 gnd
port 99 nsew
rlabel metal3 s 25341 108 25341 108 4 gnd
port 99 nsew
rlabel metal3 s 34077 108 34077 108 4 gnd
port 99 nsew
rlabel metal3 s 24093 108 24093 108 4 gnd
port 99 nsew
rlabel metal3 s 22845 108 22845 108 4 gnd
port 99 nsew
rlabel metal3 s 36573 108 36573 108 4 gnd
port 99 nsew
rlabel metal3 s 30333 108 30333 108 4 gnd
port 99 nsew
rlabel metal3 s 32829 108 32829 108 4 gnd
port 99 nsew
rlabel metal3 s 26589 108 26589 108 4 gnd
port 99 nsew
rlabel metal3 s 20349 108 20349 108 4 gnd
port 99 nsew
<< properties >>
string FIXED_BBOX 0 0 39936 2256
string GDS_END 3453270
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sram_1rw1r_32_256_8_sky130.gds
string GDS_START 3403286
<< end >>
