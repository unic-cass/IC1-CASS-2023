magic
tech sky130B
magscale 1 2
timestamp 1676037725
<< metal1 >>
rect 115 1333 1048 1426
rect 115 1269 984 1333
tri 984 1269 1048 1333 nw
tri 1048 1269 1073 1294 se
rect 1073 1269 2061 1294
rect 115 1230 945 1269
tri 945 1230 984 1269 nw
tri 1009 1230 1048 1269 se
rect 1048 1254 2061 1269
rect 1048 1236 1073 1254
tri 1073 1236 1091 1254 nw
rect 1048 1230 1067 1236
tri 1067 1230 1073 1236 nw
tri 981 1202 1009 1230 se
rect 1009 1202 1039 1230
tri 1039 1202 1067 1230 nw
tri 2028 1221 2061 1254 ne
tri 1086 1202 1102 1218 se
rect 1102 1202 1163 1218
rect 258 1162 999 1202
tri 999 1162 1039 1202 nw
tri 258 1156 264 1162 nw
tri 1040 1156 1086 1202 se
rect 1086 1172 1163 1202
rect 1086 1156 1129 1172
tri 1018 1134 1040 1156 se
rect 1040 1134 1129 1156
tri 1129 1140 1161 1172 nw
tri 53 1099 80 1126 se
rect 80 1099 326 1126
rect 53 1080 326 1099
rect 1165 1090 2125 1136
rect 53 403 99 1080
tri 99 1046 133 1080 nw
tri 2045 1056 2079 1090 ne
tri 532 1012 563 1043 se
rect 563 1012 1019 1043
tri 1019 1012 1050 1043 sw
tri 489 969 532 1012 se
rect 532 997 1050 1012
rect 532 969 555 997
tri 555 969 583 997 nw
rect 275 938 524 969
tri 524 938 555 969 nw
tri 564 938 595 969 se
rect 595 946 972 969
tri 972 946 995 969 sw
tri 999 946 1050 997 ne
tri 1050 946 1116 1012 sw
rect 595 938 995 946
rect 275 923 509 938
tri 509 923 524 938 nw
tri 549 923 564 938 se
rect 564 923 995 938
tri 519 893 549 923 se
rect 549 893 564 923
rect 343 872 564 893
tri 564 872 615 923 nw
tri 952 903 972 923 ne
rect 972 911 995 923
tri 995 911 1030 946 sw
tri 1050 911 1085 946 ne
rect 1085 911 1496 946
rect 972 903 1030 911
rect 343 765 515 872
tri 515 823 564 872 nw
tri 972 845 1030 903 ne
tri 1030 872 1069 911 sw
tri 1085 900 1096 911 ne
rect 1096 900 1496 911
tri 2040 872 2079 911 se
rect 2079 891 2125 1090
tri 2125 1056 2159 1090 nw
rect 2079 872 2106 891
tri 2106 872 2125 891 nw
rect 1030 845 2064 872
tri 687 811 721 845 sw
tri 779 811 813 845 se
tri 859 811 893 845 sw
tri 1030 830 1045 845 ne
rect 1045 830 2064 845
tri 2064 830 2106 872 nw
rect 343 763 513 765
tri 513 763 515 765 nw
rect 641 801 1023 811
tri 1023 801 1033 811 sw
rect 641 763 1257 801
tri 1005 755 1013 763 ne
rect 1013 755 1257 763
rect 150 605 899 735
rect 150 440 196 605
tri 196 563 238 605 nw
rect 267 529 550 575
rect 1018 530 1500 576
tri 297 523 303 529 ne
tri 1466 496 1500 530 ne
tri 196 440 216 460 sw
tri 53 357 99 403 ne
tri 99 374 148 423 sw
tri 150 374 216 440 ne
tri 216 376 280 440 sw
rect 216 374 810 376
rect 99 367 148 374
tri 148 367 155 374 sw
rect 99 357 155 367
tri 99 301 155 357 ne
tri 155 330 192 367 sw
tri 216 330 260 374 ne
rect 260 330 810 374
rect 155 301 192 330
tri 192 301 221 330 sw
tri 1341 301 1425 385 se
tri 1905 345 1936 376 se
rect 1936 356 1982 417
rect 1936 345 1960 356
tri 155 255 201 301 ne
rect 201 255 1425 301
rect 1834 334 1960 345
tri 1960 334 1982 356 nw
rect 1834 299 1925 334
tri 1925 299 1960 334 nw
tri 2027 300 2061 334 se
tri 2113 300 2140 327 sw
use sky130_fd_pr__nfet_01v8__example_55959141808463  sky130_fd_pr__nfet_01v8__example_55959141808463_0
timestamp 1676037725
transform 1 0 736 0 1 163
box -1 0 569 1
use sky130_fd_pr__nfet_01v8__example_55959141808464  sky130_fd_pr__nfet_01v8__example_55959141808464_0
timestamp 1676037725
transform -1 0 2110 0 -1 1288
box -1 0 889 1
use sky130_fd_pr__nfet_01v8__example_55959141808465  sky130_fd_pr__nfet_01v8__example_55959141808465_0
timestamp 1676037725
transform 1 0 1632 0 -1 363
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808465  sky130_fd_pr__nfet_01v8__example_55959141808465_1
timestamp 1676037725
transform -1 0 1576 0 -1 363
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808465  sky130_fd_pr__nfet_01v8__example_55959141808465_2
timestamp 1676037725
transform 1 0 1911 0 -1 363
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808466  sky130_fd_pr__nfet_01v8__example_55959141808466_0
timestamp 1676037725
transform -1 0 550 0 -1 817
box -1 0 289 1
use sky130_fd_pr__nfet_01v8__example_55959141808467  sky130_fd_pr__nfet_01v8__example_55959141808467_0
timestamp 1676037725
transform -1 0 894 0 -1 817
box -1 0 289 1
use sky130_fd_pr__nfet_01v8__example_55959141808468  sky130_fd_pr__nfet_01v8__example_55959141808468_0
timestamp 1676037725
transform -1 0 2110 0 1 758
box -1 0 889 1
use sky130_fd_pr__pfet_01v8__example_55959141808460  sky130_fd_pr__pfet_01v8__example_55959141808460_0
timestamp 1676037725
transform 1 0 863 0 -1 1297
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808460  sky130_fd_pr__pfet_01v8__example_55959141808460_1
timestamp 1676037725
transform 1 0 597 0 -1 1297
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808590  sky130_fd_pr__pfet_01v8__example_55959141808590_0
timestamp 1676037725
transform 1 0 331 0 -1 1297
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808590  sky130_fd_pr__pfet_01v8__example_55959141808590_1
timestamp 1676037725
transform -1 0 275 0 -1 1297
box -1 0 101 1
<< properties >>
string GDS_END 43785774
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 43756086
<< end >>
