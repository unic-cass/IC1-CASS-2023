magic
tech sky130A
magscale 1 2
timestamp 1676037725
<< poly >>
rect 12348 -90 12535 -57
rect 12348 -124 12365 -90
rect 12399 -124 12433 -90
rect 12467 -124 12501 -90
rect 12348 -157 12535 -124
rect 14575 -90 14762 -57
rect 14609 -124 14643 -90
rect 14677 -124 14711 -90
rect 14745 -124 14762 -90
rect 14575 -157 14762 -124
<< polycont >>
rect 12365 -124 12399 -90
rect 12433 -124 12467 -90
rect 12501 -124 12535 -90
rect 14575 -124 14609 -90
rect 14643 -124 14677 -90
rect 14711 -124 14745 -90
<< npolyres >>
rect 12535 -157 14575 -57
<< locali >>
rect 9117 215 9175 249
rect 9209 215 9267 249
rect 9083 175 9301 215
rect 9117 141 9175 175
rect 9209 141 9267 175
rect 9083 101 9301 141
rect 9117 67 9175 101
rect 9209 67 9267 101
rect 9083 27 9301 67
rect 9117 -7 9175 27
rect 9209 -7 9267 27
rect 9083 -47 9301 -7
rect 9117 -81 9175 -47
rect 9209 -81 9267 -47
rect 14559 -43 14761 -37
rect 9083 -121 9301 -81
rect 9117 -155 9175 -121
rect 9209 -155 9267 -121
rect 12349 -90 12551 -74
rect 12349 -100 12365 -90
rect 12349 -134 12362 -100
rect 12399 -124 12433 -90
rect 12467 -100 12501 -90
rect 12535 -94 12551 -90
rect 14559 -77 14571 -43
rect 14605 -77 14643 -43
rect 14677 -77 14715 -43
rect 14749 -77 14761 -43
rect 14559 -90 14761 -77
rect 12535 -100 12552 -94
rect 12468 -124 12501 -100
rect 12396 -134 12434 -124
rect 12468 -134 12506 -124
rect 12540 -134 12552 -100
rect 12349 -140 12552 -134
rect 14559 -124 14575 -90
rect 14609 -124 14643 -90
rect 14677 -124 14711 -90
rect 14745 -124 14761 -90
rect 14559 -125 14761 -124
rect 14559 -159 14571 -125
rect 14605 -159 14643 -125
rect 14677 -159 14715 -125
rect 14749 -159 14761 -125
rect 14559 -165 14761 -159
<< viali >>
rect 9083 215 9117 249
rect 9175 215 9209 249
rect 9267 215 9301 249
rect 9083 141 9117 175
rect 9175 141 9209 175
rect 9267 141 9301 175
rect 9083 67 9117 101
rect 9175 67 9209 101
rect 9267 67 9301 101
rect 9083 -7 9117 27
rect 9175 -7 9209 27
rect 9267 -7 9301 27
rect 9083 -81 9117 -47
rect 9175 -81 9209 -47
rect 9267 -81 9301 -47
rect 9083 -155 9117 -121
rect 9175 -155 9209 -121
rect 9267 -155 9301 -121
rect 12362 -124 12365 -100
rect 12365 -124 12396 -100
rect 14571 -77 14605 -43
rect 14643 -77 14677 -43
rect 14715 -77 14749 -43
rect 12434 -124 12467 -100
rect 12467 -124 12468 -100
rect 12506 -124 12535 -100
rect 12535 -124 12540 -100
rect 12362 -134 12396 -124
rect 12434 -134 12468 -124
rect 12506 -134 12540 -124
rect 14571 -159 14605 -125
rect 14643 -159 14677 -125
rect 14715 -159 14749 -125
<< metal1 >>
rect 1427 1478 2325 1608
rect 2455 1478 2755 1608
rect 2885 1602 3863 1608
rect 2885 1550 3733 1602
rect 3785 1550 3811 1602
rect 2885 1536 3863 1550
rect 2885 1484 3733 1536
rect 3785 1484 3811 1536
rect 2885 1478 3863 1484
rect 4439 1478 5301 1608
rect 5431 1478 7285 1608
rect 7367 1556 8282 1608
rect 8334 1556 8349 1608
rect 8401 1556 8407 1608
rect 7367 1530 8407 1556
rect 7367 1478 8282 1530
rect 8334 1478 8349 1530
rect 8401 1478 8407 1530
rect 8837 1562 9733 1608
rect 8837 1510 9132 1562
rect 9184 1510 9199 1562
rect 9251 1510 9267 1562
rect 9319 1510 9335 1562
rect 9387 1510 9403 1562
rect 9455 1510 9471 1562
rect 9523 1510 9539 1562
rect 9591 1510 9607 1562
rect 9659 1510 9675 1562
rect 9727 1510 9733 1562
rect 8837 1479 9733 1510
rect 10391 1556 10950 1608
rect 11002 1556 11025 1608
rect 11077 1556 11100 1608
rect 11152 1556 11175 1608
rect 11227 1556 11250 1608
rect 11302 1556 11325 1608
rect 11377 1556 11383 1608
rect 10391 1530 11383 1556
rect 8837 1478 9699 1479
rect 10391 1478 10950 1530
rect 11002 1478 11025 1530
rect 11077 1478 11100 1530
rect 11152 1478 11175 1530
rect 11227 1478 11250 1530
rect 11302 1478 11325 1530
rect 11377 1478 11383 1530
rect 11745 1556 12371 1608
rect 12423 1556 12441 1608
rect 12493 1556 12511 1608
rect 12563 1556 12581 1608
rect 12633 1556 12651 1608
rect 12703 1556 12709 1608
rect 11745 1530 12709 1556
rect 11745 1478 12371 1530
rect 12423 1478 12441 1530
rect 12493 1478 12511 1530
rect 12563 1478 12581 1530
rect 12633 1478 12651 1530
rect 12703 1478 12709 1530
rect 13237 1601 13367 1608
rect 13237 1549 13243 1601
rect 13295 1549 13309 1601
rect 13361 1549 13367 1601
rect 13237 1537 13367 1549
rect 13237 1485 13243 1537
rect 13295 1485 13309 1537
rect 13361 1485 13367 1537
rect 13237 1478 13367 1485
rect 13667 1601 13797 1608
rect 13667 1549 13673 1601
rect 13725 1549 13739 1601
rect 13791 1549 13797 1601
rect 13667 1537 13797 1549
rect 13667 1485 13673 1537
rect 13725 1485 13739 1537
rect 13791 1485 13797 1537
rect 13667 1478 13797 1485
rect 14229 1601 14587 1608
rect 14229 1549 14235 1601
rect 14287 1549 14301 1601
rect 14353 1549 14587 1601
rect 14229 1537 14587 1549
rect 14229 1485 14235 1537
rect 14287 1485 14301 1537
rect 14353 1485 14587 1537
rect 14229 1478 14587 1485
rect 12712 661 12811 745
rect 1330 403 1336 455
rect 1388 403 1423 455
rect 1475 403 1510 455
rect 1562 403 1597 455
rect 1649 403 1684 455
rect 1736 403 1742 455
rect 1330 339 1742 403
rect 1330 287 1336 339
rect 1388 287 1423 339
rect 1475 287 1510 339
rect 1562 287 1597 339
rect 1649 287 1684 339
rect 1736 287 1742 339
rect 2410 403 2416 455
rect 2468 403 2503 455
rect 2555 403 2590 455
rect 2642 403 2677 455
rect 2729 403 2764 455
rect 2816 403 2822 455
rect 2410 339 2822 403
rect 2410 287 2416 339
rect 2468 287 2503 339
rect 2555 287 2590 339
rect 2642 287 2677 339
rect 2729 287 2764 339
rect 2816 287 2822 339
tri 3028 333 3150 455 sw
tri 6027 281 6033 287 ne
rect 6033 281 6039 333
rect 6091 281 6109 333
rect 6161 281 6179 333
rect 6231 281 6249 333
rect 6301 281 6319 333
rect 6371 281 6388 333
rect 6440 281 6457 333
rect 6509 281 6515 333
tri 6515 281 6521 287 nw
tri 6652 281 6658 287 ne
rect 6658 281 6664 333
rect 6716 281 6733 333
rect 6785 281 6802 333
rect 6854 281 6872 333
rect 6924 281 6942 333
rect 6994 281 7012 333
rect 7064 281 7082 333
rect 7134 281 7140 333
tri 7140 281 7146 287 nw
rect 9077 255 9307 261
rect 9077 203 9078 255
rect 9130 203 9166 255
rect 9218 203 9254 255
rect 9306 203 9307 255
rect 9077 183 9307 203
rect 9077 131 9078 183
rect 9130 131 9166 183
rect 9218 131 9254 183
rect 9306 131 9307 183
rect 9077 110 9307 131
tri 3418 98 3422 102 se
rect 3422 98 3429 102
rect 3423 54 3429 98
tri 3418 50 3422 54 ne
rect 3422 50 3429 54
rect 3481 50 3493 102
rect 3545 98 3552 102
tri 3552 98 3556 102 sw
rect 3545 54 3551 98
rect 9077 58 9078 110
rect 9130 58 9166 110
rect 9218 58 9254 110
rect 9306 58 9307 110
rect 12076 151 12082 203
rect 12134 151 12155 203
rect 12207 151 12227 203
rect 12279 151 14108 203
rect 12076 145 14108 151
tri 14108 145 14166 203 sw
rect 12076 123 14166 145
rect 12076 71 12082 123
rect 12134 71 12155 123
rect 12207 71 12227 123
rect 12279 71 14166 123
rect 3545 50 3552 54
tri 3552 50 3556 54 nw
rect 9077 37 9307 58
rect 1330 -31 1336 21
rect 1388 -31 1423 21
rect 1475 -31 1510 21
rect 1562 -31 1597 21
rect 1649 -31 1684 21
rect 1736 -31 1742 21
rect 1330 -45 1742 -31
rect 1330 -97 1336 -45
rect 1388 -97 1423 -45
rect 1475 -97 1510 -45
rect 1562 -97 1597 -45
rect 1649 -97 1684 -45
rect 1736 -97 1742 -45
rect 2410 -31 2416 21
rect 2468 -31 2503 21
rect 2555 -31 2590 21
rect 2642 -31 2677 21
rect 2729 -31 2764 21
rect 2816 -31 2822 21
rect 2410 -45 2822 -31
rect 2410 -97 2416 -45
rect 2468 -97 2503 -45
rect 2555 -97 2590 -45
rect 2642 -97 2677 -45
rect 2729 -97 2764 -45
rect 2816 -97 2822 -45
rect 6033 -31 6039 21
rect 6091 -31 6123 21
rect 6175 -31 6207 21
rect 6259 -31 6291 21
rect 6343 -31 6374 21
rect 6426 -31 6457 21
rect 6509 -31 6515 21
rect 6033 -45 6515 -31
rect 6033 -97 6039 -45
rect 6091 -97 6123 -45
rect 6175 -97 6207 -45
rect 6259 -97 6291 -45
rect 6343 -97 6374 -45
rect 6426 -97 6457 -45
rect 6509 -97 6515 -45
rect 6658 -31 6664 21
rect 6716 -31 6748 21
rect 6800 -31 6832 21
rect 6884 -31 6916 21
rect 6968 -31 6999 21
rect 7051 -31 7082 21
rect 7134 -31 7140 21
rect 6658 -45 7140 -31
rect 6658 -97 6664 -45
rect 6716 -97 6748 -45
rect 6800 -97 6832 -45
rect 6884 -97 6916 -45
rect 6968 -97 6999 -45
rect 7051 -97 7082 -45
rect 7134 -97 7140 -45
rect 9077 -15 9078 37
rect 9130 -15 9166 37
rect 9218 -15 9254 37
rect 9306 -15 9307 37
rect 9077 -36 9307 -15
rect 9077 -88 9078 -36
rect 9130 -88 9166 -36
rect 9218 -88 9254 -36
rect 9306 -88 9307 -36
tri 14058 -37 14166 71 ne
tri 14166 -37 14348 145 sw
rect 9077 -109 9307 -88
rect 9077 -161 9078 -109
rect 9130 -161 9166 -109
rect 9218 -161 9254 -109
rect 9306 -161 9307 -109
rect 12003 -146 12009 -94
rect 12061 -146 12073 -94
rect 12125 -100 12552 -94
rect 12125 -134 12362 -100
rect 12396 -134 12434 -100
rect 12468 -134 12506 -100
rect 12540 -134 12552 -100
rect 12125 -146 12552 -134
rect 9077 -167 9307 -161
tri 14166 -165 14294 -37 ne
rect 14294 -43 14761 -37
rect 14294 -77 14571 -43
rect 14605 -77 14643 -43
rect 14677 -77 14715 -43
rect 14749 -77 14761 -43
rect 14294 -125 14761 -77
rect 14294 -159 14571 -125
rect 14605 -159 14643 -125
rect 14677 -159 14715 -125
rect 14749 -159 14761 -125
rect 14294 -165 14761 -159
rect 1330 -343 1336 -291
rect 1388 -343 1423 -291
rect 1475 -343 1510 -291
rect 1562 -343 1597 -291
rect 1649 -343 1684 -291
rect 1736 -343 1742 -291
rect 1330 -407 1742 -343
rect 1330 -459 1336 -407
rect 1388 -459 1423 -407
rect 1475 -459 1510 -407
rect 1562 -459 1597 -407
rect 1649 -459 1684 -407
rect 1736 -459 1742 -407
rect 2410 -344 2416 -292
rect 2468 -344 2503 -292
rect 2555 -344 2590 -292
rect 2642 -344 2677 -292
rect 2729 -344 2764 -292
rect 2816 -344 2822 -292
rect 2410 -358 2822 -344
rect 2410 -410 2416 -358
rect 2468 -410 2503 -358
rect 2555 -410 2590 -358
rect 2642 -410 2677 -358
rect 2729 -410 2764 -358
rect 2816 -410 2822 -358
rect 6033 -343 6039 -291
rect 6091 -343 6109 -291
rect 6161 -343 6179 -291
rect 6231 -343 6249 -291
rect 6301 -343 6319 -291
rect 6371 -343 6388 -291
rect 6440 -343 6457 -291
rect 6509 -343 6515 -291
rect 6033 -407 6515 -343
rect 6033 -459 6039 -407
rect 6091 -459 6109 -407
rect 6161 -459 6179 -407
rect 6231 -459 6249 -407
rect 6301 -459 6319 -407
rect 6371 -459 6388 -407
rect 6440 -459 6457 -407
rect 6509 -459 6515 -407
rect 6658 -343 6664 -291
rect 6716 -343 6734 -291
rect 6786 -343 6804 -291
rect 6856 -343 6874 -291
rect 6926 -343 6944 -291
rect 6996 -343 7013 -291
rect 7065 -343 7082 -291
rect 7134 -343 7140 -291
tri 14471 -317 14498 -290 se
rect 14498 -317 14737 -290
rect 6658 -407 7140 -343
tri 8126 -391 8200 -317 se
rect 8200 -369 10681 -317
rect 10733 -369 10745 -317
rect 10797 -369 11429 -317
rect 11481 -369 11493 -317
rect 11545 -369 12856 -317
rect 12908 -369 12920 -317
rect 12972 -369 13141 -317
rect 13193 -369 13207 -317
rect 13259 -369 14082 -317
rect 14134 -369 14146 -317
rect 14198 -342 14737 -317
rect 14789 -342 14801 -290
rect 14853 -342 14865 -290
rect 14917 -342 14929 -290
rect 14981 -342 14993 -290
rect 15045 -342 15057 -290
rect 15109 -342 15115 -290
rect 14198 -369 14550 -342
tri 14550 -369 14577 -342 nw
tri 8200 -391 8222 -369 nw
tri 8115 -402 8126 -391 se
rect 8126 -402 8137 -391
rect 6658 -459 6664 -407
rect 6716 -459 6734 -407
rect 6786 -459 6804 -407
rect 6856 -459 6874 -407
rect 6926 -459 6944 -407
rect 6996 -459 7013 -407
rect 7065 -459 7082 -407
rect 7134 -459 7140 -407
rect 7755 -454 7761 -402
rect 7813 -454 7825 -402
rect 7877 -454 8137 -402
tri 8137 -454 8200 -391 nw
tri 14602 -402 14629 -375 se
rect 14629 -402 15041 -375
rect 8246 -454 8252 -402
rect 8304 -454 8360 -402
rect 8412 -454 10446 -402
rect 10498 -454 10510 -402
rect 10562 -454 11194 -402
rect 11246 -454 11258 -402
rect 11310 -454 12615 -402
rect 12667 -454 12679 -402
rect 12731 -454 13845 -402
rect 13897 -454 13909 -402
rect 13961 -454 14539 -402
rect 14591 -454 14603 -402
rect 14655 -427 15041 -402
rect 15093 -427 15106 -375
rect 15158 -427 15164 -375
rect 14655 -454 14665 -427
tri 14665 -454 14692 -427 nw
tri 14689 -482 14716 -455 se
rect 14716 -461 15094 -455
rect 14716 -482 15042 -461
rect 7755 -534 7761 -482
rect 7813 -534 7825 -482
rect 7877 -534 7883 -482
rect 9839 -534 10204 -482
rect 10256 -534 10268 -482
rect 10320 -534 10952 -482
rect 11004 -534 11016 -482
rect 11068 -534 12006 -482
rect 12058 -534 12070 -482
rect 12122 -534 12373 -482
rect 12425 -534 12437 -482
rect 12489 -534 13600 -482
rect 13652 -534 13664 -482
rect 13716 -534 14294 -482
rect 14346 -534 14358 -482
rect 14410 -507 15042 -482
rect 14410 -534 14893 -507
tri 14893 -534 14920 -507 nw
tri 7797 -568 7831 -534 ne
rect 7831 -658 7883 -534
tri 14998 -551 15042 -507 ne
rect 15042 -525 15094 -513
rect 14880 -614 14886 -562
rect 14938 -614 14950 -562
rect 15002 -614 15008 -562
rect 15042 -583 15094 -577
tri 7831 -710 7883 -658 ne
tri 7883 -710 7957 -636 sw
tri 14316 -710 14383 -643 se
rect 14383 -695 14806 -643
rect 14858 -695 14870 -643
rect 14922 -695 14928 -643
rect 14383 -710 14390 -695
tri 14390 -710 14405 -695 nw
tri 7883 -762 7935 -710 ne
rect 7935 -762 14338 -710
tri 14338 -762 14390 -710 nw
<< via1 >>
rect 3733 1550 3785 1602
rect 3811 1550 3863 1602
rect 3733 1484 3785 1536
rect 3811 1484 3863 1536
rect 8282 1556 8334 1608
rect 8349 1556 8401 1608
rect 8282 1478 8334 1530
rect 8349 1478 8401 1530
rect 9132 1510 9184 1562
rect 9199 1510 9251 1562
rect 9267 1510 9319 1562
rect 9335 1510 9387 1562
rect 9403 1510 9455 1562
rect 9471 1510 9523 1562
rect 9539 1510 9591 1562
rect 9607 1510 9659 1562
rect 9675 1510 9727 1562
rect 10950 1556 11002 1608
rect 11025 1556 11077 1608
rect 11100 1556 11152 1608
rect 11175 1556 11227 1608
rect 11250 1556 11302 1608
rect 11325 1556 11377 1608
rect 10950 1478 11002 1530
rect 11025 1478 11077 1530
rect 11100 1478 11152 1530
rect 11175 1478 11227 1530
rect 11250 1478 11302 1530
rect 11325 1478 11377 1530
rect 12371 1556 12423 1608
rect 12441 1556 12493 1608
rect 12511 1556 12563 1608
rect 12581 1556 12633 1608
rect 12651 1556 12703 1608
rect 12371 1478 12423 1530
rect 12441 1478 12493 1530
rect 12511 1478 12563 1530
rect 12581 1478 12633 1530
rect 12651 1478 12703 1530
rect 13243 1549 13295 1601
rect 13309 1549 13361 1601
rect 13243 1485 13295 1537
rect 13309 1485 13361 1537
rect 13673 1549 13725 1601
rect 13739 1549 13791 1601
rect 13673 1485 13725 1537
rect 13739 1485 13791 1537
rect 14235 1549 14287 1601
rect 14301 1549 14353 1601
rect 14235 1485 14287 1537
rect 14301 1485 14353 1537
rect 1336 403 1388 455
rect 1423 403 1475 455
rect 1510 403 1562 455
rect 1597 403 1649 455
rect 1684 403 1736 455
rect 1336 287 1388 339
rect 1423 287 1475 339
rect 1510 287 1562 339
rect 1597 287 1649 339
rect 1684 287 1736 339
rect 2416 403 2468 455
rect 2503 403 2555 455
rect 2590 403 2642 455
rect 2677 403 2729 455
rect 2764 403 2816 455
rect 2416 287 2468 339
rect 2503 287 2555 339
rect 2590 287 2642 339
rect 2677 287 2729 339
rect 2764 287 2816 339
rect 6039 281 6091 333
rect 6109 281 6161 333
rect 6179 281 6231 333
rect 6249 281 6301 333
rect 6319 281 6371 333
rect 6388 281 6440 333
rect 6457 281 6509 333
rect 6664 281 6716 333
rect 6733 281 6785 333
rect 6802 281 6854 333
rect 6872 281 6924 333
rect 6942 281 6994 333
rect 7012 281 7064 333
rect 7082 281 7134 333
rect 9078 249 9130 255
rect 9078 215 9083 249
rect 9083 215 9117 249
rect 9117 215 9130 249
rect 9078 203 9130 215
rect 9166 249 9218 255
rect 9166 215 9175 249
rect 9175 215 9209 249
rect 9209 215 9218 249
rect 9166 203 9218 215
rect 9254 249 9306 255
rect 9254 215 9267 249
rect 9267 215 9301 249
rect 9301 215 9306 249
rect 9254 203 9306 215
rect 9078 175 9130 183
rect 9078 141 9083 175
rect 9083 141 9117 175
rect 9117 141 9130 175
rect 9078 131 9130 141
rect 9166 175 9218 183
rect 9166 141 9175 175
rect 9175 141 9209 175
rect 9209 141 9218 175
rect 9166 131 9218 141
rect 9254 175 9306 183
rect 9254 141 9267 175
rect 9267 141 9301 175
rect 9301 141 9306 175
rect 9254 131 9306 141
rect 3429 50 3481 102
rect 3493 50 3545 102
rect 9078 101 9130 110
rect 9078 67 9083 101
rect 9083 67 9117 101
rect 9117 67 9130 101
rect 9078 58 9130 67
rect 9166 101 9218 110
rect 9166 67 9175 101
rect 9175 67 9209 101
rect 9209 67 9218 101
rect 9166 58 9218 67
rect 9254 101 9306 110
rect 9254 67 9267 101
rect 9267 67 9301 101
rect 9301 67 9306 101
rect 9254 58 9306 67
rect 12082 151 12134 203
rect 12155 151 12207 203
rect 12227 151 12279 203
rect 12082 71 12134 123
rect 12155 71 12207 123
rect 12227 71 12279 123
rect 1336 -31 1388 21
rect 1423 -31 1475 21
rect 1510 -31 1562 21
rect 1597 -31 1649 21
rect 1684 -31 1736 21
rect 1336 -97 1388 -45
rect 1423 -97 1475 -45
rect 1510 -97 1562 -45
rect 1597 -97 1649 -45
rect 1684 -97 1736 -45
rect 2416 -31 2468 21
rect 2503 -31 2555 21
rect 2590 -31 2642 21
rect 2677 -31 2729 21
rect 2764 -31 2816 21
rect 2416 -97 2468 -45
rect 2503 -97 2555 -45
rect 2590 -97 2642 -45
rect 2677 -97 2729 -45
rect 2764 -97 2816 -45
rect 6039 -31 6091 21
rect 6123 -31 6175 21
rect 6207 -31 6259 21
rect 6291 -31 6343 21
rect 6374 -31 6426 21
rect 6457 -31 6509 21
rect 6039 -97 6091 -45
rect 6123 -97 6175 -45
rect 6207 -97 6259 -45
rect 6291 -97 6343 -45
rect 6374 -97 6426 -45
rect 6457 -97 6509 -45
rect 6664 -31 6716 21
rect 6748 -31 6800 21
rect 6832 -31 6884 21
rect 6916 -31 6968 21
rect 6999 -31 7051 21
rect 7082 -31 7134 21
rect 6664 -97 6716 -45
rect 6748 -97 6800 -45
rect 6832 -97 6884 -45
rect 6916 -97 6968 -45
rect 6999 -97 7051 -45
rect 7082 -97 7134 -45
rect 9078 27 9130 37
rect 9078 -7 9083 27
rect 9083 -7 9117 27
rect 9117 -7 9130 27
rect 9078 -15 9130 -7
rect 9166 27 9218 37
rect 9166 -7 9175 27
rect 9175 -7 9209 27
rect 9209 -7 9218 27
rect 9166 -15 9218 -7
rect 9254 27 9306 37
rect 9254 -7 9267 27
rect 9267 -7 9301 27
rect 9301 -7 9306 27
rect 9254 -15 9306 -7
rect 9078 -47 9130 -36
rect 9078 -81 9083 -47
rect 9083 -81 9117 -47
rect 9117 -81 9130 -47
rect 9078 -88 9130 -81
rect 9166 -47 9218 -36
rect 9166 -81 9175 -47
rect 9175 -81 9209 -47
rect 9209 -81 9218 -47
rect 9166 -88 9218 -81
rect 9254 -47 9306 -36
rect 9254 -81 9267 -47
rect 9267 -81 9301 -47
rect 9301 -81 9306 -47
rect 9254 -88 9306 -81
rect 9078 -121 9130 -109
rect 9078 -155 9083 -121
rect 9083 -155 9117 -121
rect 9117 -155 9130 -121
rect 9078 -161 9130 -155
rect 9166 -121 9218 -109
rect 9166 -155 9175 -121
rect 9175 -155 9209 -121
rect 9209 -155 9218 -121
rect 9166 -161 9218 -155
rect 9254 -121 9306 -109
rect 9254 -155 9267 -121
rect 9267 -155 9301 -121
rect 9301 -155 9306 -121
rect 9254 -161 9306 -155
rect 12009 -146 12061 -94
rect 12073 -146 12125 -94
rect 1336 -343 1388 -291
rect 1423 -343 1475 -291
rect 1510 -343 1562 -291
rect 1597 -343 1649 -291
rect 1684 -343 1736 -291
rect 1336 -459 1388 -407
rect 1423 -459 1475 -407
rect 1510 -459 1562 -407
rect 1597 -459 1649 -407
rect 1684 -459 1736 -407
rect 2416 -344 2468 -292
rect 2503 -344 2555 -292
rect 2590 -344 2642 -292
rect 2677 -344 2729 -292
rect 2764 -344 2816 -292
rect 2416 -410 2468 -358
rect 2503 -410 2555 -358
rect 2590 -410 2642 -358
rect 2677 -410 2729 -358
rect 2764 -410 2816 -358
rect 6039 -343 6091 -291
rect 6109 -343 6161 -291
rect 6179 -343 6231 -291
rect 6249 -343 6301 -291
rect 6319 -343 6371 -291
rect 6388 -343 6440 -291
rect 6457 -343 6509 -291
rect 6039 -459 6091 -407
rect 6109 -459 6161 -407
rect 6179 -459 6231 -407
rect 6249 -459 6301 -407
rect 6319 -459 6371 -407
rect 6388 -459 6440 -407
rect 6457 -459 6509 -407
rect 6664 -343 6716 -291
rect 6734 -343 6786 -291
rect 6804 -343 6856 -291
rect 6874 -343 6926 -291
rect 6944 -343 6996 -291
rect 7013 -343 7065 -291
rect 7082 -343 7134 -291
rect 10681 -369 10733 -317
rect 10745 -369 10797 -317
rect 11429 -369 11481 -317
rect 11493 -369 11545 -317
rect 12856 -369 12908 -317
rect 12920 -369 12972 -317
rect 13141 -369 13193 -317
rect 13207 -369 13259 -317
rect 14082 -369 14134 -317
rect 14146 -369 14198 -317
rect 14737 -342 14789 -290
rect 14801 -342 14853 -290
rect 14865 -342 14917 -290
rect 14929 -342 14981 -290
rect 14993 -342 15045 -290
rect 15057 -342 15109 -290
rect 6664 -459 6716 -407
rect 6734 -459 6786 -407
rect 6804 -459 6856 -407
rect 6874 -459 6926 -407
rect 6944 -459 6996 -407
rect 7013 -459 7065 -407
rect 7082 -459 7134 -407
rect 7761 -454 7813 -402
rect 7825 -454 7877 -402
rect 8252 -454 8304 -402
rect 8360 -454 8412 -402
rect 10446 -454 10498 -402
rect 10510 -454 10562 -402
rect 11194 -454 11246 -402
rect 11258 -454 11310 -402
rect 12615 -454 12667 -402
rect 12679 -454 12731 -402
rect 13845 -454 13897 -402
rect 13909 -454 13961 -402
rect 14539 -454 14591 -402
rect 14603 -454 14655 -402
rect 15041 -427 15093 -375
rect 15106 -427 15158 -375
rect 7761 -534 7813 -482
rect 7825 -534 7877 -482
rect 10204 -534 10256 -482
rect 10268 -534 10320 -482
rect 10952 -534 11004 -482
rect 11016 -534 11068 -482
rect 12006 -534 12058 -482
rect 12070 -534 12122 -482
rect 12373 -534 12425 -482
rect 12437 -534 12489 -482
rect 13600 -534 13652 -482
rect 13664 -534 13716 -482
rect 14294 -534 14346 -482
rect 14358 -534 14410 -482
rect 15042 -513 15094 -461
rect 14886 -614 14938 -562
rect 14950 -614 15002 -562
rect 15042 -577 15094 -525
rect 14806 -695 14858 -643
rect 14870 -695 14922 -643
<< metal2 >>
rect 11366 3389 13325 4498
rect 13565 1988 14578 2981
rect 3733 1602 3863 1608
rect 3785 1550 3811 1602
rect 3733 1536 3863 1550
rect 3785 1484 3811 1536
rect 1330 403 1336 455
rect 1388 403 1423 455
rect 1475 403 1510 455
rect 1562 403 1597 455
rect 1649 403 1684 455
rect 1736 403 1742 455
rect 1330 339 1742 403
rect 1330 287 1336 339
rect 1388 287 1423 339
rect 1475 287 1510 339
rect 1562 287 1597 339
rect 1649 287 1684 339
rect 1736 287 1742 339
rect 1330 21 1742 287
rect 1330 -31 1336 21
rect 1388 -31 1423 21
rect 1475 -31 1510 21
rect 1562 -31 1597 21
rect 1649 -31 1684 21
rect 1736 -31 1742 21
rect 1330 -45 1742 -31
rect 1330 -97 1336 -45
rect 1388 -97 1423 -45
rect 1475 -97 1510 -45
rect 1562 -97 1597 -45
rect 1649 -97 1684 -45
rect 1736 -97 1742 -45
rect 1330 -291 1742 -97
rect 1330 -343 1336 -291
rect 1388 -343 1423 -291
rect 1475 -343 1510 -291
rect 1562 -343 1597 -291
rect 1649 -343 1684 -291
rect 1736 -343 1742 -291
rect 1330 -407 1742 -343
rect 1330 -459 1336 -407
rect 1388 -459 1423 -407
rect 1475 -459 1510 -407
rect 1562 -459 1597 -407
rect 1649 -459 1684 -407
rect 1736 -459 1742 -407
rect 2410 403 2416 455
rect 2468 403 2503 455
rect 2555 403 2590 455
rect 2642 403 2677 455
rect 2729 403 2764 455
rect 2816 403 2822 455
rect 2410 339 2822 403
rect 2410 287 2416 339
rect 2468 287 2503 339
rect 2555 287 2590 339
rect 2642 287 2677 339
rect 2729 287 2764 339
rect 2816 287 2822 339
rect 2410 21 2822 287
rect 3423 50 3429 102
rect 3481 50 3493 102
rect 3545 50 3551 102
rect 2410 -31 2416 21
rect 2468 -31 2503 21
rect 2555 -31 2590 21
rect 2642 -31 2677 21
rect 2729 -31 2764 21
rect 2816 -31 2822 21
tri 3438 16 3472 50 ne
rect 2410 -45 2822 -31
rect 2410 -97 2416 -45
rect 2468 -97 2503 -45
rect 2555 -97 2590 -45
rect 2642 -97 2677 -45
rect 2729 -97 2764 -45
rect 2816 -97 2822 -45
rect 2410 -292 2822 -97
rect 2410 -344 2416 -292
rect 2468 -344 2503 -292
rect 2555 -344 2590 -292
rect 2642 -344 2677 -292
rect 2729 -344 2764 -292
rect 2816 -344 2822 -292
rect 2410 -358 2822 -344
rect 2410 -410 2416 -358
rect 2468 -410 2503 -358
rect 2555 -410 2590 -358
rect 2642 -410 2677 -358
rect 2729 -410 2764 -358
rect 2816 -410 2822 -358
rect 2410 -440 2822 -410
rect 3472 -687 3524 50
tri 3524 23 3551 50 nw
rect 3733 -664 3863 1484
rect 8246 1556 8282 1608
rect 8334 1556 8349 1608
rect 8401 1556 8418 1608
rect 8246 1530 8418 1556
rect 8246 1478 8282 1530
rect 8334 1478 8349 1530
rect 8401 1478 8418 1530
rect 9126 1562 10531 1593
rect 9126 1510 9132 1562
rect 9184 1510 9199 1562
rect 9251 1510 9267 1562
rect 9319 1510 9335 1562
rect 9387 1510 9403 1562
rect 9455 1510 9471 1562
rect 9523 1510 9539 1562
rect 9591 1510 9607 1562
rect 9659 1510 9675 1562
rect 9727 1510 10531 1562
rect 9126 1479 10531 1510
rect 6033 281 6039 333
rect 6091 317 6109 333
rect 6161 317 6179 333
rect 6231 317 6249 333
rect 6100 281 6109 317
rect 6231 281 6244 317
rect 6301 281 6319 333
rect 6371 317 6388 333
rect 6440 317 6457 333
rect 6440 281 6444 317
rect 6509 281 6515 333
rect 6033 261 6044 281
rect 6100 261 6144 281
rect 6200 261 6244 281
rect 6300 261 6344 281
rect 6400 261 6444 281
rect 6500 261 6515 281
rect 6033 177 6515 261
rect 6033 121 6044 177
rect 6100 121 6144 177
rect 6200 121 6244 177
rect 6300 121 6344 177
rect 6400 121 6444 177
rect 6500 121 6515 177
rect 6033 37 6515 121
rect 6033 21 6044 37
rect 6100 21 6144 37
rect 6200 21 6244 37
rect 6300 21 6344 37
rect 6400 21 6444 37
rect 6500 21 6515 37
rect 6033 -31 6039 21
rect 6100 -19 6123 21
rect 6200 -19 6207 21
rect 6343 -19 6344 21
rect 6426 -19 6444 21
rect 6091 -31 6123 -19
rect 6175 -31 6207 -19
rect 6259 -31 6291 -19
rect 6343 -31 6374 -19
rect 6426 -31 6457 -19
rect 6509 -31 6515 21
rect 6033 -45 6515 -31
rect 6033 -97 6039 -45
rect 6091 -97 6123 -45
rect 6175 -97 6207 -45
rect 6259 -97 6291 -45
rect 6343 -97 6374 -45
rect 6426 -97 6457 -45
rect 6509 -97 6515 -45
rect 6033 -103 6515 -97
rect 6033 -159 6044 -103
rect 6100 -159 6144 -103
rect 6200 -159 6244 -103
rect 6300 -159 6344 -103
rect 6400 -159 6444 -103
rect 6500 -159 6515 -103
rect 6033 -244 6515 -159
rect 6033 -291 6044 -244
rect 6100 -291 6144 -244
rect 6200 -291 6244 -244
rect 6300 -291 6344 -244
rect 6400 -291 6444 -244
rect 6500 -291 6515 -244
rect 6033 -343 6039 -291
rect 6100 -300 6109 -291
rect 6231 -300 6244 -291
rect 6091 -343 6109 -300
rect 6161 -343 6179 -300
rect 6231 -343 6249 -300
rect 6301 -343 6319 -291
rect 6440 -300 6444 -291
rect 6371 -343 6388 -300
rect 6440 -343 6457 -300
rect 6509 -343 6515 -291
rect 6033 -385 6515 -343
rect 6033 -407 6044 -385
rect 6100 -407 6144 -385
rect 6200 -407 6244 -385
rect 6300 -407 6344 -385
rect 6400 -407 6444 -385
rect 6500 -407 6515 -385
rect 6033 -459 6039 -407
rect 6100 -441 6109 -407
rect 6231 -441 6244 -407
rect 6091 -459 6109 -441
rect 6161 -459 6179 -441
rect 6231 -459 6249 -441
rect 6301 -459 6319 -407
rect 6440 -441 6444 -407
rect 6371 -459 6388 -441
rect 6440 -459 6457 -441
rect 6509 -459 6515 -407
rect 6658 281 6664 333
rect 6716 317 6733 333
rect 6785 317 6802 333
rect 6854 317 6872 333
rect 6924 317 6942 333
rect 6994 317 7012 333
rect 7064 317 7082 333
rect 6727 281 6733 317
rect 6854 281 6871 317
rect 6927 281 6942 317
rect 7064 281 7071 317
rect 7134 281 7140 333
rect 6658 261 6671 281
rect 6727 261 6771 281
rect 6827 261 6871 281
rect 6927 261 6971 281
rect 7027 261 7071 281
rect 7127 261 7140 281
rect 6658 177 7140 261
rect 6658 121 6671 177
rect 6727 121 6771 177
rect 6827 121 6871 177
rect 6927 121 6971 177
rect 7027 121 7071 177
rect 7127 121 7140 177
rect 6658 37 7140 121
rect 6658 21 6671 37
rect 6727 21 6771 37
rect 6827 21 6871 37
rect 6927 21 6971 37
rect 7027 21 7071 37
rect 7127 21 7140 37
rect 6658 -31 6664 21
rect 6727 -19 6748 21
rect 6827 -19 6832 21
rect 6968 -19 6971 21
rect 7051 -19 7071 21
rect 6716 -31 6748 -19
rect 6800 -31 6832 -19
rect 6884 -31 6916 -19
rect 6968 -31 6999 -19
rect 7051 -31 7082 -19
rect 7134 -31 7140 21
rect 6658 -45 7140 -31
rect 6658 -97 6664 -45
rect 6716 -97 6748 -45
rect 6800 -97 6832 -45
rect 6884 -97 6916 -45
rect 6968 -97 6999 -45
rect 7051 -97 7082 -45
rect 7134 -97 7140 -45
rect 6658 -103 7140 -97
rect 6658 -159 6671 -103
rect 6727 -159 6771 -103
rect 6827 -159 6871 -103
rect 6927 -159 6971 -103
rect 7027 -159 7071 -103
rect 7127 -159 7140 -103
rect 6658 -244 7140 -159
rect 6658 -291 6671 -244
rect 6727 -291 6771 -244
rect 6827 -291 6871 -244
rect 6927 -291 6971 -244
rect 7027 -291 7071 -244
rect 7127 -291 7140 -244
rect 6658 -343 6664 -291
rect 6727 -300 6734 -291
rect 6856 -300 6871 -291
rect 6927 -300 6944 -291
rect 7065 -300 7071 -291
rect 6716 -343 6734 -300
rect 6786 -343 6804 -300
rect 6856 -343 6874 -300
rect 6926 -343 6944 -300
rect 6996 -343 7013 -300
rect 7065 -343 7082 -300
rect 7134 -343 7140 -291
rect 6658 -385 7140 -343
rect 6658 -407 6671 -385
rect 6727 -407 6771 -385
rect 6827 -407 6871 -385
rect 6927 -407 6971 -385
rect 7027 -407 7071 -385
rect 7127 -407 7140 -385
rect 8246 -402 8418 1478
tri 9938 1221 10196 1479 ne
rect 9078 321 9306 330
rect 9134 265 9164 321
rect 9220 265 9250 321
rect 9078 255 9306 265
rect 9130 230 9166 255
rect 9218 230 9254 255
rect 9134 174 9164 230
rect 9220 174 9250 230
rect 9130 139 9166 174
rect 9218 139 9254 174
rect 9134 83 9164 139
rect 9220 83 9250 139
rect 10196 172 10531 1479
rect 10944 1556 10950 1608
rect 11002 1556 11025 1608
rect 11077 1556 11100 1608
rect 11152 1556 11175 1608
rect 11227 1556 11250 1608
rect 11302 1556 11325 1608
rect 11377 1556 11383 1608
rect 10944 1530 11383 1556
rect 10944 1478 10950 1530
rect 11002 1478 11025 1530
rect 11077 1478 11100 1530
rect 11152 1478 11175 1530
rect 11227 1478 11250 1530
rect 11302 1478 11325 1530
rect 11377 1478 11383 1530
tri 10531 172 10803 444 sw
rect 10196 146 10803 172
rect 10196 94 10326 146
tri 10326 114 10358 146 nw
tri 10405 113 10438 146 ne
rect 10197 92 10325 93
rect 10438 94 10568 146
tri 10568 114 10600 146 nw
tri 10639 112 10673 146 ne
rect 10439 92 10567 93
rect 10673 94 10803 146
rect 10674 92 10802 93
rect 10944 260 11383 1478
rect 12365 1556 12371 1608
rect 12423 1556 12441 1608
rect 12493 1556 12511 1608
rect 12563 1556 12581 1608
rect 12633 1556 12651 1608
rect 12703 1556 12709 1608
rect 12365 1530 12709 1556
rect 12365 1478 12371 1530
rect 12423 1478 12441 1530
rect 12493 1478 12511 1530
rect 12563 1478 12581 1530
rect 12633 1478 12651 1530
rect 12703 1478 12709 1530
tri 11383 260 11492 369 sw
rect 12365 284 12709 1478
tri 13135 1538 13205 1608 se
rect 13205 1601 13367 1608
rect 13205 1549 13243 1601
rect 13295 1549 13309 1601
rect 13361 1549 13367 1601
rect 13205 1538 13367 1549
rect 13135 1537 13367 1538
rect 13135 1485 13243 1537
rect 13295 1485 13309 1537
rect 13361 1485 13367 1537
rect 13135 1478 13367 1485
rect 13667 1601 13797 1608
rect 13667 1549 13673 1601
rect 13725 1549 13739 1601
rect 13791 1549 13797 1601
rect 13667 1537 13797 1549
rect 13667 1485 13673 1537
rect 13725 1485 13739 1537
rect 13791 1485 13797 1537
tri 12709 284 12858 433 sw
rect 10944 146 11551 260
rect 10944 94 11074 146
tri 11074 114 11106 146 nw
tri 11153 113 11186 146 ne
rect 10945 92 11073 93
rect 11186 94 11316 146
tri 11316 114 11348 146 nw
tri 11387 112 11421 146 ne
rect 11187 92 11315 93
rect 11421 94 11551 146
rect 11422 92 11550 93
rect 12071 151 12080 207
rect 12136 203 12223 207
rect 12136 151 12155 203
rect 12207 151 12223 203
rect 12279 151 12288 207
rect 12071 123 12288 151
rect 12071 121 12082 123
rect 12134 121 12155 123
rect 9130 58 9166 83
rect 9218 58 9254 83
rect 9078 48 9306 58
rect 9134 -8 9164 48
rect 9220 -8 9250 48
rect 9130 -15 9166 -8
rect 9218 -15 9254 -8
rect 9078 -36 9306 -15
rect 9130 -43 9166 -36
rect 9218 -43 9254 -36
rect 9134 -99 9164 -43
rect 9220 -99 9250 -43
rect 9078 -109 9306 -99
rect 9130 -135 9166 -109
rect 9218 -135 9254 -109
rect 9134 -191 9164 -135
rect 9220 -191 9250 -135
rect 9078 -227 9306 -191
rect 10673 -208 10803 92
rect 11186 -208 11316 92
rect 12071 65 12080 121
rect 12136 71 12155 121
rect 12207 121 12227 123
rect 12207 71 12223 121
rect 12136 65 12223 71
rect 12279 65 12288 123
rect 12365 170 12978 284
rect 12365 118 12495 170
tri 12495 136 12529 170 nw
tri 12573 136 12607 170 ne
rect 12366 116 12494 117
rect 12607 118 12737 170
tri 12737 136 12771 170 nw
tri 12814 136 12848 170 ne
rect 12608 116 12736 117
rect 12848 118 12978 170
rect 12849 116 12977 117
rect 12003 -146 12009 -94
rect 12061 -146 12073 -94
rect 12125 -146 12131 -94
tri 12003 -184 12041 -146 ne
rect 9134 -283 9164 -227
rect 9220 -283 9250 -227
rect 9078 -292 9306 -283
rect 10197 -209 10325 -208
rect 6658 -459 6664 -407
rect 6727 -441 6734 -407
rect 6856 -441 6871 -407
rect 6927 -441 6944 -407
rect 7065 -441 7071 -407
rect 6716 -459 6734 -441
rect 6786 -459 6804 -441
rect 6856 -459 6874 -441
rect 6926 -459 6944 -441
rect 6996 -459 7013 -441
rect 7065 -459 7082 -441
rect 7134 -459 7140 -407
tri 7402 -476 7476 -402 se
rect 7476 -454 7761 -402
rect 7813 -454 7825 -402
rect 7877 -454 7883 -402
rect 8246 -454 8252 -402
rect 8304 -454 8360 -402
rect 8412 -454 8418 -402
tri 7476 -476 7498 -454 nw
tri 7382 -496 7402 -476 se
rect 7402 -496 7404 -476
tri 4525 -570 4599 -496 se
rect 4599 -548 7404 -496
tri 7404 -548 7476 -476 nw
rect 10196 -482 10326 -210
rect 10439 -209 10567 -208
rect 10438 -402 10568 -210
rect 10674 -209 10802 -208
rect 10673 -317 10803 -210
rect 10673 -369 10681 -317
rect 10733 -369 10745 -317
rect 10797 -369 10803 -317
rect 10945 -209 11073 -208
rect 10438 -454 10446 -402
rect 10498 -454 10510 -402
rect 10562 -454 10568 -402
tri 4599 -570 4621 -548 nw
tri 7479 -556 7553 -482 se
rect 7553 -534 7761 -482
rect 7813 -534 7825 -482
rect 7877 -534 7883 -482
rect 10196 -534 10204 -482
rect 10256 -534 10268 -482
rect 10320 -534 10326 -482
rect 10944 -482 11074 -210
rect 11187 -209 11315 -208
rect 11186 -402 11316 -210
rect 11422 -209 11550 -208
rect 11421 -317 11551 -210
rect 11421 -369 11429 -317
rect 11481 -369 11493 -317
rect 11545 -369 11551 -317
rect 11186 -454 11194 -402
rect 11246 -454 11258 -402
rect 11310 -454 11316 -402
rect 10944 -534 10952 -482
rect 11004 -534 11016 -482
rect 11068 -534 11074 -482
tri 12000 -482 12041 -441 se
rect 12041 -482 12093 -146
tri 12093 -184 12131 -146 nw
rect 12365 -184 12495 116
rect 12366 -185 12494 -184
tri 12093 -482 12128 -447 sw
rect 12000 -534 12006 -482
rect 12058 -534 12070 -482
rect 12122 -534 12128 -482
rect 12365 -482 12495 -186
rect 12608 -185 12736 -184
rect 12607 -402 12737 -186
rect 12849 -185 12977 -184
rect 12848 -317 12978 -186
rect 12848 -369 12856 -317
rect 12908 -369 12920 -317
rect 12972 -369 12978 -317
rect 13135 -317 13265 1478
tri 13265 1408 13335 1478 nw
tri 13592 1147 13667 1222 se
rect 13667 1147 13797 1485
rect 14229 1601 14359 1608
rect 14229 1549 14235 1601
rect 14287 1549 14301 1601
rect 14353 1549 14359 1601
rect 14229 1537 14359 1549
rect 14229 1485 14235 1537
rect 14287 1485 14301 1537
rect 14353 1485 14359 1537
rect 14229 1357 14359 1485
tri 14229 1300 14286 1357 ne
rect 14286 1328 14359 1357
tri 14359 1328 14442 1411 sw
rect 13592 1126 13797 1147
tri 13797 1126 13893 1222 sw
rect 14286 1126 14442 1328
tri 14442 1126 14563 1247 sw
rect 13592 1012 14204 1126
rect 13592 960 13722 1012
tri 13722 978 13756 1012 nw
tri 13803 978 13837 1012 ne
rect 13593 958 13721 959
rect 13837 960 13967 1012
tri 13967 978 14001 1012 nw
tri 14040 978 14074 1012 ne
rect 13838 958 13966 959
rect 14074 960 14204 1012
rect 14075 958 14203 959
rect 14286 1012 14898 1126
rect 14286 960 14416 1012
tri 14416 978 14450 1012 nw
tri 14497 978 14531 1012 ne
rect 14287 958 14415 959
rect 14531 960 14661 1012
tri 14661 978 14695 1012 nw
tri 14734 978 14768 1012 ne
rect 14532 958 14660 959
rect 14768 960 14898 1012
rect 14769 958 14897 959
rect 13837 658 13967 958
rect 14286 658 14416 958
rect 13135 -369 13141 -317
rect 13193 -369 13207 -317
rect 13259 -369 13265 -317
rect 13593 657 13721 658
rect 12607 -454 12615 -402
rect 12667 -454 12679 -402
rect 12731 -454 12737 -402
rect 12365 -534 12373 -482
rect 12425 -534 12437 -482
rect 12489 -534 12495 -482
rect 13592 -482 13722 656
rect 13838 657 13966 658
rect 13837 -402 13967 656
rect 14075 657 14203 658
rect 14074 -317 14204 656
rect 14074 -369 14082 -317
rect 14134 -369 14146 -317
rect 14198 -369 14204 -317
rect 14287 657 14415 658
rect 13837 -454 13845 -402
rect 13897 -454 13909 -402
rect 13961 -454 13967 -402
rect 13592 -534 13600 -482
rect 13652 -534 13664 -482
rect 13716 -534 13722 -482
rect 14286 -482 14416 656
rect 14532 657 14660 658
rect 14531 -402 14661 656
rect 14769 657 14897 658
tri 14712 -290 14768 -234 se
rect 14768 -290 14898 656
tri 14898 -290 14972 -216 sw
rect 14712 -342 14737 -290
rect 14789 -342 14801 -290
rect 14853 -342 14865 -290
rect 14917 -342 14929 -290
rect 14981 -342 14993 -290
rect 15045 -342 15057 -290
rect 15109 -342 15115 -290
rect 14531 -454 14539 -402
rect 14591 -454 14603 -402
rect 14655 -454 14661 -402
rect 15035 -427 15041 -375
rect 15093 -427 15106 -375
rect 15158 -427 15164 -375
rect 14286 -534 14294 -482
rect 14346 -534 14358 -482
rect 14410 -534 14416 -482
rect 15042 -461 15094 -455
rect 15042 -525 15094 -513
tri 7553 -556 7575 -534 nw
tri 3472 -739 3524 -687 ne
tri 3524 -724 3583 -665 sw
rect 3524 -739 3583 -724
tri 3524 -776 3561 -739 ne
rect 3561 -776 3583 -739
tri 3583 -776 3635 -724 sw
tri 3561 -850 3635 -776 ne
tri 3635 -850 3709 -776 sw
tri 3733 -790 3859 -664 ne
rect 3859 -738 3863 -664
tri 3863 -738 3970 -631 sw
tri 4451 -644 4525 -570 se
tri 4525 -644 4599 -570 nw
tri 7459 -576 7479 -556 se
rect 7479 -576 7481 -556
tri 4377 -718 4451 -644 se
tri 4451 -718 4525 -644 nw
tri 4602 -650 4676 -576 se
rect 4676 -628 7481 -576
tri 7481 -628 7553 -556 nw
rect 14880 -614 14886 -562
rect 14938 -614 14950 -562
rect 15002 -614 15008 -562
rect 15042 -583 15094 -577
tri 4676 -650 4698 -628 nw
tri 4357 -738 4377 -718 se
rect 4377 -738 4379 -718
rect 3859 -790 4379 -738
tri 4379 -790 4451 -718 nw
tri 4528 -724 4602 -650 se
tri 4602 -724 4676 -650 nw
rect 14800 -695 14806 -643
rect 14858 -695 14870 -643
rect 14922 -695 14928 -643
tri 4454 -798 4528 -724 se
tri 4528 -798 4602 -724 nw
tri 4402 -850 4454 -798 se
rect 4454 -850 4476 -798
tri 4476 -850 4528 -798 nw
tri 3635 -902 3687 -850 ne
rect 3687 -902 4424 -850
tri 4424 -902 4476 -850 nw
<< rmetal2 >>
rect 10196 93 10326 94
rect 10196 92 10197 93
rect 10325 92 10326 93
rect 10438 93 10568 94
rect 10438 92 10439 93
rect 10567 92 10568 93
rect 10673 93 10803 94
rect 10673 92 10674 93
rect 10802 92 10803 93
rect 10944 93 11074 94
rect 10944 92 10945 93
rect 11073 92 11074 93
rect 11186 93 11316 94
rect 11186 92 11187 93
rect 11315 92 11316 93
rect 11421 93 11551 94
rect 11421 92 11422 93
rect 11550 92 11551 93
rect 12365 117 12495 118
rect 12365 116 12366 117
rect 12494 116 12495 117
rect 12607 117 12737 118
rect 12607 116 12608 117
rect 12736 116 12737 117
rect 12848 117 12978 118
rect 12848 116 12849 117
rect 12977 116 12978 117
rect 10196 -209 10197 -208
rect 10325 -209 10326 -208
rect 10196 -210 10326 -209
rect 10438 -209 10439 -208
rect 10567 -209 10568 -208
rect 10438 -210 10568 -209
rect 10673 -209 10674 -208
rect 10802 -209 10803 -208
rect 10673 -210 10803 -209
rect 10944 -209 10945 -208
rect 11073 -209 11074 -208
rect 10944 -210 11074 -209
rect 11186 -209 11187 -208
rect 11315 -209 11316 -208
rect 11186 -210 11316 -209
rect 11421 -209 11422 -208
rect 11550 -209 11551 -208
rect 11421 -210 11551 -209
rect 12365 -185 12366 -184
rect 12494 -185 12495 -184
rect 12365 -186 12495 -185
rect 12607 -185 12608 -184
rect 12736 -185 12737 -184
rect 12607 -186 12737 -185
rect 12848 -185 12849 -184
rect 12977 -185 12978 -184
rect 12848 -186 12978 -185
rect 13592 959 13722 960
rect 13592 958 13593 959
rect 13721 958 13722 959
rect 13837 959 13967 960
rect 13837 958 13838 959
rect 13966 958 13967 959
rect 14074 959 14204 960
rect 14074 958 14075 959
rect 14203 958 14204 959
rect 14286 959 14416 960
rect 14286 958 14287 959
rect 14415 958 14416 959
rect 14531 959 14661 960
rect 14531 958 14532 959
rect 14660 958 14661 959
rect 14768 959 14898 960
rect 14768 958 14769 959
rect 14897 958 14898 959
rect 13592 657 13593 658
rect 13721 657 13722 658
rect 13592 656 13722 657
rect 13837 657 13838 658
rect 13966 657 13967 658
rect 13837 656 13967 657
rect 14074 657 14075 658
rect 14203 657 14204 658
rect 14074 656 14204 657
rect 14286 657 14287 658
rect 14415 657 14416 658
rect 14286 656 14416 657
rect 14531 657 14532 658
rect 14660 657 14661 658
rect 14531 656 14661 657
rect 14768 657 14769 658
rect 14897 657 14898 658
rect 14768 656 14898 657
<< via2 >>
rect 6044 281 6091 317
rect 6091 281 6100 317
rect 6144 281 6161 317
rect 6161 281 6179 317
rect 6179 281 6200 317
rect 6244 281 6249 317
rect 6249 281 6300 317
rect 6344 281 6371 317
rect 6371 281 6388 317
rect 6388 281 6400 317
rect 6444 281 6457 317
rect 6457 281 6500 317
rect 6044 261 6100 281
rect 6144 261 6200 281
rect 6244 261 6300 281
rect 6344 261 6400 281
rect 6444 261 6500 281
rect 6044 121 6100 177
rect 6144 121 6200 177
rect 6244 121 6300 177
rect 6344 121 6400 177
rect 6444 121 6500 177
rect 6044 21 6100 37
rect 6144 21 6200 37
rect 6244 21 6300 37
rect 6344 21 6400 37
rect 6444 21 6500 37
rect 6044 -19 6091 21
rect 6091 -19 6100 21
rect 6144 -19 6175 21
rect 6175 -19 6200 21
rect 6244 -19 6259 21
rect 6259 -19 6291 21
rect 6291 -19 6300 21
rect 6344 -19 6374 21
rect 6374 -19 6400 21
rect 6444 -19 6457 21
rect 6457 -19 6500 21
rect 6044 -159 6100 -103
rect 6144 -159 6200 -103
rect 6244 -159 6300 -103
rect 6344 -159 6400 -103
rect 6444 -159 6500 -103
rect 6044 -291 6100 -244
rect 6144 -291 6200 -244
rect 6244 -291 6300 -244
rect 6344 -291 6400 -244
rect 6444 -291 6500 -244
rect 6044 -300 6091 -291
rect 6091 -300 6100 -291
rect 6144 -300 6161 -291
rect 6161 -300 6179 -291
rect 6179 -300 6200 -291
rect 6244 -300 6249 -291
rect 6249 -300 6300 -291
rect 6344 -300 6371 -291
rect 6371 -300 6388 -291
rect 6388 -300 6400 -291
rect 6444 -300 6457 -291
rect 6457 -300 6500 -291
rect 6044 -407 6100 -385
rect 6144 -407 6200 -385
rect 6244 -407 6300 -385
rect 6344 -407 6400 -385
rect 6444 -407 6500 -385
rect 6044 -441 6091 -407
rect 6091 -441 6100 -407
rect 6144 -441 6161 -407
rect 6161 -441 6179 -407
rect 6179 -441 6200 -407
rect 6244 -441 6249 -407
rect 6249 -441 6300 -407
rect 6344 -441 6371 -407
rect 6371 -441 6388 -407
rect 6388 -441 6400 -407
rect 6444 -441 6457 -407
rect 6457 -441 6500 -407
rect 6671 281 6716 317
rect 6716 281 6727 317
rect 6771 281 6785 317
rect 6785 281 6802 317
rect 6802 281 6827 317
rect 6871 281 6872 317
rect 6872 281 6924 317
rect 6924 281 6927 317
rect 6971 281 6994 317
rect 6994 281 7012 317
rect 7012 281 7027 317
rect 7071 281 7082 317
rect 7082 281 7127 317
rect 6671 261 6727 281
rect 6771 261 6827 281
rect 6871 261 6927 281
rect 6971 261 7027 281
rect 7071 261 7127 281
rect 6671 121 6727 177
rect 6771 121 6827 177
rect 6871 121 6927 177
rect 6971 121 7027 177
rect 7071 121 7127 177
rect 6671 21 6727 37
rect 6771 21 6827 37
rect 6871 21 6927 37
rect 6971 21 7027 37
rect 7071 21 7127 37
rect 6671 -19 6716 21
rect 6716 -19 6727 21
rect 6771 -19 6800 21
rect 6800 -19 6827 21
rect 6871 -19 6884 21
rect 6884 -19 6916 21
rect 6916 -19 6927 21
rect 6971 -19 6999 21
rect 6999 -19 7027 21
rect 7071 -19 7082 21
rect 7082 -19 7127 21
rect 6671 -159 6727 -103
rect 6771 -159 6827 -103
rect 6871 -159 6927 -103
rect 6971 -159 7027 -103
rect 7071 -159 7127 -103
rect 6671 -291 6727 -244
rect 6771 -291 6827 -244
rect 6871 -291 6927 -244
rect 6971 -291 7027 -244
rect 7071 -291 7127 -244
rect 6671 -300 6716 -291
rect 6716 -300 6727 -291
rect 6771 -300 6786 -291
rect 6786 -300 6804 -291
rect 6804 -300 6827 -291
rect 6871 -300 6874 -291
rect 6874 -300 6926 -291
rect 6926 -300 6927 -291
rect 6971 -300 6996 -291
rect 6996 -300 7013 -291
rect 7013 -300 7027 -291
rect 7071 -300 7082 -291
rect 7082 -300 7127 -291
rect 6671 -407 6727 -385
rect 6771 -407 6827 -385
rect 6871 -407 6927 -385
rect 6971 -407 7027 -385
rect 7071 -407 7127 -385
rect 9078 265 9134 321
rect 9164 265 9220 321
rect 9250 265 9306 321
rect 9078 203 9130 230
rect 9130 203 9134 230
rect 9078 183 9134 203
rect 9078 174 9130 183
rect 9130 174 9134 183
rect 9164 203 9166 230
rect 9166 203 9218 230
rect 9218 203 9220 230
rect 9164 183 9220 203
rect 9164 174 9166 183
rect 9166 174 9218 183
rect 9218 174 9220 183
rect 9250 203 9254 230
rect 9254 203 9306 230
rect 9250 183 9306 203
rect 9250 174 9254 183
rect 9254 174 9306 183
rect 9078 131 9130 139
rect 9130 131 9134 139
rect 9078 110 9134 131
rect 9078 83 9130 110
rect 9130 83 9134 110
rect 9164 131 9166 139
rect 9166 131 9218 139
rect 9218 131 9220 139
rect 9164 110 9220 131
rect 9164 83 9166 110
rect 9166 83 9218 110
rect 9218 83 9220 110
rect 9250 131 9254 139
rect 9254 131 9306 139
rect 9250 110 9306 131
rect 9250 83 9254 110
rect 9254 83 9306 110
rect 12080 203 12136 207
rect 12223 203 12279 207
rect 12080 151 12082 203
rect 12082 151 12134 203
rect 12134 151 12136 203
rect 12223 151 12227 203
rect 12227 151 12279 203
rect 9078 37 9134 48
rect 9078 -8 9130 37
rect 9130 -8 9134 37
rect 9164 37 9220 48
rect 9164 -8 9166 37
rect 9166 -8 9218 37
rect 9218 -8 9220 37
rect 9250 37 9306 48
rect 9250 -8 9254 37
rect 9254 -8 9306 37
rect 9078 -88 9130 -43
rect 9130 -88 9134 -43
rect 9078 -99 9134 -88
rect 9164 -88 9166 -43
rect 9166 -88 9218 -43
rect 9218 -88 9220 -43
rect 9164 -99 9220 -88
rect 9250 -88 9254 -43
rect 9254 -88 9306 -43
rect 9250 -99 9306 -88
rect 9078 -161 9130 -135
rect 9130 -161 9134 -135
rect 9078 -191 9134 -161
rect 9164 -161 9166 -135
rect 9166 -161 9218 -135
rect 9218 -161 9220 -135
rect 9164 -191 9220 -161
rect 9250 -161 9254 -135
rect 9254 -161 9306 -135
rect 9250 -191 9306 -161
rect 12080 71 12082 121
rect 12082 71 12134 121
rect 12134 71 12136 121
rect 12223 71 12227 121
rect 12227 71 12279 121
rect 12080 65 12136 71
rect 12223 65 12279 71
rect 9078 -283 9134 -227
rect 9164 -283 9220 -227
rect 9250 -283 9306 -227
rect 6671 -441 6716 -407
rect 6716 -441 6727 -407
rect 6771 -441 6786 -407
rect 6786 -441 6804 -407
rect 6804 -441 6827 -407
rect 6871 -441 6874 -407
rect 6874 -441 6926 -407
rect 6926 -441 6927 -407
rect 6971 -441 6996 -407
rect 6996 -441 7013 -407
rect 7013 -441 7027 -407
rect 7071 -441 7082 -407
rect 7082 -441 7127 -407
<< metal3 >>
rect 9073 326 9311 332
rect 6036 317 6508 322
rect 6036 261 6044 317
rect 6100 261 6144 317
rect 6200 261 6244 317
rect 6300 261 6344 317
rect 6400 261 6444 317
rect 6500 261 6508 317
rect 6036 177 6508 261
rect 6036 121 6044 177
rect 6100 121 6144 177
rect 6200 121 6244 177
rect 6300 121 6344 177
rect 6400 121 6444 177
rect 6500 121 6508 177
rect 6036 37 6508 121
rect 6036 -19 6044 37
rect 6100 -19 6144 37
rect 6200 -19 6244 37
rect 6300 -19 6344 37
rect 6400 -19 6444 37
rect 6500 -19 6508 37
rect 6036 -103 6508 -19
rect 6036 -159 6044 -103
rect 6100 -159 6144 -103
rect 6200 -159 6244 -103
rect 6300 -159 6344 -103
rect 6400 -159 6444 -103
rect 6500 -159 6508 -103
rect 6036 -244 6508 -159
rect 6036 -300 6044 -244
rect 6100 -300 6144 -244
rect 6200 -300 6244 -244
rect 6300 -300 6344 -244
rect 6400 -300 6444 -244
rect 6500 -300 6508 -244
rect 6036 -385 6508 -300
rect 6036 -441 6044 -385
rect 6100 -441 6144 -385
rect 6200 -441 6244 -385
rect 6300 -441 6344 -385
rect 6400 -441 6444 -385
rect 6500 -441 6508 -385
rect 6036 -446 6508 -441
rect 6663 317 7135 322
rect 6663 261 6671 317
rect 6727 261 6771 317
rect 6827 261 6871 317
rect 6927 261 6971 317
rect 7027 261 7071 317
rect 7127 261 7135 317
rect 6663 177 7135 261
rect 6663 121 6671 177
rect 6727 121 6771 177
rect 6827 121 6871 177
rect 6927 121 6971 177
rect 7027 121 7071 177
rect 7127 121 7135 177
rect 6663 37 7135 121
rect 6663 -19 6671 37
rect 6727 -19 6771 37
rect 6827 -19 6871 37
rect 6927 -19 6971 37
rect 7027 -19 7071 37
rect 7127 -19 7135 37
rect 6663 -103 7135 -19
rect 6663 -159 6671 -103
rect 6727 -159 6771 -103
rect 6827 -159 6871 -103
rect 6927 -159 6971 -103
rect 7027 -159 7071 -103
rect 7127 -159 7135 -103
rect 6663 -244 7135 -159
rect 6663 -300 6671 -244
rect 6727 -300 6771 -244
rect 6827 -300 6871 -244
rect 6927 -300 6971 -244
rect 7027 -300 7071 -244
rect 7127 -300 7135 -244
rect 9073 262 9074 326
rect 9138 262 9160 326
rect 9224 262 9246 326
rect 9310 262 9311 326
rect 9073 235 9311 262
rect 9073 171 9074 235
rect 9138 171 9160 235
rect 9224 171 9246 235
rect 9310 171 9311 235
rect 9073 143 9311 171
rect 9073 79 9074 143
rect 9138 79 9160 143
rect 9224 79 9246 143
rect 9310 79 9311 143
rect 9073 51 9311 79
rect 12075 207 12284 212
rect 12075 151 12080 207
rect 12136 151 12223 207
rect 12279 151 12284 207
rect 12075 121 12284 151
rect 12075 65 12080 121
rect 12136 65 12223 121
rect 12279 65 12284 121
rect 12075 60 12284 65
rect 9073 -13 9074 51
rect 9138 -13 9160 51
rect 9224 -13 9246 51
rect 9310 -13 9311 51
rect 9073 -41 9311 -13
rect 9073 -105 9074 -41
rect 9138 -105 9160 -41
rect 9224 -105 9246 -41
rect 9310 -105 9311 -41
rect 9073 -133 9311 -105
rect 9073 -197 9074 -133
rect 9138 -197 9160 -133
rect 9224 -197 9246 -133
rect 9310 -197 9311 -133
rect 9073 -227 9311 -197
rect 9073 -283 9078 -227
rect 9134 -283 9164 -227
rect 9220 -283 9250 -227
rect 9306 -283 9311 -227
rect 9073 -288 9311 -283
rect 6663 -385 7135 -300
rect 6663 -441 6671 -385
rect 6727 -441 6771 -385
rect 6827 -441 6871 -385
rect 6927 -441 6971 -385
rect 7027 -441 7071 -385
rect 7127 -441 7135 -385
rect 6663 -446 7135 -441
<< via3 >>
rect 9074 321 9138 326
rect 9074 265 9078 321
rect 9078 265 9134 321
rect 9134 265 9138 321
rect 9074 262 9138 265
rect 9160 321 9224 326
rect 9160 265 9164 321
rect 9164 265 9220 321
rect 9220 265 9224 321
rect 9160 262 9224 265
rect 9246 321 9310 326
rect 9246 265 9250 321
rect 9250 265 9306 321
rect 9306 265 9310 321
rect 9246 262 9310 265
rect 9074 230 9138 235
rect 9074 174 9078 230
rect 9078 174 9134 230
rect 9134 174 9138 230
rect 9074 171 9138 174
rect 9160 230 9224 235
rect 9160 174 9164 230
rect 9164 174 9220 230
rect 9220 174 9224 230
rect 9160 171 9224 174
rect 9246 230 9310 235
rect 9246 174 9250 230
rect 9250 174 9306 230
rect 9306 174 9310 230
rect 9246 171 9310 174
rect 9074 139 9138 143
rect 9074 83 9078 139
rect 9078 83 9134 139
rect 9134 83 9138 139
rect 9074 79 9138 83
rect 9160 139 9224 143
rect 9160 83 9164 139
rect 9164 83 9220 139
rect 9220 83 9224 139
rect 9160 79 9224 83
rect 9246 139 9310 143
rect 9246 83 9250 139
rect 9250 83 9306 139
rect 9306 83 9310 139
rect 9246 79 9310 83
rect 9074 48 9138 51
rect 9074 -8 9078 48
rect 9078 -8 9134 48
rect 9134 -8 9138 48
rect 9074 -13 9138 -8
rect 9160 48 9224 51
rect 9160 -8 9164 48
rect 9164 -8 9220 48
rect 9220 -8 9224 48
rect 9160 -13 9224 -8
rect 9246 48 9310 51
rect 9246 -8 9250 48
rect 9250 -8 9306 48
rect 9306 -8 9310 48
rect 9246 -13 9310 -8
rect 9074 -43 9138 -41
rect 9074 -99 9078 -43
rect 9078 -99 9134 -43
rect 9134 -99 9138 -43
rect 9074 -105 9138 -99
rect 9160 -43 9224 -41
rect 9160 -99 9164 -43
rect 9164 -99 9220 -43
rect 9220 -99 9224 -43
rect 9160 -105 9224 -99
rect 9246 -43 9310 -41
rect 9246 -99 9250 -43
rect 9250 -99 9306 -43
rect 9306 -99 9310 -43
rect 9246 -105 9310 -99
rect 9074 -135 9138 -133
rect 9074 -191 9078 -135
rect 9078 -191 9134 -135
rect 9134 -191 9138 -135
rect 9074 -197 9138 -191
rect 9160 -135 9224 -133
rect 9160 -191 9164 -135
rect 9164 -191 9220 -135
rect 9220 -191 9224 -135
rect 9160 -197 9224 -191
rect 9246 -135 9310 -133
rect 9246 -191 9250 -135
rect 9250 -191 9306 -135
rect 9306 -191 9310 -135
rect 9246 -197 9310 -191
<< metal4 >>
rect 9072 326 9312 327
rect 9072 262 9074 326
rect 9138 262 9160 326
rect 9224 262 9246 326
rect 9310 262 9312 326
rect 9072 235 9312 262
rect 9072 171 9074 235
rect 9138 171 9160 235
rect 9224 171 9246 235
rect 9310 171 9312 235
rect 9072 143 9312 171
rect 9072 79 9074 143
rect 9138 79 9160 143
rect 9224 79 9246 143
rect 9310 79 9312 143
rect 9072 51 9312 79
rect 9072 -13 9074 51
rect 9138 -13 9160 51
rect 9224 -13 9246 51
rect 9310 -13 9312 51
rect 9072 -41 9312 -13
rect 9072 -105 9074 -41
rect 9138 -105 9160 -41
rect 9224 -105 9246 -41
rect 9310 -105 9312 -41
rect 9072 -133 9312 -105
rect 9072 -197 9074 -133
rect 9138 -197 9160 -133
rect 9224 -197 9246 -133
rect 9310 -197 9312 -133
rect 9072 -198 9312 -197
use sky130_fd_io__pfet_con_diff_wo_abt_270v2  sky130_fd_io__pfet_con_diff_wo_abt_270v2_0
timestamp 1676037725
transform 1 0 457 0 1 346
box 10 288 15126 5118
use sky130_fd_io__tk_em2o_cdns_55959141808653  sky130_fd_io__tk_em2o_cdns_55959141808653_0
timestamp 1676037725
transform 0 1 14074 1 0 604
box 0 0 1 1
use sky130_fd_io__tk_em2o_cdns_55959141808653  sky130_fd_io__tk_em2o_cdns_55959141808653_1
timestamp 1676037725
transform 0 1 14531 1 0 604
box 0 0 1 1
use sky130_fd_io__tk_em2o_cdns_55959141808653  sky130_fd_io__tk_em2o_cdns_55959141808653_2
timestamp 1676037725
transform 0 1 13592 1 0 604
box 0 0 1 1
use sky130_fd_io__tk_em2o_cdns_55959141808653  sky130_fd_io__tk_em2o_cdns_55959141808653_3
timestamp 1676037725
transform 0 1 10196 1 0 -262
box 0 0 1 1
use sky130_fd_io__tk_em2o_cdns_55959141808653  sky130_fd_io__tk_em2o_cdns_55959141808653_4
timestamp 1676037725
transform 0 1 10438 1 0 -262
box 0 0 1 1
use sky130_fd_io__tk_em2o_cdns_55959141808653  sky130_fd_io__tk_em2o_cdns_55959141808653_5
timestamp 1676037725
transform 0 1 11421 1 0 -262
box 0 0 1 1
use sky130_fd_io__tk_em2o_cdns_55959141808653  sky130_fd_io__tk_em2o_cdns_55959141808653_6
timestamp 1676037725
transform 0 1 10944 1 0 -262
box 0 0 1 1
use sky130_fd_io__tk_em2o_cdns_55959141808653  sky130_fd_io__tk_em2o_cdns_55959141808653_7
timestamp 1676037725
transform 0 1 12848 1 0 -238
box 0 0 1 1
use sky130_fd_io__tk_em2o_cdns_55959141808653  sky130_fd_io__tk_em2o_cdns_55959141808653_8
timestamp 1676037725
transform 0 1 14768 1 0 604
box 0 0 1 1
use sky130_fd_io__tk_em2o_cdns_55959141808653  sky130_fd_io__tk_em2o_cdns_55959141808653_9
timestamp 1676037725
transform 0 1 12607 1 0 -238
box 0 0 1 1
use sky130_fd_io__tk_em2s_cdns_55959141808652  sky130_fd_io__tk_em2s_cdns_55959141808652_0
timestamp 1676037725
transform 0 1 14286 1 0 604
box 0 0 1 1
use sky130_fd_io__tk_em2s_cdns_55959141808652  sky130_fd_io__tk_em2s_cdns_55959141808652_1
timestamp 1676037725
transform 0 1 13837 1 0 604
box 0 0 1 1
use sky130_fd_io__tk_em2s_cdns_55959141808652  sky130_fd_io__tk_em2s_cdns_55959141808652_2
timestamp 1676037725
transform 0 1 10673 1 0 -262
box 0 0 1 1
use sky130_fd_io__tk_em2s_cdns_55959141808652  sky130_fd_io__tk_em2s_cdns_55959141808652_3
timestamp 1676037725
transform 0 1 11186 1 0 -262
box 0 0 1 1
use sky130_fd_io__tk_em2s_cdns_55959141808652  sky130_fd_io__tk_em2s_cdns_55959141808652_4
timestamp 1676037725
transform 0 1 12365 1 0 -238
box 0 0 1 1
use sky130_fd_pr__res_generic_po__example_5595914180838  sky130_fd_pr__res_generic_po__example_5595914180838_0
timestamp 1676037725
transform 1 0 12535 0 1 -157
box 15 17 2025 18
use sky130_fd_pr__via_pol1_centered__example_559591418081  sky130_fd_pr__via_pol1_centered__example_559591418081_0
timestamp 1676037725
transform -1 0 14660 0 -1 -107
box 0 0 1 1
use sky130_fd_pr__via_pol1_centered__example_559591418081  sky130_fd_pr__via_pol1_centered__example_559591418081_1
timestamp 1676037725
transform 1 0 12450 0 -1 -107
box 0 0 1 1
<< labels >>
flabel comment s 13504 -98 13504 -98 0 FreeSans 440 0 0 0 LEAKER
flabel metal1 s 10483 -454 10635 -402 0 FreeSans 400 180 0 0 PU_H_N[3]
port 2 nsew
flabel metal1 s 10299 -369 10384 -317 0 FreeSans 400 180 0 0 PU_H_N[2]
port 3 nsew
flabel metal1 s 2636 391 2636 391 0 FreeSans 400 0 0 0 VCC_IO
flabel metal1 s 9905 -508 9905 -508 0 FreeSans 400 180 0 0 TIE_HI_ESD
flabel metal1 s 12712 661 12811 745 3 FreeSans 520 0 0 0 VNB
port 4 nsew
flabel metal2 s 13565 1988 14578 2981 0 FreeSans 400 180 0 0 VCC_IO
port 5 nsew
flabel metal2 s 11366 3389 13325 4498 3 FreeSans 520 0 0 0 PAD
port 6 nsew
<< properties >>
string GDS_END 47383350
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 47342654
<< end >>
