* NGSPICE file created from sky130_fd_pr__rf_npn_11v0_W1p00L1p00.ext - technology: sky130A

.subckt sky130_fd_pr__rf_npn_11v0_W1p00L1p00 E B C
X0 C B a_425_425# VSUBS sky130_fd_pr__npn_11v0 area=8.01025e+13p
.ends

