magic
tech sky130A
magscale 1 2
timestamp 1676037725
<< nwell >>
rect -38 261 682 582
<< pwell >>
rect 416 157 643 203
rect 1 21 643 157
rect 29 -17 63 21
<< scnmos >>
rect 79 47 109 131
rect 167 47 197 131
rect 273 47 303 131
rect 369 47 399 131
rect 535 47 565 177
<< scpmoshvt >>
rect 79 413 109 497
rect 179 413 209 497
rect 283 413 313 497
rect 369 413 399 497
rect 535 297 565 497
<< ndiff >>
rect 442 161 535 177
rect 442 131 476 161
rect 27 101 79 131
rect 27 67 35 101
rect 69 67 79 101
rect 27 47 79 67
rect 109 47 167 131
rect 197 47 273 131
rect 303 47 369 131
rect 399 127 476 131
rect 510 127 535 161
rect 399 93 535 127
rect 399 59 476 93
rect 510 59 535 93
rect 399 47 535 59
rect 565 161 617 177
rect 565 127 575 161
rect 609 127 617 161
rect 565 93 617 127
rect 565 59 575 93
rect 609 59 617 93
rect 565 47 617 59
<< pdiff >>
rect 27 485 79 497
rect 27 451 35 485
rect 69 451 79 485
rect 27 413 79 451
rect 109 477 179 497
rect 109 443 127 477
rect 161 443 179 477
rect 109 413 179 443
rect 209 485 283 497
rect 209 451 229 485
rect 263 451 283 485
rect 209 413 283 451
rect 313 477 369 497
rect 313 443 324 477
rect 358 443 369 477
rect 313 413 369 443
rect 399 485 535 497
rect 399 451 475 485
rect 509 451 535 485
rect 399 417 535 451
rect 399 413 475 417
rect 418 383 475 413
rect 509 383 535 417
rect 418 297 535 383
rect 565 485 617 497
rect 565 451 575 485
rect 609 451 617 485
rect 565 417 617 451
rect 565 383 575 417
rect 609 383 617 417
rect 565 349 617 383
rect 565 315 575 349
rect 609 315 617 349
rect 565 297 617 315
<< ndiffc >>
rect 35 67 69 101
rect 476 127 510 161
rect 476 59 510 93
rect 575 127 609 161
rect 575 59 609 93
<< pdiffc >>
rect 35 451 69 485
rect 127 443 161 477
rect 229 451 263 485
rect 324 443 358 477
rect 475 451 509 485
rect 475 383 509 417
rect 575 451 609 485
rect 575 383 609 417
rect 575 315 609 349
<< poly >>
rect 79 497 109 523
rect 179 497 209 523
rect 283 497 313 523
rect 369 497 399 523
rect 535 497 565 523
rect 79 265 109 413
rect 179 265 209 413
rect 283 265 313 413
rect 369 265 399 413
rect 535 265 565 297
rect 21 249 109 265
rect 21 215 31 249
rect 65 215 109 249
rect 21 199 109 215
rect 79 131 109 199
rect 167 249 221 265
rect 167 215 177 249
rect 211 215 221 249
rect 167 199 221 215
rect 273 249 327 265
rect 273 215 283 249
rect 317 215 327 249
rect 273 199 327 215
rect 369 249 433 265
rect 369 215 379 249
rect 413 215 433 249
rect 369 199 433 215
rect 480 249 565 265
rect 480 215 490 249
rect 524 215 565 249
rect 480 199 565 215
rect 167 131 197 199
rect 273 131 303 199
rect 369 131 399 199
rect 535 177 565 199
rect 79 21 109 47
rect 167 21 197 47
rect 273 21 303 47
rect 369 21 399 47
rect 535 21 565 47
<< polycont >>
rect 31 215 65 249
rect 177 215 211 249
rect 283 215 317 249
rect 379 215 413 249
rect 490 215 524 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 18 485 85 527
rect 18 451 35 485
rect 69 451 85 485
rect 119 477 169 493
rect 119 443 127 477
rect 161 443 169 477
rect 17 249 65 415
rect 119 333 169 443
rect 213 485 279 527
rect 213 451 229 485
rect 263 451 279 485
rect 213 383 279 451
rect 316 477 366 493
rect 316 443 324 477
rect 358 443 366 477
rect 316 333 366 443
rect 459 485 525 527
rect 459 451 475 485
rect 509 451 525 485
rect 459 417 525 451
rect 559 485 627 493
rect 559 451 575 485
rect 609 451 627 485
rect 559 441 627 451
rect 459 383 475 417
rect 509 383 525 417
rect 459 367 525 383
rect 575 417 627 441
rect 609 383 627 417
rect 575 349 627 383
rect 17 215 31 249
rect 17 153 65 215
rect 99 299 537 333
rect 99 117 133 299
rect 474 265 537 299
rect 609 315 627 349
rect 34 101 133 117
rect 34 67 35 101
rect 69 67 133 101
rect 177 249 247 265
rect 211 215 247 249
rect 177 72 247 215
rect 283 249 343 265
rect 317 215 343 249
rect 283 71 343 215
rect 379 249 435 265
rect 413 215 435 249
rect 474 249 540 265
rect 474 215 490 249
rect 524 215 540 249
rect 379 71 435 215
rect 471 161 525 177
rect 575 161 627 315
rect 471 127 476 161
rect 510 127 525 161
rect 471 93 525 127
rect 34 51 133 67
rect 471 59 476 93
rect 510 59 525 93
rect 559 127 575 161
rect 609 127 627 161
rect 559 93 627 127
rect 559 59 575 93
rect 609 59 627 93
rect 471 17 525 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
flabel locali s 581 425 615 459 0 FreeSans 200 0 0 0 X
port 9 nsew signal output
flabel locali s 305 85 339 119 0 FreeSans 200 0 0 0 C
port 3 nsew signal input
flabel locali s 305 153 339 187 0 FreeSans 200 0 0 0 C
port 3 nsew signal input
flabel locali s 29 221 63 255 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 305 221 339 255 0 FreeSans 200 0 0 0 C
port 3 nsew signal input
flabel locali s 213 85 247 119 0 FreeSans 200 0 0 0 B
port 2 nsew signal input
flabel locali s 213 153 247 187 0 FreeSans 200 0 0 0 B
port 2 nsew signal input
flabel locali s 397 221 431 255 0 FreeSans 200 0 0 0 D
port 4 nsew signal input
flabel locali s 581 85 615 119 0 FreeSans 200 0 0 0 X
port 9 nsew signal output
flabel locali s 581 153 615 187 0 FreeSans 200 0 0 0 X
port 9 nsew signal output
flabel locali s 581 221 615 255 0 FreeSans 200 0 0 0 X
port 9 nsew signal output
flabel locali s 581 289 615 323 0 FreeSans 200 0 0 0 X
port 9 nsew signal output
flabel locali s 581 357 615 391 0 FreeSans 200 0 0 0 X
port 9 nsew signal output
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional abutment
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
rlabel comment s 0 0 0 0 4 and4_1
rlabel metal1 s 0 -48 644 48 1 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 496 644 592 1 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 644 544
string GDS_END 3904386
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3898032
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 16.100 0.000 
<< end >>
