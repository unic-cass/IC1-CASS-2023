magic
tech sky130B
magscale 1 2
timestamp 1676037725
<< nwell >>
rect -38 261 682 582
<< pwell >>
rect 1 21 643 203
rect 29 -17 63 21
<< locali >>
rect 17 73 73 493
rect 489 323 529 481
rect 463 289 529 323
rect 463 265 499 289
rect 196 215 267 265
rect 306 215 399 265
rect 433 215 499 265
rect 534 215 627 255
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 111 375 268 527
rect 347 361 424 493
rect 347 341 429 361
rect 107 299 429 341
rect 107 179 162 299
rect 563 291 627 527
rect 107 143 357 179
rect 284 129 357 143
rect 391 139 627 173
rect 119 17 153 109
rect 391 95 457 139
rect 207 59 457 95
rect 491 17 525 105
rect 559 56 627 139
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
rlabel locali s 534 215 627 255 6 A1
port 1 nsew signal input
rlabel locali s 433 215 499 265 6 A2
port 2 nsew signal input
rlabel locali s 463 265 499 289 6 A2
port 2 nsew signal input
rlabel locali s 463 289 529 323 6 A2
port 2 nsew signal input
rlabel locali s 489 323 529 481 6 A2
port 2 nsew signal input
rlabel locali s 196 215 267 265 6 B1
port 3 nsew signal input
rlabel locali s 306 215 399 265 6 B2
port 4 nsew signal input
rlabel metal1 s 0 -48 644 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 1 21 643 203 6 VNB
port 6 nsew ground bidirectional
rlabel nwell s -38 261 682 582 6 VPB
port 7 nsew power bidirectional
rlabel metal1 s 0 496 644 592 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 17 73 73 493 6 X
port 9 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 644 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 1358900
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1352882
<< end >>
