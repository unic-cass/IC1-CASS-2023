magic
tech sky130B
magscale 1 2
timestamp 1676037725
<< pwell >>
rect 15 163 1035 1225
<< mvnmos >>
rect 241 189 341 1199
rect 397 189 497 1199
rect 553 189 653 1199
rect 709 189 809 1199
<< mvndiff >>
rect 181 1187 241 1199
rect 181 1153 196 1187
rect 230 1153 241 1187
rect 181 1119 241 1153
rect 181 1085 196 1119
rect 230 1085 241 1119
rect 181 1051 241 1085
rect 181 1017 196 1051
rect 230 1017 241 1051
rect 181 983 241 1017
rect 181 949 196 983
rect 230 949 241 983
rect 181 915 241 949
rect 181 881 196 915
rect 230 881 241 915
rect 181 847 241 881
rect 181 813 196 847
rect 230 813 241 847
rect 181 779 241 813
rect 181 745 196 779
rect 230 745 241 779
rect 181 711 241 745
rect 181 677 196 711
rect 230 677 241 711
rect 181 643 241 677
rect 181 609 196 643
rect 230 609 241 643
rect 181 575 241 609
rect 181 541 196 575
rect 230 541 241 575
rect 181 507 241 541
rect 181 473 196 507
rect 230 473 241 507
rect 181 439 241 473
rect 181 405 196 439
rect 230 405 241 439
rect 181 371 241 405
rect 181 337 196 371
rect 230 337 241 371
rect 181 303 241 337
rect 181 269 196 303
rect 230 269 241 303
rect 181 235 241 269
rect 181 201 196 235
rect 230 201 241 235
rect 181 189 241 201
rect 341 1187 397 1199
rect 341 1153 352 1187
rect 386 1153 397 1187
rect 341 1119 397 1153
rect 341 1085 352 1119
rect 386 1085 397 1119
rect 341 1051 397 1085
rect 341 1017 352 1051
rect 386 1017 397 1051
rect 341 983 397 1017
rect 341 949 352 983
rect 386 949 397 983
rect 341 915 397 949
rect 341 881 352 915
rect 386 881 397 915
rect 341 847 397 881
rect 341 813 352 847
rect 386 813 397 847
rect 341 779 397 813
rect 341 745 352 779
rect 386 745 397 779
rect 341 711 397 745
rect 341 677 352 711
rect 386 677 397 711
rect 341 643 397 677
rect 341 609 352 643
rect 386 609 397 643
rect 341 575 397 609
rect 341 541 352 575
rect 386 541 397 575
rect 341 507 397 541
rect 341 473 352 507
rect 386 473 397 507
rect 341 439 397 473
rect 341 405 352 439
rect 386 405 397 439
rect 341 371 397 405
rect 341 337 352 371
rect 386 337 397 371
rect 341 303 397 337
rect 341 269 352 303
rect 386 269 397 303
rect 341 235 397 269
rect 341 201 352 235
rect 386 201 397 235
rect 341 189 397 201
rect 497 1187 553 1199
rect 497 1153 508 1187
rect 542 1153 553 1187
rect 497 1119 553 1153
rect 497 1085 508 1119
rect 542 1085 553 1119
rect 497 1051 553 1085
rect 497 1017 508 1051
rect 542 1017 553 1051
rect 497 983 553 1017
rect 497 949 508 983
rect 542 949 553 983
rect 497 915 553 949
rect 497 881 508 915
rect 542 881 553 915
rect 497 847 553 881
rect 497 813 508 847
rect 542 813 553 847
rect 497 779 553 813
rect 497 745 508 779
rect 542 745 553 779
rect 497 711 553 745
rect 497 677 508 711
rect 542 677 553 711
rect 497 643 553 677
rect 497 609 508 643
rect 542 609 553 643
rect 497 575 553 609
rect 497 541 508 575
rect 542 541 553 575
rect 497 507 553 541
rect 497 473 508 507
rect 542 473 553 507
rect 497 439 553 473
rect 497 405 508 439
rect 542 405 553 439
rect 497 371 553 405
rect 497 337 508 371
rect 542 337 553 371
rect 497 303 553 337
rect 497 269 508 303
rect 542 269 553 303
rect 497 235 553 269
rect 497 201 508 235
rect 542 201 553 235
rect 497 189 553 201
rect 653 1187 709 1199
rect 653 1153 664 1187
rect 698 1153 709 1187
rect 653 1119 709 1153
rect 653 1085 664 1119
rect 698 1085 709 1119
rect 653 1051 709 1085
rect 653 1017 664 1051
rect 698 1017 709 1051
rect 653 983 709 1017
rect 653 949 664 983
rect 698 949 709 983
rect 653 915 709 949
rect 653 881 664 915
rect 698 881 709 915
rect 653 847 709 881
rect 653 813 664 847
rect 698 813 709 847
rect 653 779 709 813
rect 653 745 664 779
rect 698 745 709 779
rect 653 711 709 745
rect 653 677 664 711
rect 698 677 709 711
rect 653 643 709 677
rect 653 609 664 643
rect 698 609 709 643
rect 653 575 709 609
rect 653 541 664 575
rect 698 541 709 575
rect 653 507 709 541
rect 653 473 664 507
rect 698 473 709 507
rect 653 439 709 473
rect 653 405 664 439
rect 698 405 709 439
rect 653 371 709 405
rect 653 337 664 371
rect 698 337 709 371
rect 653 303 709 337
rect 653 269 664 303
rect 698 269 709 303
rect 653 235 709 269
rect 653 201 664 235
rect 698 201 709 235
rect 653 189 709 201
rect 809 1187 869 1199
rect 809 1153 820 1187
rect 854 1153 869 1187
rect 809 1119 869 1153
rect 809 1085 820 1119
rect 854 1085 869 1119
rect 809 1051 869 1085
rect 809 1017 820 1051
rect 854 1017 869 1051
rect 809 983 869 1017
rect 809 949 820 983
rect 854 949 869 983
rect 809 915 869 949
rect 809 881 820 915
rect 854 881 869 915
rect 809 847 869 881
rect 809 813 820 847
rect 854 813 869 847
rect 809 779 869 813
rect 809 745 820 779
rect 854 745 869 779
rect 809 711 869 745
rect 809 677 820 711
rect 854 677 869 711
rect 809 643 869 677
rect 809 609 820 643
rect 854 609 869 643
rect 809 575 869 609
rect 809 541 820 575
rect 854 541 869 575
rect 809 507 869 541
rect 809 473 820 507
rect 854 473 869 507
rect 809 439 869 473
rect 809 405 820 439
rect 854 405 869 439
rect 809 371 869 405
rect 809 337 820 371
rect 854 337 869 371
rect 809 303 869 337
rect 809 269 820 303
rect 854 269 869 303
rect 809 235 869 269
rect 809 201 820 235
rect 854 201 869 235
rect 809 189 869 201
<< mvndiffc >>
rect 196 1153 230 1187
rect 196 1085 230 1119
rect 196 1017 230 1051
rect 196 949 230 983
rect 196 881 230 915
rect 196 813 230 847
rect 196 745 230 779
rect 196 677 230 711
rect 196 609 230 643
rect 196 541 230 575
rect 196 473 230 507
rect 196 405 230 439
rect 196 337 230 371
rect 196 269 230 303
rect 196 201 230 235
rect 352 1153 386 1187
rect 352 1085 386 1119
rect 352 1017 386 1051
rect 352 949 386 983
rect 352 881 386 915
rect 352 813 386 847
rect 352 745 386 779
rect 352 677 386 711
rect 352 609 386 643
rect 352 541 386 575
rect 352 473 386 507
rect 352 405 386 439
rect 352 337 386 371
rect 352 269 386 303
rect 352 201 386 235
rect 508 1153 542 1187
rect 508 1085 542 1119
rect 508 1017 542 1051
rect 508 949 542 983
rect 508 881 542 915
rect 508 813 542 847
rect 508 745 542 779
rect 508 677 542 711
rect 508 609 542 643
rect 508 541 542 575
rect 508 473 542 507
rect 508 405 542 439
rect 508 337 542 371
rect 508 269 542 303
rect 508 201 542 235
rect 664 1153 698 1187
rect 664 1085 698 1119
rect 664 1017 698 1051
rect 664 949 698 983
rect 664 881 698 915
rect 664 813 698 847
rect 664 745 698 779
rect 664 677 698 711
rect 664 609 698 643
rect 664 541 698 575
rect 664 473 698 507
rect 664 405 698 439
rect 664 337 698 371
rect 664 269 698 303
rect 664 201 698 235
rect 820 1153 854 1187
rect 820 1085 854 1119
rect 820 1017 854 1051
rect 820 949 854 983
rect 820 881 854 915
rect 820 813 854 847
rect 820 745 854 779
rect 820 677 854 711
rect 820 609 854 643
rect 820 541 854 575
rect 820 473 854 507
rect 820 405 854 439
rect 820 337 854 371
rect 820 269 854 303
rect 820 201 854 235
<< mvpsubdiff >>
rect 41 1187 181 1199
rect 41 201 60 1187
rect 162 201 181 1187
rect 41 189 181 201
rect 869 1187 1009 1199
rect 869 201 888 1187
rect 990 201 1009 1187
rect 869 189 1009 201
<< mvpsubdiffcont >>
rect 60 201 162 1187
rect 888 201 990 1187
<< poly >>
rect 383 1367 667 1388
rect 190 1275 341 1291
rect 190 1241 206 1275
rect 240 1241 341 1275
rect 383 1265 406 1367
rect 644 1265 667 1367
rect 383 1249 667 1265
rect 709 1275 860 1291
rect 190 1225 341 1241
rect 241 1199 341 1225
rect 397 1199 497 1249
rect 553 1199 653 1249
rect 709 1241 810 1275
rect 844 1241 860 1275
rect 709 1225 860 1241
rect 709 1199 809 1225
rect 241 163 341 189
rect 190 147 341 163
rect 190 113 206 147
rect 240 113 341 147
rect 397 139 497 189
rect 553 139 653 189
rect 709 163 809 189
rect 709 147 860 163
rect 190 97 341 113
rect 383 123 667 139
rect 383 21 406 123
rect 644 21 667 123
rect 709 113 810 147
rect 844 113 860 147
rect 709 97 860 113
rect 383 0 667 21
<< polycont >>
rect 206 1241 240 1275
rect 406 1265 644 1367
rect 810 1241 844 1275
rect 206 113 240 147
rect 406 21 644 123
rect 810 113 844 147
<< locali >>
rect 383 1369 667 1388
rect 190 1275 256 1291
rect 190 1241 206 1275
rect 240 1241 256 1275
rect 383 1263 400 1369
rect 650 1263 667 1369
rect 383 1251 667 1263
rect 794 1275 860 1291
rect 190 1225 256 1241
rect 794 1241 810 1275
rect 844 1241 860 1275
rect 794 1225 860 1241
rect 190 1203 230 1225
rect 820 1203 860 1225
rect 41 1187 230 1203
rect 41 201 60 1187
rect 162 1153 196 1187
rect 162 1119 230 1153
rect 162 1085 196 1119
rect 162 1051 230 1085
rect 162 1017 196 1051
rect 162 983 230 1017
rect 162 949 196 983
rect 162 915 230 949
rect 162 881 196 915
rect 162 847 230 881
rect 162 813 196 847
rect 162 779 230 813
rect 162 745 196 779
rect 162 711 230 745
rect 162 677 196 711
rect 162 643 230 677
rect 162 609 196 643
rect 162 575 230 609
rect 162 541 196 575
rect 162 507 230 541
rect 162 473 196 507
rect 162 439 230 473
rect 162 405 196 439
rect 162 371 230 405
rect 162 337 196 371
rect 162 303 230 337
rect 162 269 196 303
rect 162 235 230 269
rect 162 201 196 235
rect 41 185 230 201
rect 352 1187 386 1203
rect 352 1119 386 1145
rect 352 1051 386 1073
rect 352 983 386 1001
rect 352 915 386 929
rect 352 847 386 857
rect 352 779 386 785
rect 352 711 386 713
rect 352 675 386 677
rect 352 603 386 609
rect 352 531 386 541
rect 352 459 386 473
rect 352 387 386 405
rect 352 315 386 337
rect 352 243 386 269
rect 352 185 386 201
rect 508 1187 542 1203
rect 508 1119 542 1145
rect 508 1051 542 1073
rect 508 983 542 1001
rect 508 915 542 929
rect 508 847 542 857
rect 508 779 542 785
rect 508 711 542 713
rect 508 675 542 677
rect 508 603 542 609
rect 508 531 542 541
rect 508 459 542 473
rect 508 387 542 405
rect 508 315 542 337
rect 508 243 542 269
rect 508 185 542 201
rect 664 1187 698 1203
rect 664 1119 698 1145
rect 664 1051 698 1073
rect 664 983 698 1001
rect 664 915 698 929
rect 664 847 698 857
rect 664 779 698 785
rect 664 711 698 713
rect 664 675 698 677
rect 664 603 698 609
rect 664 531 698 541
rect 664 459 698 473
rect 664 387 698 405
rect 664 315 698 337
rect 664 243 698 269
rect 664 185 698 201
rect 820 1187 1009 1203
rect 854 1153 888 1187
rect 820 1119 888 1153
rect 854 1085 888 1119
rect 820 1051 888 1085
rect 854 1017 888 1051
rect 820 983 888 1017
rect 854 949 888 983
rect 820 915 888 949
rect 854 881 888 915
rect 820 847 888 881
rect 854 813 888 847
rect 820 779 888 813
rect 854 745 888 779
rect 820 711 888 745
rect 854 677 888 711
rect 820 643 888 677
rect 854 609 888 643
rect 820 575 888 609
rect 854 541 888 575
rect 820 507 888 541
rect 854 473 888 507
rect 820 439 888 473
rect 854 405 888 439
rect 820 371 888 405
rect 854 337 888 371
rect 820 303 888 337
rect 854 269 888 303
rect 820 235 888 269
rect 854 201 888 235
rect 990 201 1009 1187
rect 820 185 1009 201
rect 190 163 230 185
rect 820 163 860 185
rect 190 147 256 163
rect 190 113 206 147
rect 240 113 256 147
rect 794 147 860 163
rect 190 97 256 113
rect 383 125 667 137
rect 383 19 400 125
rect 650 19 667 125
rect 794 113 810 147
rect 844 113 860 147
rect 794 97 860 113
rect 383 0 667 19
<< viali >>
rect 400 1367 650 1369
rect 400 1265 406 1367
rect 406 1265 644 1367
rect 644 1265 650 1367
rect 400 1263 650 1265
rect 60 1145 94 1179
rect 60 1073 94 1107
rect 60 1001 94 1035
rect 60 929 94 963
rect 60 857 94 891
rect 60 785 94 819
rect 60 713 94 747
rect 60 641 94 675
rect 60 569 94 603
rect 60 497 94 531
rect 60 425 94 459
rect 60 353 94 387
rect 60 281 94 315
rect 60 209 94 243
rect 352 1153 386 1179
rect 352 1145 386 1153
rect 352 1085 386 1107
rect 352 1073 386 1085
rect 352 1017 386 1035
rect 352 1001 386 1017
rect 352 949 386 963
rect 352 929 386 949
rect 352 881 386 891
rect 352 857 386 881
rect 352 813 386 819
rect 352 785 386 813
rect 352 745 386 747
rect 352 713 386 745
rect 352 643 386 675
rect 352 641 386 643
rect 352 575 386 603
rect 352 569 386 575
rect 352 507 386 531
rect 352 497 386 507
rect 352 439 386 459
rect 352 425 386 439
rect 352 371 386 387
rect 352 353 386 371
rect 352 303 386 315
rect 352 281 386 303
rect 352 235 386 243
rect 352 209 386 235
rect 508 1153 542 1179
rect 508 1145 542 1153
rect 508 1085 542 1107
rect 508 1073 542 1085
rect 508 1017 542 1035
rect 508 1001 542 1017
rect 508 949 542 963
rect 508 929 542 949
rect 508 881 542 891
rect 508 857 542 881
rect 508 813 542 819
rect 508 785 542 813
rect 508 745 542 747
rect 508 713 542 745
rect 508 643 542 675
rect 508 641 542 643
rect 508 575 542 603
rect 508 569 542 575
rect 508 507 542 531
rect 508 497 542 507
rect 508 439 542 459
rect 508 425 542 439
rect 508 371 542 387
rect 508 353 542 371
rect 508 303 542 315
rect 508 281 542 303
rect 508 235 542 243
rect 508 209 542 235
rect 664 1153 698 1179
rect 664 1145 698 1153
rect 664 1085 698 1107
rect 664 1073 698 1085
rect 664 1017 698 1035
rect 664 1001 698 1017
rect 664 949 698 963
rect 664 929 698 949
rect 664 881 698 891
rect 664 857 698 881
rect 664 813 698 819
rect 664 785 698 813
rect 664 745 698 747
rect 664 713 698 745
rect 664 643 698 675
rect 664 641 698 643
rect 664 575 698 603
rect 664 569 698 575
rect 664 507 698 531
rect 664 497 698 507
rect 664 439 698 459
rect 664 425 698 439
rect 664 371 698 387
rect 664 353 698 371
rect 664 303 698 315
rect 664 281 698 303
rect 664 235 698 243
rect 664 209 698 235
rect 956 1145 990 1179
rect 956 1073 990 1107
rect 956 1001 990 1035
rect 956 929 990 963
rect 956 857 990 891
rect 956 785 990 819
rect 956 713 990 747
rect 956 641 990 675
rect 956 569 990 603
rect 956 497 990 531
rect 956 425 990 459
rect 956 353 990 387
rect 956 281 990 315
rect 956 209 990 243
rect 400 123 650 125
rect 400 21 406 123
rect 406 21 644 123
rect 644 21 650 123
rect 400 19 650 21
<< metal1 >>
rect 380 1369 670 1388
rect 380 1263 400 1369
rect 650 1263 670 1369
rect 380 1251 670 1263
rect 41 1179 100 1191
rect 41 1145 60 1179
rect 94 1145 100 1179
rect 41 1107 100 1145
rect 41 1073 60 1107
rect 94 1073 100 1107
rect 41 1035 100 1073
rect 41 1001 60 1035
rect 94 1001 100 1035
rect 41 963 100 1001
rect 41 929 60 963
rect 94 929 100 963
rect 41 891 100 929
rect 41 857 60 891
rect 94 857 100 891
rect 41 819 100 857
rect 41 785 60 819
rect 94 785 100 819
rect 41 747 100 785
rect 41 713 60 747
rect 94 713 100 747
rect 41 675 100 713
rect 41 641 60 675
rect 94 641 100 675
rect 41 603 100 641
rect 41 569 60 603
rect 94 569 100 603
rect 41 531 100 569
rect 41 497 60 531
rect 94 497 100 531
rect 41 459 100 497
rect 41 425 60 459
rect 94 425 100 459
rect 41 387 100 425
rect 41 353 60 387
rect 94 353 100 387
rect 41 315 100 353
rect 41 281 60 315
rect 94 281 100 315
rect 41 243 100 281
rect 41 209 60 243
rect 94 209 100 243
rect 41 197 100 209
rect 343 1179 395 1191
rect 343 1145 352 1179
rect 386 1145 395 1179
rect 343 1107 395 1145
rect 343 1073 352 1107
rect 386 1073 395 1107
rect 343 1035 395 1073
rect 343 1001 352 1035
rect 386 1001 395 1035
rect 343 963 395 1001
rect 343 929 352 963
rect 386 929 395 963
rect 343 891 395 929
rect 343 857 352 891
rect 386 857 395 891
rect 343 819 395 857
rect 343 785 352 819
rect 386 785 395 819
rect 343 747 395 785
rect 343 713 352 747
rect 386 713 395 747
rect 343 675 395 713
rect 343 641 352 675
rect 386 641 395 675
rect 343 639 395 641
rect 343 575 352 587
rect 386 575 395 587
rect 343 511 352 523
rect 386 511 395 523
rect 343 447 352 459
rect 386 447 395 459
rect 343 387 395 395
rect 343 383 352 387
rect 386 383 395 387
rect 343 319 395 331
rect 343 255 395 267
rect 343 197 395 203
rect 499 1185 551 1191
rect 499 1121 551 1133
rect 499 1057 551 1069
rect 499 1001 508 1005
rect 542 1001 551 1005
rect 499 993 551 1001
rect 499 929 508 941
rect 542 929 551 941
rect 499 865 508 877
rect 542 865 551 877
rect 499 801 508 813
rect 542 801 551 813
rect 499 747 551 749
rect 499 713 508 747
rect 542 713 551 747
rect 499 675 551 713
rect 499 641 508 675
rect 542 641 551 675
rect 499 603 551 641
rect 499 569 508 603
rect 542 569 551 603
rect 499 531 551 569
rect 499 497 508 531
rect 542 497 551 531
rect 499 459 551 497
rect 499 425 508 459
rect 542 425 551 459
rect 499 387 551 425
rect 499 353 508 387
rect 542 353 551 387
rect 499 315 551 353
rect 499 281 508 315
rect 542 281 551 315
rect 499 243 551 281
rect 499 209 508 243
rect 542 209 551 243
rect 499 197 551 209
rect 655 1179 707 1191
rect 655 1145 664 1179
rect 698 1145 707 1179
rect 655 1107 707 1145
rect 655 1073 664 1107
rect 698 1073 707 1107
rect 655 1035 707 1073
rect 655 1001 664 1035
rect 698 1001 707 1035
rect 655 963 707 1001
rect 655 929 664 963
rect 698 929 707 963
rect 655 891 707 929
rect 655 857 664 891
rect 698 857 707 891
rect 655 819 707 857
rect 655 785 664 819
rect 698 785 707 819
rect 655 747 707 785
rect 655 713 664 747
rect 698 713 707 747
rect 655 675 707 713
rect 655 641 664 675
rect 698 641 707 675
rect 655 639 707 641
rect 655 575 664 587
rect 698 575 707 587
rect 655 511 664 523
rect 698 511 707 523
rect 655 447 664 459
rect 698 447 707 459
rect 655 387 707 395
rect 655 383 664 387
rect 698 383 707 387
rect 655 319 707 331
rect 655 255 707 267
rect 655 197 707 203
rect 950 1179 1009 1191
rect 950 1145 956 1179
rect 990 1145 1009 1179
rect 950 1107 1009 1145
rect 950 1073 956 1107
rect 990 1073 1009 1107
rect 950 1035 1009 1073
rect 950 1001 956 1035
rect 990 1001 1009 1035
rect 950 963 1009 1001
rect 950 929 956 963
rect 990 929 1009 963
rect 950 891 1009 929
rect 950 857 956 891
rect 990 857 1009 891
rect 950 819 1009 857
rect 950 785 956 819
rect 990 785 1009 819
rect 950 747 1009 785
rect 950 713 956 747
rect 990 713 1009 747
rect 950 675 1009 713
rect 950 641 956 675
rect 990 641 1009 675
rect 950 603 1009 641
rect 950 569 956 603
rect 990 569 1009 603
rect 950 531 1009 569
rect 950 497 956 531
rect 990 497 1009 531
rect 950 459 1009 497
rect 950 425 956 459
rect 990 425 1009 459
rect 950 387 1009 425
rect 950 353 956 387
rect 990 353 1009 387
rect 950 315 1009 353
rect 950 281 956 315
rect 990 281 1009 315
rect 950 243 1009 281
rect 950 209 956 243
rect 990 209 1009 243
rect 950 197 1009 209
rect 380 125 670 137
rect 380 19 400 125
rect 650 19 670 125
rect 380 0 670 19
<< via1 >>
rect 343 603 395 639
rect 343 587 352 603
rect 352 587 386 603
rect 386 587 395 603
rect 343 569 352 575
rect 352 569 386 575
rect 386 569 395 575
rect 343 531 395 569
rect 343 523 352 531
rect 352 523 386 531
rect 386 523 395 531
rect 343 497 352 511
rect 352 497 386 511
rect 386 497 395 511
rect 343 459 395 497
rect 343 425 352 447
rect 352 425 386 447
rect 386 425 395 447
rect 343 395 395 425
rect 343 353 352 383
rect 352 353 386 383
rect 386 353 395 383
rect 343 331 395 353
rect 343 315 395 319
rect 343 281 352 315
rect 352 281 386 315
rect 386 281 395 315
rect 343 267 395 281
rect 343 243 395 255
rect 343 209 352 243
rect 352 209 386 243
rect 386 209 395 243
rect 343 203 395 209
rect 499 1179 551 1185
rect 499 1145 508 1179
rect 508 1145 542 1179
rect 542 1145 551 1179
rect 499 1133 551 1145
rect 499 1107 551 1121
rect 499 1073 508 1107
rect 508 1073 542 1107
rect 542 1073 551 1107
rect 499 1069 551 1073
rect 499 1035 551 1057
rect 499 1005 508 1035
rect 508 1005 542 1035
rect 542 1005 551 1035
rect 499 963 551 993
rect 499 941 508 963
rect 508 941 542 963
rect 542 941 551 963
rect 499 891 551 929
rect 499 877 508 891
rect 508 877 542 891
rect 542 877 551 891
rect 499 857 508 865
rect 508 857 542 865
rect 542 857 551 865
rect 499 819 551 857
rect 499 813 508 819
rect 508 813 542 819
rect 542 813 551 819
rect 499 785 508 801
rect 508 785 542 801
rect 542 785 551 801
rect 499 749 551 785
rect 655 603 707 639
rect 655 587 664 603
rect 664 587 698 603
rect 698 587 707 603
rect 655 569 664 575
rect 664 569 698 575
rect 698 569 707 575
rect 655 531 707 569
rect 655 523 664 531
rect 664 523 698 531
rect 698 523 707 531
rect 655 497 664 511
rect 664 497 698 511
rect 698 497 707 511
rect 655 459 707 497
rect 655 425 664 447
rect 664 425 698 447
rect 698 425 707 447
rect 655 395 707 425
rect 655 353 664 383
rect 664 353 698 383
rect 698 353 707 383
rect 655 331 707 353
rect 655 315 707 319
rect 655 281 664 315
rect 664 281 698 315
rect 698 281 707 315
rect 655 267 707 281
rect 655 243 707 255
rect 655 209 664 243
rect 664 209 698 243
rect 698 209 707 243
rect 655 203 707 209
<< metal2 >>
rect 14 1185 1036 1191
rect 14 1133 499 1185
rect 551 1133 1036 1185
rect 14 1121 1036 1133
rect 14 1069 499 1121
rect 551 1069 1036 1121
rect 14 1057 1036 1069
rect 14 1005 499 1057
rect 551 1005 1036 1057
rect 14 993 1036 1005
rect 14 941 499 993
rect 551 941 1036 993
rect 14 929 1036 941
rect 14 877 499 929
rect 551 877 1036 929
rect 14 865 1036 877
rect 14 813 499 865
rect 551 813 1036 865
rect 14 801 1036 813
rect 14 749 499 801
rect 551 749 1036 801
rect 14 719 1036 749
rect 14 639 1036 669
rect 14 587 343 639
rect 395 587 655 639
rect 707 587 1036 639
rect 14 575 1036 587
rect 14 523 343 575
rect 395 523 655 575
rect 707 523 1036 575
rect 14 511 1036 523
rect 14 459 343 511
rect 395 459 655 511
rect 707 459 1036 511
rect 14 447 1036 459
rect 14 395 343 447
rect 395 395 655 447
rect 707 395 1036 447
rect 14 383 1036 395
rect 14 331 343 383
rect 395 331 655 383
rect 707 331 1036 383
rect 14 319 1036 331
rect 14 267 343 319
rect 395 267 655 319
rect 707 267 1036 319
rect 14 255 1036 267
rect 14 203 343 255
rect 395 203 655 255
rect 707 203 1036 255
rect 14 197 1036 203
<< labels >>
flabel metal1 s 470 85 568 119 0 FreeSans 200 0 0 0 GATE
port 2 nsew
flabel metal1 s 470 1263 568 1297 0 FreeSans 400 0 0 0 GATE
port 2 nsew
flabel metal1 s 950 679 1009 709 0 FreeSans 200 90 0 0 SUBSTRATE
port 4 nsew
flabel metal1 s 41 675 100 705 0 FreeSans 200 90 0 0 SUBSTRATE
port 4 nsew
flabel comment s 369 694 369 694 0 FreeSans 300 0 0 0 S
flabel comment s 369 694 369 694 0 FreeSans 300 0 0 0 S
flabel comment s 525 694 525 694 0 FreeSans 300 0 0 0 S
flabel comment s 525 694 525 694 0 FreeSans 300 0 0 0 D
flabel comment s 681 694 681 694 0 FreeSans 300 0 0 0 S
flabel comment s 681 694 681 694 0 FreeSans 300 0 0 0 S
flabel comment s 283 681 283 681 0 FreeSans 400 90 0 0 dummy_poly
flabel comment s 751 707 751 707 0 FreeSans 400 90 0 0 dummy_poly
flabel metal2 s 26 442 128 488 0 FreeSans 200 0 0 0 SOURCE
port 3 nsew
flabel metal2 s 26 991 137 1048 0 FreeSans 200 0 0 0 DRAIN
port 1 nsew
<< properties >>
string GDS_END 8463040
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 8440388
string device primitive
<< end >>
