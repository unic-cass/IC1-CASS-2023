magic
tech sky130A
magscale 1 2
timestamp 1676037725
use sky130_fd_pr__hvdfl1sd__example_55959141808100  sky130_fd_pr__hvdfl1sd__example_55959141808100_0
timestamp 1676037725
transform -1 0 0 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 32491180
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 32490324
<< end >>
