magic
tech sky130A
magscale 1 2
timestamp 1676037725
<< nwell >>
rect -54 784 204 1454
rect -59 616 209 784
rect -54 -54 204 616
<< scpmos >>
rect 60 0 90 1400
<< pdiff >>
rect 0 717 60 1400
rect 0 683 8 717
rect 42 683 60 717
rect 0 0 60 683
rect 90 717 150 1400
rect 90 683 108 717
rect 142 683 150 717
rect 90 0 150 683
<< pdiffc >>
rect 8 683 42 717
rect 108 683 142 717
<< poly >>
rect 60 1400 90 1426
rect 60 -26 90 0
<< locali >>
rect 8 717 42 733
rect 8 667 42 683
rect 108 717 142 733
rect 108 667 142 683
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_12  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_12_0
timestamp 1676037725
transform 1 0 100 0 1 667
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_12  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_12_1
timestamp 1676037725
transform 1 0 0 0 1 667
box 0 0 1 1
<< labels >>
rlabel locali s 25 700 25 700 4 S
rlabel locali s 125 700 125 700 4 D
rlabel poly s 75 700 75 700 4 G
<< properties >>
string FIXED_BBOX -54 -54 204 616
string GDS_END 9932
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_1kbyte_1rw1r_8x1024_8.gds
string GDS_START 9072
<< end >>
