magic
tech sky130A
magscale 1 2
timestamp 1676037725
<< locali >>
rect 165 752 177 786
rect 211 752 249 786
rect 283 752 321 786
rect 355 752 393 786
rect 427 752 439 786
rect 48 672 82 674
rect 48 600 82 638
rect 48 528 82 566
rect 48 456 82 494
rect 48 384 82 422
rect 48 312 82 350
rect 48 240 82 278
rect 48 168 82 206
rect 48 132 82 134
rect 522 672 556 674
rect 522 600 556 638
rect 522 528 556 566
rect 522 456 556 494
rect 522 384 556 422
rect 522 312 556 350
rect 522 240 556 278
rect 522 168 556 206
rect 522 132 556 134
rect 165 20 177 54
rect 211 20 249 54
rect 283 20 321 54
rect 355 20 393 54
rect 427 20 439 54
<< viali >>
rect 177 752 211 786
rect 249 752 283 786
rect 321 752 355 786
rect 393 752 427 786
rect 48 638 82 672
rect 48 566 82 600
rect 48 494 82 528
rect 48 422 82 456
rect 48 350 82 384
rect 48 278 82 312
rect 48 206 82 240
rect 48 134 82 168
rect 522 638 556 672
rect 522 566 556 600
rect 522 494 556 528
rect 522 422 556 456
rect 522 350 556 384
rect 522 278 556 312
rect 522 206 556 240
rect 522 134 556 168
rect 177 20 211 54
rect 249 20 283 54
rect 321 20 355 54
rect 393 20 427 54
<< obsli1 >>
rect 159 98 193 708
rect 285 98 319 708
rect 411 98 445 708
<< metal1 >>
rect 165 786 439 806
rect 165 752 177 786
rect 211 752 249 786
rect 283 752 321 786
rect 355 752 393 786
rect 427 752 439 786
rect 165 740 439 752
rect 36 672 94 684
rect 36 638 48 672
rect 82 638 94 672
rect 36 600 94 638
rect 36 566 48 600
rect 82 566 94 600
rect 36 528 94 566
rect 36 494 48 528
rect 82 494 94 528
rect 36 456 94 494
rect 36 422 48 456
rect 82 422 94 456
rect 36 384 94 422
rect 36 350 48 384
rect 82 350 94 384
rect 36 312 94 350
rect 36 278 48 312
rect 82 278 94 312
rect 36 240 94 278
rect 36 206 48 240
rect 82 206 94 240
rect 36 168 94 206
rect 36 134 48 168
rect 82 134 94 168
rect 36 122 94 134
rect 510 672 568 684
rect 510 638 522 672
rect 556 638 568 672
rect 510 600 568 638
rect 510 566 522 600
rect 556 566 568 600
rect 510 528 568 566
rect 510 494 522 528
rect 556 494 568 528
rect 510 456 568 494
rect 510 422 522 456
rect 556 422 568 456
rect 510 384 568 422
rect 510 350 522 384
rect 556 350 568 384
rect 510 312 568 350
rect 510 278 522 312
rect 556 278 568 312
rect 510 240 568 278
rect 510 206 522 240
rect 556 206 568 240
rect 510 168 568 206
rect 510 134 522 168
rect 556 134 568 168
rect 510 122 568 134
rect 165 54 439 66
rect 165 20 177 54
rect 211 20 249 54
rect 283 20 321 54
rect 355 20 393 54
rect 427 20 439 54
rect 165 0 439 20
<< obsm1 >>
rect 150 122 202 684
rect 276 122 328 684
rect 402 122 454 684
<< metal2 >>
rect 10 428 594 684
rect 10 122 594 378
<< labels >>
rlabel viali s 522 638 556 672 6 BULK
port 1 nsew
rlabel viali s 522 566 556 600 6 BULK
port 1 nsew
rlabel viali s 522 494 556 528 6 BULK
port 1 nsew
rlabel viali s 522 422 556 456 6 BULK
port 1 nsew
rlabel viali s 522 350 556 384 6 BULK
port 1 nsew
rlabel viali s 522 278 556 312 6 BULK
port 1 nsew
rlabel viali s 522 206 556 240 6 BULK
port 1 nsew
rlabel viali s 522 134 556 168 6 BULK
port 1 nsew
rlabel viali s 48 638 82 672 6 BULK
port 1 nsew
rlabel viali s 48 566 82 600 6 BULK
port 1 nsew
rlabel viali s 48 494 82 528 6 BULK
port 1 nsew
rlabel viali s 48 422 82 456 6 BULK
port 1 nsew
rlabel viali s 48 350 82 384 6 BULK
port 1 nsew
rlabel viali s 48 278 82 312 6 BULK
port 1 nsew
rlabel viali s 48 206 82 240 6 BULK
port 1 nsew
rlabel viali s 48 134 82 168 6 BULK
port 1 nsew
rlabel locali s 522 132 556 674 6 BULK
port 1 nsew
rlabel locali s 48 132 82 674 6 BULK
port 1 nsew
rlabel metal1 s 510 122 568 684 6 BULK
port 1 nsew
rlabel metal1 s 36 122 94 684 6 BULK
port 1 nsew
rlabel metal2 s 10 428 594 684 6 DRAIN
port 2 nsew
rlabel viali s 393 752 427 786 6 GATE
port 3 nsew
rlabel viali s 393 20 427 54 6 GATE
port 3 nsew
rlabel viali s 321 752 355 786 6 GATE
port 3 nsew
rlabel viali s 321 20 355 54 6 GATE
port 3 nsew
rlabel viali s 249 752 283 786 6 GATE
port 3 nsew
rlabel viali s 249 20 283 54 6 GATE
port 3 nsew
rlabel viali s 177 752 211 786 6 GATE
port 3 nsew
rlabel viali s 177 20 211 54 6 GATE
port 3 nsew
rlabel locali s 165 752 439 786 6 GATE
port 3 nsew
rlabel locali s 165 20 439 54 6 GATE
port 3 nsew
rlabel metal1 s 165 740 439 806 6 GATE
port 3 nsew
rlabel metal1 s 165 0 439 66 6 GATE
port 3 nsew
rlabel metal2 s 10 122 594 378 6 SOURCE
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 604 806
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 9849686
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 9838578
<< end >>
