magic
tech sky130A
magscale 1 2
timestamp 1676037725
<< locali >>
rect 12165 1381 12231 1473
rect 12178 1347 12216 1381
<< viali >>
rect 12144 1347 12178 1381
rect 12216 1347 12250 1381
<< metal1 >>
rect 2787 2731 3539 2732
rect 2787 2679 2793 2731
rect 2845 2679 2892 2731
rect 2944 2679 2991 2731
rect 3043 2679 3089 2731
rect 3141 2679 3187 2731
rect 3239 2679 3285 2731
rect 3337 2679 3383 2731
rect 3435 2679 3481 2731
rect 3533 2679 3539 2731
rect 2787 2643 3539 2679
rect 2787 2591 2793 2643
rect 2845 2591 2892 2643
rect 2944 2591 2991 2643
rect 3043 2591 3089 2643
rect 3141 2591 3187 2643
rect 3239 2591 3285 2643
rect 3337 2591 3383 2643
rect 3435 2591 3481 2643
rect 3533 2591 3539 2643
rect 2787 2555 3539 2591
rect 5273 2579 5506 2710
rect 2787 2503 2793 2555
rect 2845 2503 2892 2555
rect 2944 2503 2991 2555
rect 3043 2503 3089 2555
rect 3141 2503 3187 2555
rect 3239 2503 3285 2555
rect 3337 2503 3383 2555
rect 3435 2503 3481 2555
rect 3533 2503 3539 2555
rect 2787 2502 3539 2503
rect 11522 2498 11542 2700
rect 12400 2498 12458 2700
rect 14371 2498 14400 2700
rect 11522 2424 11542 2470
rect 12400 2424 12458 2470
rect 14371 2424 14400 2470
rect 3224 2201 3334 2247
rect 3689 2037 3741 2043
rect 3689 1973 3741 1985
rect 2858 1906 2864 1958
rect 2916 1906 2928 1958
rect 2980 1906 2986 1958
rect 3122 1905 3128 1957
rect 3180 1905 3198 1957
rect 3250 1905 3267 1957
rect 3319 1905 3336 1957
rect 3388 1905 3394 1957
rect 11555 1972 11581 2248
rect 12400 1972 12429 2248
rect 14371 1972 14400 2248
tri 3667 1895 3689 1917 se
rect 3689 1895 3741 1921
rect 3879 1906 3885 1958
rect 3937 1906 3949 1958
rect 4001 1906 4007 1958
tri 3638 1866 3667 1895 se
rect 3236 1814 3242 1866
rect 3294 1814 3306 1866
rect 3358 1821 3667 1866
tri 3667 1821 3741 1895 nw
rect 4887 1880 4893 1932
rect 4945 1880 4957 1932
rect 5009 1880 5015 1932
rect 11142 1904 12092 1944
rect 10588 1821 10594 1873
rect 10646 1821 10658 1873
rect 10710 1821 10716 1873
rect 10843 1821 10849 1873
rect 10901 1821 10913 1873
rect 10965 1821 10971 1873
rect 3358 1814 3660 1821
tri 3660 1814 3667 1821 nw
rect 7703 1643 7781 1749
rect 10633 1720 10685 1821
rect 10578 1668 10584 1720
rect 10636 1668 10648 1720
rect 10700 1668 10706 1720
rect 10843 1707 10971 1821
rect 2773 1578 2779 1630
rect 2831 1578 2864 1630
rect 2916 1578 2949 1630
rect 3001 1578 3007 1630
rect 2773 1558 3007 1578
rect 2773 1506 2779 1558
rect 2831 1506 2864 1558
rect 2916 1506 2949 1558
rect 3001 1506 3007 1558
rect 3061 1511 3294 1626
rect 7685 1591 7691 1643
rect 7743 1591 7755 1643
rect 7807 1591 7813 1643
rect 10843 1639 10942 1707
tri 10942 1678 10971 1707 nw
rect 4449 1500 4455 1552
rect 4507 1500 4525 1552
rect 4577 1500 4595 1552
rect 4647 1500 4665 1552
rect 4717 1500 4735 1552
rect 4787 1500 4805 1552
rect 4857 1500 4875 1552
rect 4927 1500 4944 1552
rect 4996 1500 5002 1552
rect 8613 1547 8663 1593
rect 10814 1587 10820 1639
rect 10872 1587 10884 1639
rect 10936 1587 10942 1639
rect 5354 1505 5412 1547
rect 10820 1452 10872 1458
rect 11142 1427 11182 1904
rect 10872 1400 11182 1427
rect 10820 1388 11182 1400
rect 10872 1387 11182 1388
rect 11248 1837 11300 1843
rect 13410 1819 13416 1871
rect 13468 1819 13480 1871
rect 13532 1819 13538 1871
rect 11248 1773 11300 1785
rect 13467 1734 13473 1786
rect 13525 1734 13537 1786
rect 13589 1734 13595 1786
rect 11248 1387 11300 1721
rect 13467 1654 13473 1706
rect 13525 1654 13537 1706
rect 13589 1654 13595 1706
rect 14219 1574 14225 1626
rect 14277 1574 14289 1626
rect 14341 1574 14347 1626
rect 12939 1520 12978 1541
rect 12679 1475 12721 1503
rect 12911 1492 13039 1520
rect 14236 1415 14338 1447
rect 11248 1381 12262 1387
rect 11248 1354 12144 1381
rect 12132 1347 12144 1354
rect 12178 1347 12216 1381
rect 12250 1347 12262 1381
rect 12132 1341 12262 1347
rect 10820 1330 10872 1336
rect 9612 1287 9670 1329
rect 4800 823 5019 1016
<< via1 >>
rect 2793 2679 2845 2731
rect 2892 2679 2944 2731
rect 2991 2679 3043 2731
rect 3089 2679 3141 2731
rect 3187 2679 3239 2731
rect 3285 2679 3337 2731
rect 3383 2679 3435 2731
rect 3481 2679 3533 2731
rect 2793 2591 2845 2643
rect 2892 2591 2944 2643
rect 2991 2591 3043 2643
rect 3089 2591 3141 2643
rect 3187 2591 3239 2643
rect 3285 2591 3337 2643
rect 3383 2591 3435 2643
rect 3481 2591 3533 2643
rect 2793 2503 2845 2555
rect 2892 2503 2944 2555
rect 2991 2503 3043 2555
rect 3089 2503 3141 2555
rect 3187 2503 3239 2555
rect 3285 2503 3337 2555
rect 3383 2503 3435 2555
rect 3481 2503 3533 2555
rect 3689 1985 3741 2037
rect 2864 1906 2916 1958
rect 2928 1906 2980 1958
rect 3128 1905 3180 1957
rect 3198 1905 3250 1957
rect 3267 1905 3319 1957
rect 3336 1905 3388 1957
rect 3689 1921 3741 1973
rect 3885 1906 3937 1958
rect 3949 1906 4001 1958
rect 3242 1814 3294 1866
rect 3306 1814 3358 1866
rect 4893 1880 4945 1932
rect 4957 1880 5009 1932
rect 10594 1821 10646 1873
rect 10658 1821 10710 1873
rect 10849 1821 10901 1873
rect 10913 1821 10965 1873
rect 10584 1668 10636 1720
rect 10648 1668 10700 1720
rect 2779 1578 2831 1630
rect 2864 1578 2916 1630
rect 2949 1578 3001 1630
rect 2779 1506 2831 1558
rect 2864 1506 2916 1558
rect 2949 1506 3001 1558
rect 7691 1591 7743 1643
rect 7755 1591 7807 1643
rect 4455 1500 4507 1552
rect 4525 1500 4577 1552
rect 4595 1500 4647 1552
rect 4665 1500 4717 1552
rect 4735 1500 4787 1552
rect 4805 1500 4857 1552
rect 4875 1500 4927 1552
rect 4944 1500 4996 1552
rect 10820 1587 10872 1639
rect 10884 1587 10936 1639
rect 10820 1400 10872 1452
rect 10820 1336 10872 1388
rect 11248 1785 11300 1837
rect 13416 1819 13468 1871
rect 13480 1819 13532 1871
rect 11248 1721 11300 1773
rect 13473 1734 13525 1786
rect 13537 1734 13589 1786
rect 13473 1654 13525 1706
rect 13537 1654 13589 1706
rect 14225 1574 14277 1626
rect 14289 1574 14341 1626
<< metal2 >>
rect 2779 2676 2788 2732
rect 2844 2731 2874 2732
rect 2930 2731 2960 2732
rect 3016 2731 3046 2732
rect 3102 2731 3131 2732
rect 3187 2731 3216 2732
rect 3272 2731 3301 2732
rect 3357 2731 3386 2732
rect 2845 2679 2874 2731
rect 2944 2679 2960 2731
rect 3043 2679 3046 2731
rect 3272 2679 3285 2731
rect 3357 2679 3383 2731
rect 2844 2676 2874 2679
rect 2930 2676 2960 2679
rect 3016 2676 3046 2679
rect 3102 2676 3131 2679
rect 3187 2676 3216 2679
rect 3272 2676 3301 2679
rect 3357 2676 3386 2679
rect 3442 2676 3471 2732
rect 3527 2731 3539 2732
rect 3533 2679 3539 2731
rect 3527 2676 3539 2679
rect 2779 2648 3539 2676
rect 2779 2592 2788 2648
rect 2844 2643 2874 2648
rect 2930 2643 2960 2648
rect 3016 2643 3046 2648
rect 3102 2643 3131 2648
rect 3187 2643 3216 2648
rect 3272 2643 3301 2648
rect 3357 2643 3386 2648
rect 2845 2592 2874 2643
rect 2944 2592 2960 2643
rect 3043 2592 3046 2643
rect 3272 2592 3285 2643
rect 3357 2592 3383 2643
rect 3442 2592 3471 2648
rect 3527 2643 3539 2648
rect 2779 2591 2793 2592
rect 2845 2591 2892 2592
rect 2944 2591 2991 2592
rect 3043 2591 3089 2592
rect 3141 2591 3187 2592
rect 3239 2591 3285 2592
rect 3337 2591 3383 2592
rect 3435 2591 3481 2592
rect 3533 2591 3539 2643
rect 2779 2564 3539 2591
rect 2779 2508 2788 2564
rect 2844 2555 2874 2564
rect 2930 2555 2960 2564
rect 3016 2555 3046 2564
rect 3102 2555 3131 2564
rect 3187 2555 3216 2564
rect 3272 2555 3301 2564
rect 3357 2555 3386 2564
rect 2845 2508 2874 2555
rect 2944 2508 2960 2555
rect 3043 2508 3046 2555
rect 3272 2508 3285 2555
rect 3357 2508 3383 2555
rect 3442 2508 3471 2564
rect 3527 2555 3539 2564
rect 2787 2503 2793 2508
rect 2845 2503 2892 2508
rect 2944 2503 2991 2508
rect 3043 2503 3089 2508
rect 3141 2503 3187 2508
rect 3239 2503 3285 2508
rect 3337 2503 3383 2508
rect 3435 2503 3481 2508
rect 3533 2503 3539 2555
rect 2787 2502 3539 2503
tri 3007 2041 3010 2044 se
rect 3010 2041 3518 2044
tri 3518 2041 3521 2044 sw
tri 2924 1958 3007 2041 se
rect 3007 2004 3521 2041
rect 3007 1958 3009 2004
rect 2858 1906 2864 1958
rect 2916 1906 2928 1958
rect 2980 1957 3009 1958
tri 3009 1957 3056 2004 nw
tri 3476 1959 3521 2004 ne
tri 3521 1959 3603 2041 sw
rect 3689 2040 4181 2073
tri 4181 2040 4214 2073 sw
rect 3689 2037 6615 2040
rect 3741 2031 6615 2037
tri 4165 1998 4198 2031 ne
rect 4198 2002 6615 2031
tri 6615 2002 6653 2040 sw
rect 4198 1998 6653 2002
rect 3689 1973 3741 1985
tri 3521 1957 3523 1959 ne
rect 3523 1957 3603 1959
rect 2980 1906 2986 1957
tri 2986 1934 3009 1957 nw
rect 3122 1905 3128 1957
rect 3180 1905 3198 1957
rect 3250 1905 3267 1957
rect 3319 1905 3336 1957
rect 3388 1906 3471 1957
tri 3471 1906 3522 1957 sw
tri 3523 1906 3574 1957 ne
rect 3574 1906 3603 1957
rect 3388 1905 3522 1906
rect 3236 1814 3242 1866
rect 3294 1814 3306 1866
rect 3358 1862 3434 1866
tri 3434 1862 3438 1866 sw
tri 3465 1862 3508 1905 ne
rect 3508 1873 3522 1905
tri 3522 1873 3555 1906 sw
tri 3574 1877 3603 1906 ne
tri 3603 1877 3685 1959 sw
rect 3689 1915 3741 1921
rect 3879 1906 3885 1958
rect 3937 1906 3949 1958
rect 4001 1906 4007 1958
tri 6599 1944 6653 1998 ne
tri 6653 1944 6711 2002 sw
rect 3508 1862 3555 1873
rect 3358 1814 3438 1862
tri 3412 1792 3434 1814 ne
rect 3434 1792 3438 1814
tri 3438 1792 3508 1862 sw
tri 3508 1818 3552 1862 ne
rect 3552 1825 3555 1862
tri 3555 1825 3603 1873 sw
tri 3603 1825 3655 1877 ne
rect 3655 1825 3685 1877
rect 3552 1818 3603 1825
tri 3552 1795 3575 1818 ne
rect 3575 1795 3603 1818
tri 3603 1795 3633 1825 sw
tri 3655 1795 3685 1825 ne
tri 3685 1795 3767 1877 sw
rect 3939 1816 3979 1906
rect 4887 1880 4893 1932
rect 4945 1880 4957 1932
rect 5009 1880 6572 1932
tri 6550 1858 6572 1880 ne
tri 6572 1873 6631 1932 sw
tri 6653 1902 6695 1944 ne
rect 6695 1902 11181 1944
rect 6572 1858 10594 1873
tri 3434 1718 3508 1792 ne
tri 3508 1788 3512 1792 sw
rect 3508 1760 3512 1788
tri 3512 1760 3540 1788 sw
tri 3575 1760 3610 1795 ne
rect 3610 1760 3633 1795
tri 3633 1760 3668 1795 sw
rect 3508 1718 3540 1760
tri 3540 1718 3582 1760 sw
rect 2767 1593 2776 1649
rect 2832 1593 2859 1649
rect 2915 1630 2941 1649
rect 2997 1630 3006 1649
tri 3508 1644 3582 1718 ne
tri 3582 1714 3586 1718 sw
rect 3582 1702 3586 1714
tri 3586 1702 3598 1714 sw
tri 3610 1702 3668 1760 ne
tri 3668 1743 3685 1760 sw
tri 3685 1743 3737 1795 ne
rect 3737 1743 3767 1795
rect 3668 1702 3685 1743
tri 3685 1702 3726 1743 sw
tri 3737 1713 3767 1743 ne
tri 3767 1713 3849 1795 sw
tri 3939 1776 3979 1816 ne
tri 3979 1793 4020 1834 sw
tri 6572 1833 6597 1858 ne
rect 6597 1833 10594 1858
rect 10588 1821 10594 1833
rect 10646 1821 10658 1873
rect 10710 1821 10716 1873
rect 10843 1821 10849 1873
rect 10901 1821 10913 1873
rect 10965 1843 11027 1873
tri 11027 1843 11057 1873 sw
tri 11091 1843 11150 1902 ne
rect 11150 1843 11181 1902
tri 11181 1843 11282 1944 sw
rect 13410 1859 13416 1871
tri 11898 1845 11912 1859 se
rect 11912 1845 13416 1859
rect 10965 1821 11057 1843
rect 3979 1776 10991 1793
tri 3979 1753 4002 1776 ne
rect 4002 1765 10991 1776
tri 10991 1765 11019 1793 sw
tri 11021 1787 11055 1821 ne
rect 11055 1787 11057 1821
tri 11057 1787 11113 1843 sw
tri 11150 1787 11206 1843 ne
rect 11206 1837 11300 1843
rect 11206 1787 11248 1837
rect 4002 1753 11019 1765
rect 3582 1644 3598 1702
tri 3598 1644 3656 1702 sw
tri 3668 1644 3726 1702 ne
tri 3726 1673 3755 1702 sw
tri 3767 1673 3807 1713 ne
rect 3807 1673 10482 1713
rect 3726 1644 3755 1673
tri 3755 1644 3784 1673 sw
rect 2916 1593 2941 1630
rect 2767 1578 2779 1593
rect 2831 1578 2864 1593
rect 2916 1578 2949 1593
rect 3001 1578 3007 1630
rect 2767 1559 3007 1578
tri 3582 1570 3656 1644 ne
tri 3656 1577 3723 1644 sw
tri 3726 1602 3768 1644 ne
rect 3768 1635 6346 1644
tri 6346 1635 6355 1644 sw
rect 3768 1602 6355 1635
tri 6330 1577 6355 1602 ne
tri 6355 1577 6413 1635 sw
rect 7685 1591 7691 1643
rect 7743 1591 7755 1643
rect 7807 1633 7813 1643
tri 10448 1639 10482 1673 ne
tri 10482 1639 10556 1713 sw
rect 10578 1668 10584 1720
rect 10636 1668 10648 1720
rect 10700 1713 10706 1720
rect 10700 1709 10969 1713
tri 10969 1709 10973 1713 sw
tri 10973 1709 11017 1753 ne
rect 11017 1729 11019 1753
tri 11019 1729 11055 1765 sw
tri 11055 1729 11113 1787 ne
tri 11113 1729 11171 1787 sw
tri 11206 1781 11212 1787 ne
rect 11212 1785 11248 1787
tri 11854 1801 11898 1845 se
rect 11898 1819 13416 1845
rect 13468 1819 13480 1871
rect 13532 1819 13538 1871
rect 11898 1801 11912 1819
tri 11912 1801 11930 1819 nw
rect 11212 1781 11300 1785
rect 11248 1773 11300 1781
rect 11017 1709 11055 1729
rect 10700 1680 10973 1709
tri 10973 1680 11002 1709 sw
tri 11017 1680 11046 1709 ne
rect 11046 1707 11055 1709
tri 11055 1707 11077 1729 sw
rect 11046 1680 11077 1707
rect 10700 1673 11002 1680
rect 10700 1668 10706 1673
rect 7807 1598 10356 1633
tri 10356 1598 10391 1633 sw
rect 7807 1593 10391 1598
rect 7807 1591 7813 1593
rect 3656 1570 3723 1577
rect 2767 1503 2776 1559
rect 2832 1503 2859 1559
rect 2915 1558 2941 1559
rect 2997 1558 3007 1559
rect 2916 1506 2941 1558
rect 3001 1506 3007 1558
rect 2915 1503 2941 1506
rect 2997 1503 3006 1506
tri 3656 1503 3723 1570 ne
tri 3723 1552 3748 1577 sw
rect 3723 1503 4455 1552
tri 3723 1500 3726 1503 ne
rect 3726 1500 4455 1503
rect 4507 1500 4525 1552
rect 4577 1500 4595 1552
rect 4647 1500 4665 1552
rect 4717 1500 4735 1552
rect 4787 1500 4805 1552
rect 4857 1500 4875 1552
rect 4927 1500 4944 1552
rect 4996 1500 5002 1552
tri 6355 1519 6413 1577 ne
tri 6413 1519 6471 1577 sw
tri 10338 1540 10391 1593 ne
tri 10391 1540 10449 1598 sw
tri 10482 1587 10534 1639 ne
rect 10534 1587 10820 1639
rect 10872 1587 10884 1639
rect 10936 1587 10942 1639
tri 10952 1623 11002 1673 ne
tri 11002 1649 11033 1680 sw
tri 11046 1649 11077 1680 ne
tri 11077 1671 11113 1707 sw
tri 11113 1671 11171 1729 ne
tri 11171 1671 11229 1729 sw
tri 11796 1743 11854 1801 se
tri 11854 1743 11912 1801 nw
tri 11934 1765 11955 1786 se
rect 11955 1765 13473 1786
tri 11912 1743 11934 1765 se
rect 11934 1746 13473 1765
rect 11934 1743 11955 1746
rect 11248 1715 11300 1721
tri 11738 1685 11796 1743 se
tri 11796 1685 11854 1743 nw
tri 11897 1728 11912 1743 se
rect 11912 1728 11955 1743
tri 11955 1728 11973 1746 nw
rect 13467 1734 13473 1746
rect 13525 1734 13537 1786
rect 13589 1734 13595 1786
tri 11854 1685 11897 1728 se
rect 11077 1649 11113 1671
tri 11113 1649 11135 1671 sw
rect 11002 1623 11033 1649
tri 11033 1623 11059 1649 sw
tri 11002 1566 11059 1623 ne
tri 11059 1605 11077 1623 sw
tri 11077 1605 11121 1649 ne
rect 11121 1613 11135 1649
tri 11135 1613 11171 1649 sw
tri 11171 1613 11229 1671 ne
tri 11229 1613 11287 1671 sw
tri 11680 1627 11738 1685 se
tri 11738 1627 11796 1685 nw
tri 11839 1670 11854 1685 se
rect 11854 1670 11897 1685
tri 11897 1670 11955 1728 nw
tri 11965 1680 11991 1706 se
rect 11991 1680 13473 1706
tri 11955 1670 11965 1680 se
rect 11965 1670 13473 1680
tri 11796 1627 11839 1670 se
rect 11121 1605 11171 1613
rect 11059 1566 11077 1605
tri 11077 1566 11116 1605 sw
tri 11121 1566 11160 1605 ne
rect 11160 1591 11171 1605
tri 11171 1591 11193 1613 sw
rect 11160 1566 11193 1591
tri 6413 1461 6471 1519 ne
tri 6471 1461 6529 1519 sw
tri 10391 1500 10431 1540 ne
rect 10431 1509 11012 1540
tri 11012 1509 11043 1540 sw
tri 11059 1509 11116 1566 ne
tri 11116 1533 11149 1566 sw
tri 11160 1533 11193 1566 ne
tri 11193 1555 11229 1591 sw
tri 11229 1555 11287 1613 ne
tri 11287 1555 11345 1613 sw
tri 11622 1569 11680 1627 se
tri 11680 1569 11738 1627 nw
tri 11781 1612 11796 1627 se
rect 11796 1612 11839 1627
tri 11839 1612 11897 1670 nw
tri 11933 1648 11955 1670 se
rect 11955 1666 13473 1670
rect 11955 1648 11969 1666
tri 11897 1612 11933 1648 se
rect 11933 1626 11969 1648
tri 11969 1626 12009 1666 nw
tri 13316 1654 13328 1666 ne
rect 13328 1654 13473 1666
rect 13525 1654 13537 1706
rect 13589 1654 13595 1706
tri 11738 1569 11781 1612 se
tri 11608 1555 11622 1569 se
rect 11622 1555 11626 1569
rect 11193 1533 11229 1555
tri 11229 1533 11251 1555 sw
rect 11116 1509 11149 1533
tri 11149 1509 11173 1533 sw
rect 10431 1500 11043 1509
tri 6471 1419 6513 1461 ne
rect 6513 1447 10706 1461
tri 10706 1447 10720 1461 sw
rect 10820 1452 10872 1458
tri 10994 1452 11042 1500 ne
rect 11042 1452 11043 1500
tri 11043 1452 11100 1509 sw
tri 11116 1452 11173 1509 ne
tri 11173 1489 11193 1509 sw
tri 11193 1489 11237 1533 ne
rect 11237 1515 11251 1533
tri 11251 1515 11269 1533 sw
tri 11287 1515 11327 1555 ne
rect 11327 1515 11626 1555
tri 11626 1515 11680 1569 nw
tri 11723 1554 11738 1569 se
rect 11738 1554 11781 1569
tri 11781 1554 11839 1612 nw
tri 11875 1590 11897 1612 se
rect 11897 1590 11933 1612
tri 11933 1590 11969 1626 nw
tri 11999 1598 12027 1626 se
rect 12027 1598 14225 1626
tri 11839 1554 11875 1590 se
tri 11684 1515 11723 1554 se
rect 11237 1489 11269 1515
rect 11173 1452 11193 1489
tri 11193 1452 11230 1489 sw
tri 11237 1474 11252 1489 ne
rect 11252 1475 11269 1489
tri 11269 1475 11309 1515 sw
tri 11644 1475 11684 1515 se
rect 11684 1496 11723 1515
tri 11723 1496 11781 1554 nw
tri 11817 1532 11839 1554 se
rect 11839 1532 11875 1554
tri 11875 1532 11933 1590 nw
tri 11969 1568 11999 1598 se
rect 11999 1586 14225 1598
rect 11999 1568 12027 1586
tri 12027 1568 12045 1586 nw
rect 14219 1574 14225 1586
rect 14277 1574 14289 1626
rect 14341 1574 14347 1626
tri 11933 1532 11969 1568 se
tri 11781 1496 11817 1532 se
rect 11684 1475 11701 1496
rect 11252 1474 11701 1475
tri 11701 1474 11723 1496 nw
tri 11759 1474 11781 1496 se
rect 11781 1474 11817 1496
tri 11817 1474 11875 1532 nw
tri 11911 1510 11933 1532 se
rect 11933 1510 11969 1532
tri 11969 1510 12027 1568 nw
tri 11875 1474 11911 1510 se
rect 6513 1419 10820 1447
tri 10690 1400 10709 1419 ne
rect 10709 1400 10820 1419
rect 10820 1388 10872 1400
tri 11042 1395 11099 1452 ne
rect 11099 1395 11100 1452
tri 11100 1395 11157 1452 sw
tri 11173 1395 11230 1452 ne
tri 11230 1435 11247 1452 sw
tri 11252 1435 11291 1474 ne
rect 11291 1435 11662 1474
tri 11662 1435 11701 1474 nw
tri 11720 1435 11759 1474 se
rect 11230 1395 11247 1435
tri 11247 1395 11287 1435 sw
tri 11680 1395 11720 1435 se
rect 11720 1416 11759 1435
tri 11759 1416 11817 1474 nw
tri 11853 1452 11875 1474 se
rect 11875 1452 11911 1474
tri 11911 1452 11969 1510 nw
tri 11817 1416 11853 1452 se
rect 11720 1395 11738 1416
tri 11738 1395 11759 1416 nw
tri 11099 1355 11139 1395 ne
rect 11139 1355 11157 1395
tri 11157 1355 11197 1395 sw
tri 11230 1355 11270 1395 ne
rect 11270 1355 11698 1395
tri 11698 1355 11738 1395 nw
tri 11795 1394 11817 1416 se
rect 11817 1394 11853 1416
tri 11853 1394 11911 1452 nw
tri 11756 1355 11795 1394 se
rect 10820 1330 10872 1336
tri 11139 1315 11179 1355 ne
rect 11179 1315 11197 1355
tri 11197 1315 11237 1355 sw
tri 11716 1315 11756 1355 se
rect 11756 1336 11795 1355
tri 11795 1336 11853 1394 nw
rect 11756 1315 11774 1336
tri 11774 1315 11795 1336 nw
tri 11179 1275 11219 1315 ne
rect 11219 1275 11734 1315
tri 11734 1275 11774 1315 nw
<< via2 >>
rect 2788 2731 2844 2732
rect 2874 2731 2930 2732
rect 2960 2731 3016 2732
rect 3046 2731 3102 2732
rect 3131 2731 3187 2732
rect 3216 2731 3272 2732
rect 3301 2731 3357 2732
rect 3386 2731 3442 2732
rect 2788 2679 2793 2731
rect 2793 2679 2844 2731
rect 2874 2679 2892 2731
rect 2892 2679 2930 2731
rect 2960 2679 2991 2731
rect 2991 2679 3016 2731
rect 3046 2679 3089 2731
rect 3089 2679 3102 2731
rect 3131 2679 3141 2731
rect 3141 2679 3187 2731
rect 3216 2679 3239 2731
rect 3239 2679 3272 2731
rect 3301 2679 3337 2731
rect 3337 2679 3357 2731
rect 3386 2679 3435 2731
rect 3435 2679 3442 2731
rect 2788 2676 2844 2679
rect 2874 2676 2930 2679
rect 2960 2676 3016 2679
rect 3046 2676 3102 2679
rect 3131 2676 3187 2679
rect 3216 2676 3272 2679
rect 3301 2676 3357 2679
rect 3386 2676 3442 2679
rect 3471 2731 3527 2732
rect 3471 2679 3481 2731
rect 3481 2679 3527 2731
rect 3471 2676 3527 2679
rect 2788 2643 2844 2648
rect 2874 2643 2930 2648
rect 2960 2643 3016 2648
rect 3046 2643 3102 2648
rect 3131 2643 3187 2648
rect 3216 2643 3272 2648
rect 3301 2643 3357 2648
rect 3386 2643 3442 2648
rect 2788 2592 2793 2643
rect 2793 2592 2844 2643
rect 2874 2592 2892 2643
rect 2892 2592 2930 2643
rect 2960 2592 2991 2643
rect 2991 2592 3016 2643
rect 3046 2592 3089 2643
rect 3089 2592 3102 2643
rect 3131 2592 3141 2643
rect 3141 2592 3187 2643
rect 3216 2592 3239 2643
rect 3239 2592 3272 2643
rect 3301 2592 3337 2643
rect 3337 2592 3357 2643
rect 3386 2592 3435 2643
rect 3435 2592 3442 2643
rect 3471 2643 3527 2648
rect 3471 2592 3481 2643
rect 3481 2592 3527 2643
rect 2788 2555 2844 2564
rect 2874 2555 2930 2564
rect 2960 2555 3016 2564
rect 3046 2555 3102 2564
rect 3131 2555 3187 2564
rect 3216 2555 3272 2564
rect 3301 2555 3357 2564
rect 3386 2555 3442 2564
rect 2788 2508 2793 2555
rect 2793 2508 2844 2555
rect 2874 2508 2892 2555
rect 2892 2508 2930 2555
rect 2960 2508 2991 2555
rect 2991 2508 3016 2555
rect 3046 2508 3089 2555
rect 3089 2508 3102 2555
rect 3131 2508 3141 2555
rect 3141 2508 3187 2555
rect 3216 2508 3239 2555
rect 3239 2508 3272 2555
rect 3301 2508 3337 2555
rect 3337 2508 3357 2555
rect 3386 2508 3435 2555
rect 3435 2508 3442 2555
rect 3471 2555 3527 2564
rect 3471 2508 3481 2555
rect 3481 2508 3527 2555
rect 2776 1630 2832 1649
rect 2776 1593 2779 1630
rect 2779 1593 2831 1630
rect 2831 1593 2832 1630
rect 2859 1630 2915 1649
rect 2941 1630 2997 1649
rect 2859 1593 2864 1630
rect 2864 1593 2915 1630
rect 2941 1593 2949 1630
rect 2949 1593 2997 1630
rect 2776 1558 2832 1559
rect 2776 1506 2779 1558
rect 2779 1506 2831 1558
rect 2831 1506 2832 1558
rect 2776 1503 2832 1506
rect 2859 1558 2915 1559
rect 2941 1558 2997 1559
rect 2859 1506 2864 1558
rect 2864 1506 2915 1558
rect 2941 1506 2949 1558
rect 2949 1506 2997 1558
rect 2859 1503 2915 1506
rect 2941 1503 2997 1506
<< metal3 >>
tri 2771 2761 3000 2990 se
rect 3000 2761 3545 2895
rect 2771 2732 3545 2761
rect 2771 2676 2788 2732
rect 2844 2676 2874 2732
rect 2930 2676 2960 2732
rect 3016 2676 3046 2732
rect 3102 2676 3131 2732
rect 3187 2676 3216 2732
rect 3272 2676 3301 2732
rect 3357 2676 3386 2732
rect 3442 2676 3471 2732
rect 3527 2676 3545 2732
rect 2771 2648 3545 2676
rect 2771 2592 2788 2648
rect 2844 2592 2874 2648
rect 2930 2592 2960 2648
rect 3016 2592 3046 2648
rect 3102 2592 3131 2648
rect 3187 2592 3216 2648
rect 3272 2592 3301 2648
rect 3357 2592 3386 2648
rect 3442 2592 3471 2648
rect 3527 2592 3545 2648
rect 2771 2564 3545 2592
rect 2771 2508 2788 2564
rect 2844 2508 2874 2564
rect 2930 2508 2960 2564
rect 3016 2508 3046 2564
rect 3102 2508 3131 2564
rect 3187 2508 3216 2564
rect 3272 2508 3301 2564
rect 3357 2508 3386 2564
rect 3442 2508 3471 2564
rect 3527 2508 3545 2564
rect 2771 2497 3545 2508
rect 2771 1649 3009 2497
tri 3009 2400 3106 2497 nw
rect 2771 1593 2776 1649
rect 2832 1593 2859 1649
rect 2915 1593 2941 1649
rect 2997 1593 3009 1649
rect 2771 1559 3009 1593
rect 2771 1503 2776 1559
rect 2832 1503 2859 1559
rect 2915 1503 2941 1559
rect 2997 1503 3009 1559
rect 2771 1498 3009 1503
use sky130_fd_io__gpio_ovtv2_hotswap_latch_i2c_fix  sky130_fd_io__gpio_ovtv2_hotswap_latch_i2c_fix_0
timestamp 1676037725
transform 1 0 -9399 0 1 -970
box 11695 1627 37770 16163
use sky130_fd_io__sio_hotswap_log_ovtv2_i2c_fix  sky130_fd_io__sio_hotswap_log_ovtv2_i2c_fix_0
timestamp 1676037725
transform 1 0 8920 0 1 1484
box 16 -95 6374 1336
<< labels >>
flabel metal1 s 12939 1513 12978 1541 0 FreeSans 200 0 0 0 EN_H
port 1 nsew
flabel metal1 s 12679 1475 12721 1503 0 FreeSans 200 0 0 0 FORCEHI_H[1]
port 2 nsew
flabel metal1 s 14236 1415 14338 1447 0 FreeSans 200 0 0 0 OD_I_H_N
port 3 nsew
flabel metal1 s 8613 1547 8663 1593 3 FreeSans 520 0 0 0 ENHS_LAT_H_N
port 4 nsew
flabel metal1 s 3224 2201 3334 2247 3 FreeSans 520 0 0 0 PGHS_H
port 5 nsew
flabel metal1 s 12400 1972 12429 2248 0 FreeSans 200 0 0 0 VDDIO
port 6 nsew
flabel metal1 s 14371 1972 14400 2248 0 FreeSans 200 0 0 0 VDDIO
port 6 nsew
flabel metal1 s 11555 1972 11581 2248 0 FreeSans 200 0 0 0 VDDIO
port 6 nsew
flabel metal1 s 14371 2498 14400 2700 0 FreeSans 200 0 0 0 VSSD
port 7 nsew
flabel metal1 s 12400 2498 12429 2700 0 FreeSans 200 0 0 0 VSSD
port 7 nsew
flabel metal1 s 14371 2424 14400 2470 0 FreeSans 200 0 0 0 VSSD
port 7 nsew
flabel metal1 s 12400 2424 12429 2470 0 FreeSans 200 0 0 0 VSSD
port 7 nsew
flabel metal1 s 11522 2424 11542 2470 0 FreeSans 200 0 0 0 VSSD
port 7 nsew
flabel metal1 s 11522 2498 11542 2700 0 FreeSans 200 0 0 0 VSSD
port 7 nsew
flabel metal1 s 12429 2424 12458 2470 0 FreeSans 200 0 0 0 VSSD
port 7 nsew
flabel metal1 s 12429 2498 12458 2700 0 FreeSans 200 0 0 0 VSSD
port 7 nsew
flabel metal1 s 4800 823 5019 1016 3 FreeSans 520 0 0 0 VDDIO
port 6 nsew
flabel metal1 s 5273 2579 5506 2710 3 FreeSans 520 0 0 0 VSSD
port 7 nsew
flabel metal1 s 3061 1511 3294 1626 3 FreeSans 520 0 0 0 VSSD
port 7 nsew
flabel metal1 s 9612 1287 9670 1329 0 FreeSans 440 0 0 0 VPWR_KA
port 8 nsew
flabel metal1 s 5354 1505 5412 1547 0 FreeSans 440 180 0 0 PAD_ESD
port 9 nsew
<< properties >>
string GDS_END 34148584
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 34133488
<< end >>
