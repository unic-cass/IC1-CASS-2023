magic
tech sky130B
magscale 1 2
timestamp 1676037725
use sky130_fd_pr__dfl1sd2__example_55959141808104  sky130_fd_pr__dfl1sd2__example_55959141808104_0
timestamp 1676037725
transform -1 0 -32 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808104  sky130_fd_pr__dfl1sd2__example_55959141808104_1
timestamp 1676037725
transform 1 0 100 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 33978302
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 33977184
<< end >>
