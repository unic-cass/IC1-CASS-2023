magic
tech sky130B
magscale 1 2
timestamp 1676037725
<< pwell >>
rect 1176 3561 1197 3610
rect 3392 3561 3413 3610
rect 1176 1289 1197 1338
rect 3392 1289 3413 1338
rect 1179 1269 1189 1279
<< obsli1 >>
rect 0 0 4498 4610
<< obsm1 >>
rect 0 4544 4498 4610
rect 0 2338 72 4544
rect 100 3473 128 4516
rect 156 3501 184 4544
rect 212 3473 240 4516
rect 268 3501 296 4544
rect 324 3473 352 4516
rect 380 3501 408 4544
rect 436 3473 464 4516
rect 492 3501 520 4544
rect 548 3473 576 4516
rect 604 3501 632 4544
rect 660 3473 688 4516
rect 716 3501 744 4544
rect 772 3473 800 4516
rect 828 3501 856 4544
rect 884 3473 912 4516
rect 940 3501 968 4544
rect 996 3473 1024 4516
rect 1052 3501 1080 4544
rect 1108 3473 1174 4516
rect 1202 3501 1230 4544
rect 1258 3473 1286 4516
rect 1314 3501 1342 4544
rect 1370 3473 1398 4516
rect 1426 3501 1454 4544
rect 1482 3473 1510 4516
rect 1538 3501 1566 4544
rect 1594 3473 1622 4516
rect 1650 3501 1678 4544
rect 1706 3473 1734 4516
rect 1762 3501 1790 4544
rect 1818 3473 1846 4516
rect 1874 3501 1902 4544
rect 1930 3473 1958 4516
rect 1986 3501 2014 4544
rect 2042 3473 2070 4516
rect 2098 3501 2126 4544
rect 2154 3473 2182 4516
rect 100 3409 2182 3473
rect 100 2366 128 3409
rect 156 2338 184 3381
rect 212 2366 240 3409
rect 268 2338 296 3381
rect 324 2366 352 3409
rect 380 2338 408 3381
rect 436 2366 464 3409
rect 492 2338 520 3381
rect 548 2366 576 3409
rect 604 2338 632 3381
rect 660 2366 688 3409
rect 716 2338 744 3381
rect 772 2366 800 3409
rect 828 2338 856 3381
rect 884 2366 912 3409
rect 940 2338 968 3381
rect 996 2366 1024 3409
rect 1052 2338 1080 3381
rect 1108 2366 1174 3409
rect 1202 2338 1230 3381
rect 1258 2366 1286 3409
rect 1314 2338 1342 3381
rect 1370 2366 1398 3409
rect 1426 2338 1454 3381
rect 1482 2366 1510 3409
rect 1538 2338 1566 3381
rect 1594 2366 1622 3409
rect 1650 2338 1678 3381
rect 1706 2366 1734 3409
rect 1762 2338 1790 3381
rect 1818 2366 1846 3409
rect 1874 2338 1902 3381
rect 1930 2366 1958 3409
rect 1986 2338 2014 3381
rect 2042 2366 2070 3409
rect 2098 2338 2126 3381
rect 2154 2366 2182 3409
rect 2210 2338 2288 4544
rect 2316 3473 2344 4516
rect 2372 3501 2400 4544
rect 2428 3473 2456 4516
rect 2484 3501 2512 4544
rect 2540 3473 2568 4516
rect 2596 3501 2624 4544
rect 2652 3473 2680 4516
rect 2708 3501 2736 4544
rect 2764 3473 2792 4516
rect 2820 3501 2848 4544
rect 2876 3473 2904 4516
rect 2932 3501 2960 4544
rect 2988 3473 3016 4516
rect 3044 3501 3072 4544
rect 3100 3473 3128 4516
rect 3156 3501 3184 4544
rect 3212 3473 3240 4516
rect 3268 3501 3296 4544
rect 3324 3473 3390 4516
rect 3418 3501 3446 4544
rect 3474 3473 3502 4516
rect 3530 3501 3558 4544
rect 3586 3473 3614 4516
rect 3642 3501 3670 4544
rect 3698 3473 3726 4516
rect 3754 3501 3782 4544
rect 3810 3473 3838 4516
rect 3866 3501 3894 4544
rect 3922 3473 3950 4516
rect 3978 3501 4006 4544
rect 4034 3473 4062 4516
rect 4090 3501 4118 4544
rect 4146 3473 4174 4516
rect 4202 3501 4230 4544
rect 4258 3473 4286 4516
rect 4314 3501 4342 4544
rect 4370 3473 4398 4516
rect 2316 3409 4398 3473
rect 2316 2366 2344 3409
rect 2372 2338 2400 3381
rect 2428 2366 2456 3409
rect 2484 2338 2512 3381
rect 2540 2366 2568 3409
rect 2596 2338 2624 3381
rect 2652 2366 2680 3409
rect 2708 2338 2736 3381
rect 2764 2366 2792 3409
rect 2820 2338 2848 3381
rect 2876 2366 2904 3409
rect 2932 2338 2960 3381
rect 2988 2366 3016 3409
rect 3044 2338 3072 3381
rect 3100 2366 3128 3409
rect 3156 2338 3184 3381
rect 3212 2366 3240 3409
rect 3268 2338 3296 3381
rect 3324 2366 3390 3409
rect 3418 2338 3446 3381
rect 3474 2366 3502 3409
rect 3530 2338 3558 3381
rect 3586 2366 3614 3409
rect 3642 2338 3670 3381
rect 3698 2366 3726 3409
rect 3754 2338 3782 3381
rect 3810 2366 3838 3409
rect 3866 2338 3894 3381
rect 3922 2366 3950 3409
rect 3978 2338 4006 3381
rect 4034 2366 4062 3409
rect 4090 2338 4118 3381
rect 4146 2366 4174 3409
rect 4202 2338 4230 3381
rect 4258 2366 4286 3409
rect 4314 2338 4342 3381
rect 4370 2366 4398 3409
rect 4426 2338 4498 4544
rect 0 2272 4498 2338
rect 0 66 72 2272
rect 100 1201 128 2244
rect 156 1229 184 2272
rect 212 1201 240 2244
rect 268 1229 296 2272
rect 324 1201 352 2244
rect 380 1229 408 2272
rect 436 1201 464 2244
rect 492 1229 520 2272
rect 548 1201 576 2244
rect 604 1229 632 2272
rect 660 1201 688 2244
rect 716 1229 744 2272
rect 772 1201 800 2244
rect 828 1229 856 2272
rect 884 1201 912 2244
rect 940 1229 968 2272
rect 996 1201 1024 2244
rect 1052 1229 1080 2272
rect 1108 1201 1174 2244
rect 1202 1229 1230 2272
rect 1258 1201 1286 2244
rect 1314 1229 1342 2272
rect 1370 1201 1398 2244
rect 1426 1229 1454 2272
rect 1482 1201 1510 2244
rect 1538 1229 1566 2272
rect 1594 1201 1622 2244
rect 1650 1229 1678 2272
rect 1706 1201 1734 2244
rect 1762 1229 1790 2272
rect 1818 1201 1846 2244
rect 1874 1229 1902 2272
rect 1930 1201 1958 2244
rect 1986 1229 2014 2272
rect 2042 1201 2070 2244
rect 2098 1229 2126 2272
rect 2154 1201 2182 2244
rect 100 1137 2182 1201
rect 100 94 128 1137
rect 156 66 184 1109
rect 212 94 240 1137
rect 268 66 296 1109
rect 324 94 352 1137
rect 380 66 408 1109
rect 436 94 464 1137
rect 492 66 520 1109
rect 548 94 576 1137
rect 604 66 632 1109
rect 660 94 688 1137
rect 716 66 744 1109
rect 772 94 800 1137
rect 828 66 856 1109
rect 884 94 912 1137
rect 940 66 968 1109
rect 996 94 1024 1137
rect 1052 66 1080 1109
rect 1108 94 1174 1137
rect 1202 66 1230 1109
rect 1258 94 1286 1137
rect 1314 66 1342 1109
rect 1370 94 1398 1137
rect 1426 66 1454 1109
rect 1482 94 1510 1137
rect 1538 66 1566 1109
rect 1594 94 1622 1137
rect 1650 66 1678 1109
rect 1706 94 1734 1137
rect 1762 66 1790 1109
rect 1818 94 1846 1137
rect 1874 66 1902 1109
rect 1930 94 1958 1137
rect 1986 66 2014 1109
rect 2042 94 2070 1137
rect 2098 66 2126 1109
rect 2154 94 2182 1137
rect 2210 66 2288 2272
rect 2316 1201 2344 2244
rect 2372 1229 2400 2272
rect 2428 1201 2456 2244
rect 2484 1229 2512 2272
rect 2540 1201 2568 2244
rect 2596 1229 2624 2272
rect 2652 1201 2680 2244
rect 2708 1229 2736 2272
rect 2764 1201 2792 2244
rect 2820 1229 2848 2272
rect 2876 1201 2904 2244
rect 2932 1229 2960 2272
rect 2988 1201 3016 2244
rect 3044 1229 3072 2272
rect 3100 1201 3128 2244
rect 3156 1229 3184 2272
rect 3212 1201 3240 2244
rect 3268 1229 3296 2272
rect 3324 1201 3390 2244
rect 3418 1229 3446 2272
rect 3474 1201 3502 2244
rect 3530 1229 3558 2272
rect 3586 1201 3614 2244
rect 3642 1229 3670 2272
rect 3698 1201 3726 2244
rect 3754 1229 3782 2272
rect 3810 1201 3838 2244
rect 3866 1229 3894 2272
rect 3922 1201 3950 2244
rect 3978 1229 4006 2272
rect 4034 1201 4062 2244
rect 4090 1229 4118 2272
rect 4146 1201 4174 2244
rect 4202 1229 4230 2272
rect 4258 1201 4286 2244
rect 4314 1229 4342 2272
rect 4370 1201 4398 2244
rect 2316 1137 4398 1201
rect 2316 94 2344 1137
rect 2372 66 2400 1109
rect 2428 94 2456 1137
rect 2484 66 2512 1109
rect 2540 94 2568 1137
rect 2596 66 2624 1109
rect 2652 94 2680 1137
rect 2708 66 2736 1109
rect 2764 94 2792 1137
rect 2820 66 2848 1109
rect 2876 94 2904 1137
rect 2932 66 2960 1109
rect 2988 94 3016 1137
rect 3044 66 3072 1109
rect 3100 94 3128 1137
rect 3156 66 3184 1109
rect 3212 94 3240 1137
rect 3268 66 3296 1109
rect 3324 94 3390 1137
rect 3418 66 3446 1109
rect 3474 94 3502 1137
rect 3530 66 3558 1109
rect 3586 94 3614 1137
rect 3642 66 3670 1109
rect 3698 94 3726 1137
rect 3754 66 3782 1109
rect 3810 94 3838 1137
rect 3866 66 3894 1109
rect 3922 94 3950 1137
rect 3978 66 4006 1109
rect 4034 94 4062 1137
rect 4090 66 4118 1109
rect 4146 94 4174 1137
rect 4202 66 4230 1109
rect 4258 94 4286 1137
rect 4314 66 4342 1109
rect 4370 94 4398 1137
rect 4426 66 4498 2272
rect 0 0 4498 66
<< obsm2 >>
rect 0 4544 1086 4610
rect 0 4460 66 4544
rect 1114 4516 1168 4610
rect 1196 4544 3302 4610
rect 94 4488 2188 4516
rect 0 4432 1085 4460
rect 0 4348 66 4432
rect 1113 4404 1169 4488
rect 2216 4460 2282 4544
rect 3330 4516 3384 4610
rect 3412 4544 4498 4610
rect 2310 4488 4404 4516
rect 1197 4432 3301 4460
rect 94 4376 2188 4404
rect 0 4320 1085 4348
rect 0 4236 66 4320
rect 1113 4292 1169 4376
rect 2216 4348 2282 4432
rect 3329 4404 3385 4488
rect 4432 4460 4498 4544
rect 3413 4432 4498 4460
rect 2310 4376 4404 4404
rect 1197 4320 3301 4348
rect 94 4264 2188 4292
rect 0 4208 1085 4236
rect 0 4124 66 4208
rect 1113 4180 1169 4264
rect 2216 4236 2282 4320
rect 3329 4292 3385 4376
rect 4432 4348 4498 4432
rect 3413 4320 4498 4348
rect 2310 4264 4404 4292
rect 1197 4208 3301 4236
rect 94 4152 2188 4180
rect 0 4096 1085 4124
rect 0 4012 66 4096
rect 1113 4068 1169 4152
rect 2216 4124 2282 4208
rect 3329 4180 3385 4264
rect 4432 4236 4498 4320
rect 3413 4208 4498 4236
rect 2310 4152 4404 4180
rect 1197 4096 3301 4124
rect 94 4040 2188 4068
rect 0 3984 1085 4012
rect 0 3900 66 3984
rect 1113 3956 1169 4040
rect 2216 4012 2282 4096
rect 3329 4068 3385 4152
rect 4432 4124 4498 4208
rect 3413 4096 4498 4124
rect 2310 4040 4404 4068
rect 1197 3984 3301 4012
rect 94 3928 2188 3956
rect 0 3872 1085 3900
rect 0 3788 66 3872
rect 1113 3844 1169 3928
rect 2216 3900 2282 3984
rect 3329 3956 3385 4040
rect 4432 4012 4498 4096
rect 3413 3984 4498 4012
rect 2310 3928 4404 3956
rect 1197 3872 3301 3900
rect 94 3816 2188 3844
rect 0 3760 1085 3788
rect 0 3676 66 3760
rect 1113 3732 1169 3816
rect 2216 3788 2282 3872
rect 3329 3844 3385 3928
rect 4432 3900 4498 3984
rect 3413 3872 4498 3900
rect 2310 3816 4404 3844
rect 1197 3760 3301 3788
rect 94 3704 2188 3732
rect 0 3648 1085 3676
rect 0 3564 66 3648
rect 1113 3620 1169 3704
rect 2216 3676 2282 3760
rect 3329 3732 3385 3816
rect 4432 3788 4498 3872
rect 3413 3760 4498 3788
rect 2310 3704 4404 3732
rect 1197 3648 3301 3676
rect 94 3592 2188 3620
rect 0 3497 1085 3564
rect 0 3496 66 3497
rect 1113 3469 1169 3592
rect 2216 3564 2282 3648
rect 3329 3620 3385 3704
rect 4432 3676 4498 3760
rect 3413 3648 4498 3676
rect 2310 3592 4404 3620
rect 1197 3497 3301 3564
rect 2216 3496 2282 3497
rect 3329 3469 3385 3592
rect 4432 3564 4498 3648
rect 3413 3497 4498 3564
rect 4432 3496 4498 3497
rect 74 3468 2208 3469
rect 2290 3468 4424 3469
rect 0 3414 4498 3468
rect 74 3413 2208 3414
rect 2290 3413 4424 3414
rect 0 3385 66 3386
rect 0 3318 1085 3385
rect 0 3234 66 3318
rect 1113 3290 1169 3413
rect 2216 3385 2282 3386
rect 1197 3318 3301 3385
rect 94 3262 2188 3290
rect 0 3206 1085 3234
rect 0 3122 66 3206
rect 1113 3178 1169 3262
rect 2216 3234 2282 3318
rect 3329 3290 3385 3413
rect 4432 3385 4498 3386
rect 3413 3318 4498 3385
rect 2310 3262 4404 3290
rect 1197 3206 3301 3234
rect 94 3150 2188 3178
rect 0 3094 1085 3122
rect 0 3010 66 3094
rect 1113 3066 1169 3150
rect 2216 3122 2282 3206
rect 3329 3178 3385 3262
rect 4432 3234 4498 3318
rect 3413 3206 4498 3234
rect 2310 3150 4404 3178
rect 1197 3094 3301 3122
rect 94 3038 2188 3066
rect 0 2982 1085 3010
rect 0 2898 66 2982
rect 1113 2954 1169 3038
rect 2216 3010 2282 3094
rect 3329 3066 3385 3150
rect 4432 3122 4498 3206
rect 3413 3094 4498 3122
rect 2310 3038 4404 3066
rect 1197 2982 3301 3010
rect 94 2926 2188 2954
rect 0 2870 1085 2898
rect 0 2786 66 2870
rect 1113 2842 1169 2926
rect 2216 2898 2282 2982
rect 3329 2954 3385 3038
rect 4432 3010 4498 3094
rect 3413 2982 4498 3010
rect 2310 2926 4404 2954
rect 1197 2870 3301 2898
rect 94 2814 2188 2842
rect 0 2758 1085 2786
rect 0 2674 66 2758
rect 1113 2730 1169 2814
rect 2216 2786 2282 2870
rect 3329 2842 3385 2926
rect 4432 2898 4498 2982
rect 3413 2870 4498 2898
rect 2310 2814 4404 2842
rect 1197 2758 3301 2786
rect 94 2702 2188 2730
rect 0 2646 1085 2674
rect 0 2562 66 2646
rect 1113 2618 1169 2702
rect 2216 2674 2282 2758
rect 3329 2730 3385 2814
rect 4432 2786 4498 2870
rect 3413 2758 4498 2786
rect 2310 2702 4404 2730
rect 1197 2646 3301 2674
rect 94 2590 2188 2618
rect 0 2534 1085 2562
rect 0 2450 66 2534
rect 1113 2506 1169 2590
rect 2216 2562 2282 2646
rect 3329 2618 3385 2702
rect 4432 2674 4498 2758
rect 3413 2646 4498 2674
rect 2310 2590 4404 2618
rect 1197 2534 3301 2562
rect 94 2478 2188 2506
rect 0 2422 1085 2450
rect 0 2338 66 2422
rect 1113 2394 1169 2478
rect 2216 2450 2282 2534
rect 3329 2506 3385 2590
rect 4432 2562 4498 2646
rect 3413 2534 4498 2562
rect 2310 2478 4404 2506
rect 1197 2422 3301 2450
rect 94 2366 2188 2394
rect 0 2272 1086 2338
rect 0 2188 66 2272
rect 1114 2244 1168 2366
rect 2216 2338 2282 2422
rect 3329 2394 3385 2478
rect 4432 2450 4498 2534
rect 3413 2422 4498 2450
rect 2310 2366 4404 2394
rect 1196 2272 3302 2338
rect 94 2216 2188 2244
rect 0 2160 1085 2188
rect 0 2076 66 2160
rect 1113 2132 1169 2216
rect 2216 2188 2282 2272
rect 3330 2244 3384 2366
rect 4432 2338 4498 2422
rect 3412 2272 4498 2338
rect 2310 2216 4404 2244
rect 1197 2160 3301 2188
rect 94 2104 2188 2132
rect 0 2048 1085 2076
rect 0 1964 66 2048
rect 1113 2020 1169 2104
rect 2216 2076 2282 2160
rect 3329 2132 3385 2216
rect 4432 2188 4498 2272
rect 3413 2160 4498 2188
rect 2310 2104 4404 2132
rect 1197 2048 3301 2076
rect 94 1992 2188 2020
rect 0 1936 1085 1964
rect 0 1852 66 1936
rect 1113 1908 1169 1992
rect 2216 1964 2282 2048
rect 3329 2020 3385 2104
rect 4432 2076 4498 2160
rect 3413 2048 4498 2076
rect 2310 1992 4404 2020
rect 1197 1936 3301 1964
rect 94 1880 2188 1908
rect 0 1824 1085 1852
rect 0 1740 66 1824
rect 1113 1796 1169 1880
rect 2216 1852 2282 1936
rect 3329 1908 3385 1992
rect 4432 1964 4498 2048
rect 3413 1936 4498 1964
rect 2310 1880 4404 1908
rect 1197 1824 3301 1852
rect 94 1768 2188 1796
rect 0 1712 1085 1740
rect 0 1628 66 1712
rect 1113 1684 1169 1768
rect 2216 1740 2282 1824
rect 3329 1796 3385 1880
rect 4432 1852 4498 1936
rect 3413 1824 4498 1852
rect 2310 1768 4404 1796
rect 1197 1712 3301 1740
rect 94 1656 2188 1684
rect 0 1600 1085 1628
rect 0 1516 66 1600
rect 1113 1572 1169 1656
rect 2216 1628 2282 1712
rect 3329 1684 3385 1768
rect 4432 1740 4498 1824
rect 3413 1712 4498 1740
rect 2310 1656 4404 1684
rect 1197 1600 3301 1628
rect 94 1544 2188 1572
rect 0 1488 1085 1516
rect 0 1404 66 1488
rect 1113 1460 1169 1544
rect 2216 1516 2282 1600
rect 3329 1572 3385 1656
rect 4432 1628 4498 1712
rect 3413 1600 4498 1628
rect 2310 1544 4404 1572
rect 1197 1488 3301 1516
rect 94 1432 2188 1460
rect 0 1376 1085 1404
rect 0 1292 66 1376
rect 1113 1348 1169 1432
rect 2216 1404 2282 1488
rect 3329 1460 3385 1544
rect 4432 1516 4498 1600
rect 3413 1488 4498 1516
rect 2310 1432 4404 1460
rect 1197 1376 3301 1404
rect 94 1320 2188 1348
rect 0 1225 1085 1292
rect 0 1224 66 1225
rect 1113 1197 1169 1320
rect 2216 1292 2282 1376
rect 3329 1348 3385 1432
rect 4432 1404 4498 1488
rect 3413 1376 4498 1404
rect 2310 1320 4404 1348
rect 1197 1225 3301 1292
rect 2216 1224 2282 1225
rect 3329 1197 3385 1320
rect 4432 1292 4498 1376
rect 3413 1225 4498 1292
rect 4432 1224 4498 1225
rect 74 1196 2208 1197
rect 2290 1196 4424 1197
rect 0 1142 4498 1196
rect 74 1141 2208 1142
rect 2290 1141 4424 1142
rect 0 1113 66 1114
rect 0 1046 1085 1113
rect 0 962 66 1046
rect 1113 1018 1169 1141
rect 2216 1113 2282 1114
rect 1197 1046 3301 1113
rect 94 990 2188 1018
rect 0 934 1085 962
rect 0 850 66 934
rect 1113 906 1169 990
rect 2216 962 2282 1046
rect 3329 1018 3385 1141
rect 4432 1113 4498 1114
rect 3413 1046 4498 1113
rect 2310 990 4404 1018
rect 1197 934 3301 962
rect 94 878 2188 906
rect 0 822 1085 850
rect 0 738 66 822
rect 1113 794 1169 878
rect 2216 850 2282 934
rect 3329 906 3385 990
rect 4432 962 4498 1046
rect 3413 934 4498 962
rect 2310 878 4404 906
rect 1197 822 3301 850
rect 94 766 2188 794
rect 0 710 1085 738
rect 0 626 66 710
rect 1113 682 1169 766
rect 2216 738 2282 822
rect 3329 794 3385 878
rect 4432 850 4498 934
rect 3413 822 4498 850
rect 2310 766 4404 794
rect 1197 710 3301 738
rect 94 654 2188 682
rect 0 598 1085 626
rect 0 514 66 598
rect 1113 570 1169 654
rect 2216 626 2282 710
rect 3329 682 3385 766
rect 4432 738 4498 822
rect 3413 710 4498 738
rect 2310 654 4404 682
rect 1197 598 3301 626
rect 94 542 2188 570
rect 0 486 1085 514
rect 0 402 66 486
rect 1113 458 1169 542
rect 2216 514 2282 598
rect 3329 570 3385 654
rect 4432 626 4498 710
rect 3413 598 4498 626
rect 2310 542 4404 570
rect 1197 486 3301 514
rect 94 430 2188 458
rect 0 374 1085 402
rect 0 290 66 374
rect 1113 346 1169 430
rect 2216 402 2282 486
rect 3329 458 3385 542
rect 4432 514 4498 598
rect 3413 486 4498 514
rect 2310 430 4404 458
rect 1197 374 3301 402
rect 94 318 2188 346
rect 0 262 1085 290
rect 0 178 66 262
rect 1113 234 1169 318
rect 2216 290 2282 374
rect 3329 346 3385 430
rect 4432 402 4498 486
rect 3413 374 4498 402
rect 2310 318 4404 346
rect 1197 262 3301 290
rect 94 206 2188 234
rect 0 150 1085 178
rect 0 66 66 150
rect 1113 122 1169 206
rect 2216 178 2282 262
rect 3329 234 3385 318
rect 4432 290 4498 374
rect 3413 262 4498 290
rect 2310 206 4404 234
rect 1197 150 3301 178
rect 94 94 2188 122
rect 0 0 1086 66
rect 1114 0 1168 94
rect 2216 66 2282 150
rect 3329 122 3385 206
rect 4432 178 4498 262
rect 3413 150 4498 178
rect 2310 94 4404 122
rect 1196 0 3302 66
rect 3330 0 3384 94
rect 4432 66 4498 150
rect 3412 0 4498 66
<< obsm3 >>
rect 0 4544 4498 4610
rect 0 2338 66 4544
rect 126 3474 186 4484
rect 246 3534 306 4544
rect 366 3474 426 4484
rect 486 3534 546 4544
rect 606 3474 666 4484
rect 726 3534 786 4544
rect 846 3474 906 4484
rect 966 3534 1048 4544
rect 1108 3474 1174 4484
rect 1234 3534 1316 4544
rect 1376 3474 1436 4484
rect 1496 3534 1556 4544
rect 1616 3474 1676 4484
rect 1736 3534 1796 4544
rect 1856 3474 1916 4484
rect 1976 3534 2036 4544
rect 2096 3474 2156 4484
rect 126 3408 2156 3474
rect 126 2398 186 3408
rect 246 2338 306 3348
rect 366 2398 426 3408
rect 486 2338 546 3348
rect 606 2398 666 3408
rect 726 2338 786 3348
rect 846 2398 906 3408
rect 966 2338 1048 3348
rect 1108 2398 1174 3408
rect 1234 2338 1316 3348
rect 1376 2398 1436 3408
rect 1496 2338 1556 3348
rect 1616 2398 1676 3408
rect 1736 2338 1796 3348
rect 1856 2398 1916 3408
rect 1976 2338 2036 3348
rect 2096 2398 2156 3408
rect 2216 2338 2282 4544
rect 2342 3474 2402 4484
rect 2462 3534 2522 4544
rect 2582 3474 2642 4484
rect 2702 3534 2762 4544
rect 2822 3474 2882 4484
rect 2942 3534 3002 4544
rect 3062 3474 3122 4484
rect 3182 3534 3264 4544
rect 3324 3474 3390 4484
rect 3450 3534 3532 4544
rect 3592 3474 3652 4484
rect 3712 3534 3772 4544
rect 3832 3474 3892 4484
rect 3952 3534 4012 4544
rect 4072 3474 4132 4484
rect 4192 3534 4252 4544
rect 4312 3474 4372 4484
rect 2342 3408 4372 3474
rect 2342 2398 2402 3408
rect 2462 2338 2522 3348
rect 2582 2398 2642 3408
rect 2702 2338 2762 3348
rect 2822 2398 2882 3408
rect 2942 2338 3002 3348
rect 3062 2398 3122 3408
rect 3182 2338 3264 3348
rect 3324 2398 3390 3408
rect 3450 2338 3532 3348
rect 3592 2398 3652 3408
rect 3712 2338 3772 3348
rect 3832 2398 3892 3408
rect 3952 2338 4012 3348
rect 4072 2398 4132 3408
rect 4192 2338 4252 3348
rect 4312 2398 4372 3408
rect 4432 2338 4498 4544
rect 0 2272 4498 2338
rect 0 66 66 2272
rect 126 1202 186 2212
rect 246 1262 306 2272
rect 366 1202 426 2212
rect 486 1262 546 2272
rect 606 1202 666 2212
rect 726 1262 786 2272
rect 846 1202 906 2212
rect 966 1262 1048 2272
rect 1108 1202 1174 2212
rect 1234 1262 1316 2272
rect 1376 1202 1436 2212
rect 1496 1262 1556 2272
rect 1616 1202 1676 2212
rect 1736 1262 1796 2272
rect 1856 1202 1916 2212
rect 1976 1262 2036 2272
rect 2096 1202 2156 2212
rect 126 1136 2156 1202
rect 126 126 186 1136
rect 246 66 306 1076
rect 366 126 426 1136
rect 486 66 546 1076
rect 606 126 666 1136
rect 726 66 786 1076
rect 846 126 906 1136
rect 966 66 1048 1076
rect 1108 126 1174 1136
rect 1234 66 1316 1076
rect 1376 126 1436 1136
rect 1496 66 1556 1076
rect 1616 126 1676 1136
rect 1736 66 1796 1076
rect 1856 126 1916 1136
rect 1976 66 2036 1076
rect 2096 126 2156 1136
rect 2216 66 2282 2272
rect 2342 1202 2402 2212
rect 2462 1262 2522 2272
rect 2582 1202 2642 2212
rect 2702 1262 2762 2272
rect 2822 1202 2882 2212
rect 2942 1262 3002 2272
rect 3062 1202 3122 2212
rect 3182 1262 3264 2272
rect 3324 1202 3390 2212
rect 3450 1262 3532 2272
rect 3592 1202 3652 2212
rect 3712 1262 3772 2272
rect 3832 1202 3892 2212
rect 3952 1262 4012 2272
rect 4072 1202 4132 2212
rect 4192 1262 4252 2272
rect 4312 1202 4372 2212
rect 2342 1136 4372 1202
rect 2342 126 2402 1136
rect 2462 66 2522 1076
rect 2582 126 2642 1136
rect 2702 66 2762 1076
rect 2822 126 2882 1136
rect 2942 66 3002 1076
rect 3062 126 3122 1136
rect 3182 66 3264 1076
rect 3324 126 3390 1136
rect 3450 66 3532 1076
rect 3592 126 3652 1136
rect 3712 66 3772 1076
rect 3832 126 3892 1136
rect 3952 66 4012 1076
rect 4072 126 4132 1136
rect 4192 66 4252 1076
rect 4312 126 4372 1136
rect 4432 66 4498 2272
rect 0 0 4498 66
<< metal4 >>
rect 0 4544 4498 4610
rect 0 4364 66 4544
rect 126 4424 2156 4484
rect 0 4304 1048 4364
rect 0 4124 66 4304
rect 1108 4244 1174 4424
rect 2216 4364 2282 4544
rect 2342 4424 4372 4484
rect 1234 4304 3264 4364
rect 126 4184 2156 4244
rect 0 4064 1048 4124
rect 0 3884 66 4064
rect 1108 4004 1174 4184
rect 2216 4124 2282 4304
rect 3324 4244 3390 4424
rect 4432 4364 4498 4544
rect 3450 4304 4498 4364
rect 2342 4184 4372 4244
rect 1234 4064 3264 4124
rect 126 3944 2156 4004
rect 0 3804 1048 3884
rect 0 3624 66 3804
rect 1108 3744 1174 3944
rect 2216 3884 2282 4064
rect 3324 4004 3390 4184
rect 4432 4124 4498 4304
rect 3450 4064 4498 4124
rect 2342 3944 4372 4004
rect 1234 3804 3264 3884
rect 126 3684 2156 3744
rect 0 3534 1048 3624
rect 0 3348 66 3534
rect 1108 3474 1174 3684
rect 2216 3624 2282 3804
rect 3324 3744 3390 3944
rect 4432 3884 4498 4064
rect 3450 3804 4498 3884
rect 2342 3684 4372 3744
rect 1234 3534 3264 3624
rect 126 3408 2156 3474
rect 0 3258 1048 3348
rect 0 3078 66 3258
rect 1108 3198 1174 3408
rect 2216 3348 2282 3534
rect 3324 3474 3390 3684
rect 4432 3624 4498 3804
rect 3450 3534 4498 3624
rect 2342 3408 4372 3474
rect 1234 3258 3264 3348
rect 126 3138 2156 3198
rect 0 2998 1048 3078
rect 0 2818 66 2998
rect 1108 2938 1174 3138
rect 2216 3078 2282 3258
rect 3324 3198 3390 3408
rect 4432 3348 4498 3534
rect 3450 3258 4498 3348
rect 2342 3138 4372 3198
rect 1234 2998 3264 3078
rect 126 2878 2156 2938
rect 0 2758 1048 2818
rect 0 2578 66 2758
rect 1108 2698 1174 2878
rect 2216 2818 2282 2998
rect 3324 2938 3390 3138
rect 4432 3078 4498 3258
rect 3450 2998 4498 3078
rect 2342 2878 4372 2938
rect 1234 2758 3264 2818
rect 126 2638 2156 2698
rect 0 2518 1048 2578
rect 0 2338 66 2518
rect 1108 2458 1174 2638
rect 2216 2578 2282 2758
rect 3324 2698 3390 2878
rect 4432 2818 4498 2998
rect 3450 2758 4498 2818
rect 2342 2638 4372 2698
rect 1234 2518 3264 2578
rect 126 2398 2156 2458
rect 2216 2338 2282 2518
rect 3324 2458 3390 2638
rect 4432 2578 4498 2758
rect 3450 2518 4498 2578
rect 2342 2398 4372 2458
rect 4432 2338 4498 2518
rect 0 2272 4498 2338
rect 0 2092 66 2272
rect 126 2152 2156 2212
rect 0 2032 1048 2092
rect 0 1852 66 2032
rect 1108 1972 1174 2152
rect 2216 2092 2282 2272
rect 2342 2152 4372 2212
rect 1234 2032 3264 2092
rect 126 1912 2156 1972
rect 0 1792 1048 1852
rect 0 1612 66 1792
rect 1108 1732 1174 1912
rect 2216 1852 2282 2032
rect 3324 1972 3390 2152
rect 4432 2092 4498 2272
rect 3450 2032 4498 2092
rect 2342 1912 4372 1972
rect 1234 1792 3264 1852
rect 126 1672 2156 1732
rect 0 1532 1048 1612
rect 0 1352 66 1532
rect 1108 1472 1174 1672
rect 2216 1612 2282 1792
rect 3324 1732 3390 1912
rect 4432 1852 4498 2032
rect 3450 1792 4498 1852
rect 2342 1672 4372 1732
rect 1234 1532 3264 1612
rect 126 1412 2156 1472
rect 0 1262 1048 1352
rect 0 1076 66 1262
rect 1108 1202 1174 1412
rect 2216 1352 2282 1532
rect 3324 1472 3390 1672
rect 4432 1612 4498 1792
rect 3450 1532 4498 1612
rect 2342 1412 4372 1472
rect 1234 1262 3264 1352
rect 126 1136 2156 1202
rect 0 986 1048 1076
rect 0 806 66 986
rect 1108 926 1174 1136
rect 2216 1076 2282 1262
rect 3324 1202 3390 1412
rect 4432 1352 4498 1532
rect 3450 1262 4498 1352
rect 2342 1136 4372 1202
rect 1234 986 3264 1076
rect 126 866 2156 926
rect 0 726 1048 806
rect 0 546 66 726
rect 1108 666 1174 866
rect 2216 806 2282 986
rect 3324 926 3390 1136
rect 4432 1076 4498 1262
rect 3450 986 4498 1076
rect 2342 866 4372 926
rect 1234 726 3264 806
rect 126 606 2156 666
rect 0 486 1048 546
rect 0 306 66 486
rect 1108 426 1174 606
rect 2216 546 2282 726
rect 3324 666 3390 866
rect 4432 806 4498 986
rect 3450 726 4498 806
rect 2342 606 4372 666
rect 1234 486 3264 546
rect 126 366 2156 426
rect 0 246 1048 306
rect 0 66 66 246
rect 1108 186 1174 366
rect 2216 306 2282 486
rect 3324 426 3390 606
rect 4432 546 4498 726
rect 3450 486 4498 546
rect 2342 366 4372 426
rect 1234 246 3264 306
rect 126 126 2156 186
rect 2216 66 2282 246
rect 3324 186 3390 366
rect 4432 306 4498 486
rect 3450 246 4498 306
rect 2342 126 4372 186
rect 4432 66 4498 246
rect 0 0 4498 66
<< metal5 >>
rect 0 0 4498 4610
<< labels >>
rlabel metal4 s 4432 4364 4498 4544 6 C0
port 1 nsew
rlabel metal4 s 4432 4124 4498 4304 6 C0
port 1 nsew
rlabel metal4 s 4432 3884 4498 4064 6 C0
port 1 nsew
rlabel metal4 s 4432 3624 4498 3804 6 C0
port 1 nsew
rlabel metal4 s 4432 3348 4498 3534 6 C0
port 1 nsew
rlabel metal4 s 4432 3078 4498 3258 6 C0
port 1 nsew
rlabel metal4 s 4432 2818 4498 2998 6 C0
port 1 nsew
rlabel metal4 s 4432 2578 4498 2758 6 C0
port 1 nsew
rlabel metal4 s 4432 2338 4498 2518 6 C0
port 1 nsew
rlabel metal4 s 4432 2092 4498 2272 6 C0
port 1 nsew
rlabel metal4 s 4432 1852 4498 2032 6 C0
port 1 nsew
rlabel metal4 s 4432 1612 4498 1792 6 C0
port 1 nsew
rlabel metal4 s 4432 1352 4498 1532 6 C0
port 1 nsew
rlabel metal4 s 4432 1076 4498 1262 6 C0
port 1 nsew
rlabel metal4 s 4432 806 4498 986 6 C0
port 1 nsew
rlabel metal4 s 4432 546 4498 726 6 C0
port 1 nsew
rlabel metal4 s 4432 306 4498 486 6 C0
port 1 nsew
rlabel metal4 s 4432 66 4498 246 6 C0
port 1 nsew
rlabel metal4 s 3450 4304 4498 4364 6 C0
port 1 nsew
rlabel metal4 s 3450 4064 4498 4124 6 C0
port 1 nsew
rlabel metal4 s 3450 3804 4498 3884 6 C0
port 1 nsew
rlabel metal4 s 3450 3534 4498 3624 6 C0
port 1 nsew
rlabel metal4 s 3450 3258 4498 3348 6 C0
port 1 nsew
rlabel metal4 s 3450 2998 4498 3078 6 C0
port 1 nsew
rlabel metal4 s 3450 2758 4498 2818 6 C0
port 1 nsew
rlabel metal4 s 3450 2518 4498 2578 6 C0
port 1 nsew
rlabel metal4 s 3450 2032 4498 2092 6 C0
port 1 nsew
rlabel metal4 s 3450 1792 4498 1852 6 C0
port 1 nsew
rlabel metal4 s 3450 1532 4498 1612 6 C0
port 1 nsew
rlabel metal4 s 3450 1262 4498 1352 6 C0
port 1 nsew
rlabel metal4 s 3450 986 4498 1076 6 C0
port 1 nsew
rlabel metal4 s 3450 726 4498 806 6 C0
port 1 nsew
rlabel metal4 s 3450 486 4498 546 6 C0
port 1 nsew
rlabel metal4 s 3450 246 4498 306 6 C0
port 1 nsew
rlabel metal4 s 2216 4364 2282 4544 6 C0
port 1 nsew
rlabel metal4 s 2216 4124 2282 4304 6 C0
port 1 nsew
rlabel metal4 s 2216 3884 2282 4064 6 C0
port 1 nsew
rlabel metal4 s 2216 3624 2282 3804 6 C0
port 1 nsew
rlabel metal4 s 2216 3348 2282 3534 6 C0
port 1 nsew
rlabel metal4 s 2216 3078 2282 3258 6 C0
port 1 nsew
rlabel metal4 s 2216 2818 2282 2998 6 C0
port 1 nsew
rlabel metal4 s 2216 2578 2282 2758 6 C0
port 1 nsew
rlabel metal4 s 2216 2338 2282 2518 6 C0
port 1 nsew
rlabel metal4 s 2216 2092 2282 2272 6 C0
port 1 nsew
rlabel metal4 s 2216 1852 2282 2032 6 C0
port 1 nsew
rlabel metal4 s 2216 1612 2282 1792 6 C0
port 1 nsew
rlabel metal4 s 2216 1352 2282 1532 6 C0
port 1 nsew
rlabel metal4 s 2216 1076 2282 1262 6 C0
port 1 nsew
rlabel metal4 s 2216 806 2282 986 6 C0
port 1 nsew
rlabel metal4 s 2216 546 2282 726 6 C0
port 1 nsew
rlabel metal4 s 2216 306 2282 486 6 C0
port 1 nsew
rlabel metal4 s 2216 66 2282 246 6 C0
port 1 nsew
rlabel metal4 s 1234 4304 3264 4364 6 C0
port 1 nsew
rlabel metal4 s 1234 4064 3264 4124 6 C0
port 1 nsew
rlabel metal4 s 1234 3804 3264 3884 6 C0
port 1 nsew
rlabel metal4 s 1234 3534 3264 3624 6 C0
port 1 nsew
rlabel metal4 s 1234 3258 3264 3348 6 C0
port 1 nsew
rlabel metal4 s 1234 2998 3264 3078 6 C0
port 1 nsew
rlabel metal4 s 1234 2758 3264 2818 6 C0
port 1 nsew
rlabel metal4 s 1234 2518 3264 2578 6 C0
port 1 nsew
rlabel metal4 s 1234 2032 3264 2092 6 C0
port 1 nsew
rlabel metal4 s 1234 1792 3264 1852 6 C0
port 1 nsew
rlabel metal4 s 1234 1532 3264 1612 6 C0
port 1 nsew
rlabel metal4 s 1234 1262 3264 1352 6 C0
port 1 nsew
rlabel metal4 s 1234 986 3264 1076 6 C0
port 1 nsew
rlabel metal4 s 1234 726 3264 806 6 C0
port 1 nsew
rlabel metal4 s 1234 486 3264 546 6 C0
port 1 nsew
rlabel metal4 s 1234 246 3264 306 6 C0
port 1 nsew
rlabel metal4 s 0 4544 4498 4610 6 C0
port 1 nsew
rlabel metal4 s 0 4364 66 4544 6 C0
port 1 nsew
rlabel metal4 s 0 4304 1048 4364 6 C0
port 1 nsew
rlabel metal4 s 0 4124 66 4304 6 C0
port 1 nsew
rlabel metal4 s 0 4064 1048 4124 6 C0
port 1 nsew
rlabel metal4 s 0 3884 66 4064 6 C0
port 1 nsew
rlabel metal4 s 0 3804 1048 3884 6 C0
port 1 nsew
rlabel metal4 s 0 3624 66 3804 6 C0
port 1 nsew
rlabel metal4 s 0 3534 1048 3624 6 C0
port 1 nsew
rlabel metal4 s 0 3348 66 3534 6 C0
port 1 nsew
rlabel metal4 s 0 3258 1048 3348 6 C0
port 1 nsew
rlabel metal4 s 0 3078 66 3258 6 C0
port 1 nsew
rlabel metal4 s 0 2998 1048 3078 6 C0
port 1 nsew
rlabel metal4 s 0 2818 66 2998 6 C0
port 1 nsew
rlabel metal4 s 0 2758 1048 2818 6 C0
port 1 nsew
rlabel metal4 s 0 2578 66 2758 6 C0
port 1 nsew
rlabel metal4 s 0 2518 1048 2578 6 C0
port 1 nsew
rlabel metal4 s 0 2338 66 2518 6 C0
port 1 nsew
rlabel metal4 s 0 2272 4498 2338 6 C0
port 1 nsew
rlabel metal4 s 0 2092 66 2272 6 C0
port 1 nsew
rlabel metal4 s 0 2032 1048 2092 6 C0
port 1 nsew
rlabel metal4 s 0 1852 66 2032 6 C0
port 1 nsew
rlabel metal4 s 0 1792 1048 1852 6 C0
port 1 nsew
rlabel metal4 s 0 1612 66 1792 6 C0
port 1 nsew
rlabel metal4 s 0 1532 1048 1612 6 C0
port 1 nsew
rlabel metal4 s 0 1352 66 1532 6 C0
port 1 nsew
rlabel metal4 s 0 1262 1048 1352 6 C0
port 1 nsew
rlabel metal4 s 0 1076 66 1262 6 C0
port 1 nsew
rlabel metal4 s 0 986 1048 1076 6 C0
port 1 nsew
rlabel metal4 s 0 806 66 986 6 C0
port 1 nsew
rlabel metal4 s 0 726 1048 806 6 C0
port 1 nsew
rlabel metal4 s 0 546 66 726 6 C0
port 1 nsew
rlabel metal4 s 0 486 1048 546 6 C0
port 1 nsew
rlabel metal4 s 0 306 66 486 6 C0
port 1 nsew
rlabel metal4 s 0 246 1048 306 6 C0
port 1 nsew
rlabel metal4 s 0 66 66 246 6 C0
port 1 nsew
rlabel metal4 s 0 0 4498 66 6 C0
port 1 nsew
rlabel metal4 s 3324 4244 3390 4424 6 C1
port 2 nsew
rlabel metal4 s 3324 4004 3390 4184 6 C1
port 2 nsew
rlabel metal4 s 3324 3744 3390 3944 6 C1
port 2 nsew
rlabel metal4 s 3324 3474 3390 3684 6 C1
port 2 nsew
rlabel metal4 s 3324 3198 3390 3408 6 C1
port 2 nsew
rlabel metal4 s 3324 2938 3390 3138 6 C1
port 2 nsew
rlabel metal4 s 3324 2698 3390 2878 6 C1
port 2 nsew
rlabel metal4 s 3324 2458 3390 2638 6 C1
port 2 nsew
rlabel metal4 s 3324 1972 3390 2152 6 C1
port 2 nsew
rlabel metal4 s 3324 1732 3390 1912 6 C1
port 2 nsew
rlabel metal4 s 3324 1472 3390 1672 6 C1
port 2 nsew
rlabel metal4 s 3324 1202 3390 1412 6 C1
port 2 nsew
rlabel metal4 s 3324 926 3390 1136 6 C1
port 2 nsew
rlabel metal4 s 3324 666 3390 866 6 C1
port 2 nsew
rlabel metal4 s 3324 426 3390 606 6 C1
port 2 nsew
rlabel metal4 s 3324 186 3390 366 6 C1
port 2 nsew
rlabel metal4 s 2342 4424 4372 4484 6 C1
port 2 nsew
rlabel metal4 s 2342 4184 4372 4244 6 C1
port 2 nsew
rlabel metal4 s 2342 3944 4372 4004 6 C1
port 2 nsew
rlabel metal4 s 2342 3684 4372 3744 6 C1
port 2 nsew
rlabel metal4 s 2342 3408 4372 3474 6 C1
port 2 nsew
rlabel metal4 s 2342 3138 4372 3198 6 C1
port 2 nsew
rlabel metal4 s 2342 2878 4372 2938 6 C1
port 2 nsew
rlabel metal4 s 2342 2638 4372 2698 6 C1
port 2 nsew
rlabel metal4 s 2342 2398 4372 2458 6 C1
port 2 nsew
rlabel metal4 s 2342 2152 4372 2212 6 C1
port 2 nsew
rlabel metal4 s 2342 1912 4372 1972 6 C1
port 2 nsew
rlabel metal4 s 2342 1672 4372 1732 6 C1
port 2 nsew
rlabel metal4 s 2342 1412 4372 1472 6 C1
port 2 nsew
rlabel metal4 s 2342 1136 4372 1202 6 C1
port 2 nsew
rlabel metal4 s 2342 866 4372 926 6 C1
port 2 nsew
rlabel metal4 s 2342 606 4372 666 6 C1
port 2 nsew
rlabel metal4 s 2342 366 4372 426 6 C1
port 2 nsew
rlabel metal4 s 2342 126 4372 186 6 C1
port 2 nsew
rlabel metal4 s 1108 4244 1174 4424 6 C1
port 2 nsew
rlabel metal4 s 1108 4004 1174 4184 6 C1
port 2 nsew
rlabel metal4 s 1108 3744 1174 3944 6 C1
port 2 nsew
rlabel metal4 s 1108 3474 1174 3684 6 C1
port 2 nsew
rlabel metal4 s 1108 3198 1174 3408 6 C1
port 2 nsew
rlabel metal4 s 1108 2938 1174 3138 6 C1
port 2 nsew
rlabel metal4 s 1108 2698 1174 2878 6 C1
port 2 nsew
rlabel metal4 s 1108 2458 1174 2638 6 C1
port 2 nsew
rlabel metal4 s 1108 1972 1174 2152 6 C1
port 2 nsew
rlabel metal4 s 1108 1732 1174 1912 6 C1
port 2 nsew
rlabel metal4 s 1108 1472 1174 1672 6 C1
port 2 nsew
rlabel metal4 s 1108 1202 1174 1412 6 C1
port 2 nsew
rlabel metal4 s 1108 926 1174 1136 6 C1
port 2 nsew
rlabel metal4 s 1108 666 1174 866 6 C1
port 2 nsew
rlabel metal4 s 1108 426 1174 606 6 C1
port 2 nsew
rlabel metal4 s 1108 186 1174 366 6 C1
port 2 nsew
rlabel metal4 s 126 4424 2156 4484 6 C1
port 2 nsew
rlabel metal4 s 126 4184 2156 4244 6 C1
port 2 nsew
rlabel metal4 s 126 3944 2156 4004 6 C1
port 2 nsew
rlabel metal4 s 126 3684 2156 3744 6 C1
port 2 nsew
rlabel metal4 s 126 3408 2156 3474 6 C1
port 2 nsew
rlabel metal4 s 126 3138 2156 3198 6 C1
port 2 nsew
rlabel metal4 s 126 2878 2156 2938 6 C1
port 2 nsew
rlabel metal4 s 126 2638 2156 2698 6 C1
port 2 nsew
rlabel metal4 s 126 2398 2156 2458 6 C1
port 2 nsew
rlabel metal4 s 126 2152 2156 2212 6 C1
port 2 nsew
rlabel metal4 s 126 1912 2156 1972 6 C1
port 2 nsew
rlabel metal4 s 126 1672 2156 1732 6 C1
port 2 nsew
rlabel metal4 s 126 1412 2156 1472 6 C1
port 2 nsew
rlabel metal4 s 126 1136 2156 1202 6 C1
port 2 nsew
rlabel metal4 s 126 866 2156 926 6 C1
port 2 nsew
rlabel metal4 s 126 606 2156 666 6 C1
port 2 nsew
rlabel metal4 s 126 366 2156 426 6 C1
port 2 nsew
rlabel metal4 s 126 126 2156 186 6 C1
port 2 nsew
rlabel metal5 s 0 0 4498 4610 6 M5
port 3 nsew
rlabel pwell s 1179 1269 1189 1279 6 SUB
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 4498 4610
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1551524
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 1550950
<< end >>
