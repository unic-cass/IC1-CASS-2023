* NGSPICE file created from sky130_ef_sc_hd__fakediode_2.ext - technology: sky130A

.subckt sky130_ef_sc_hd__fakediode_2 DIODE VGND VPWR VPB VNB
D0 VNB a_31_39# sky130_fd_pr__diode_pw2nd_05v5 pj=2.64e+06 area=4.347e+11
.ends

