magic
tech sky130A
magscale 1 2
timestamp 1676037725
use sky130_fd_io__gnd2gnd_diff  sky130_fd_io__gnd2gnd_diff_0
array 0 3 824 0 0 3052
timestamp 1676037725
transform 1 0 632 0 1 220
box 0 0 300 3000
use sky130_fd_io__gnd2gnd_tap  sky130_fd_io__gnd2gnd_tap_0
array 0 4 824 0 0 3052
timestamp 1676037725
transform 1 0 220 0 1 220
box 0 0 300 3000
use sky130_fd_pr__tpl1__example_55959141808685  sky130_fd_pr__tpl1__example_55959141808685_0
timestamp 1676037725
transform 1 0 26 0 1 115
box 0 0 1 1
use sky130_fd_pr__tpl1__example_55959141808685  sky130_fd_pr__tpl1__example_55959141808685_1
timestamp 1676037725
transform 1 0 3928 0 1 115
box 0 0 1 1
use sky130_fd_pr__tpl1__example_55959141808686  sky130_fd_pr__tpl1__example_55959141808686_0
timestamp 1676037725
transform -1 0 3942 0 1 26
box 0 0 1 1
use sky130_fd_pr__tpl1__example_55959141808686  sky130_fd_pr__tpl1__example_55959141808686_1
timestamp 1676037725
transform -1 0 3952 0 1 3332
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808684  sky130_fd_pr__via_l1m1__example_55959141808684_0
timestamp 1676037725
transform 1 0 3955 0 1 160
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808684  sky130_fd_pr__via_l1m1__example_55959141808684_1
timestamp 1676037725
transform 1 0 53 0 1 160
box 0 0 1 1
<< properties >>
string GDS_END 8053710
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 8052078
<< end >>
