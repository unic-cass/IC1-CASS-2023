magic
tech sky130A
magscale 1 2
timestamp 1676037725
<< nwell >>
rect 2129 954 3345 1655
rect 5141 404 6151 1104
<< pwell >>
rect 2169 1974 5668 2060
rect 2169 1952 3264 1974
rect 2166 1760 3264 1952
rect 2169 -3 5107 83
<< mvnmos >>
rect 2248 1786 2368 1926
rect 2424 1786 2544 1926
rect 2713 1786 2833 1926
rect 2889 1786 3009 1926
rect 3065 1786 3185 1926
<< mvpmos >>
rect 2248 1388 2368 1588
rect 2424 1388 2544 1588
rect 2713 1388 2833 1588
rect 2889 1388 3009 1588
rect 3065 1388 3185 1588
rect 2248 1120 2368 1320
rect 2424 1120 2544 1320
rect 2713 1120 2833 1320
rect 2889 1120 3009 1320
rect 3065 1120 3185 1320
<< mvndiff >>
rect 2192 1900 2248 1926
rect 2192 1866 2203 1900
rect 2237 1866 2248 1900
rect 2192 1832 2248 1866
rect 2192 1798 2203 1832
rect 2237 1798 2248 1832
rect 2192 1786 2248 1798
rect 2368 1900 2424 1926
rect 2368 1866 2379 1900
rect 2413 1866 2424 1900
rect 2368 1832 2424 1866
rect 2368 1798 2379 1832
rect 2413 1798 2424 1832
rect 2368 1786 2424 1798
rect 2544 1900 2597 1926
rect 2544 1866 2555 1900
rect 2589 1866 2597 1900
rect 2544 1832 2597 1866
rect 2544 1798 2555 1832
rect 2589 1798 2597 1832
rect 2544 1786 2597 1798
rect 2657 1900 2713 1926
rect 2657 1866 2668 1900
rect 2702 1866 2713 1900
rect 2657 1832 2713 1866
rect 2657 1798 2668 1832
rect 2702 1798 2713 1832
rect 2657 1786 2713 1798
rect 2833 1900 2889 1926
rect 2833 1866 2844 1900
rect 2878 1866 2889 1900
rect 2833 1832 2889 1866
rect 2833 1798 2844 1832
rect 2878 1798 2889 1832
rect 2833 1786 2889 1798
rect 3009 1900 3065 1926
rect 3009 1866 3020 1900
rect 3054 1866 3065 1900
rect 3009 1832 3065 1866
rect 3009 1798 3020 1832
rect 3054 1798 3065 1832
rect 3009 1786 3065 1798
rect 3185 1900 3238 1926
rect 3185 1866 3196 1900
rect 3230 1866 3238 1900
rect 3185 1832 3238 1866
rect 3185 1798 3196 1832
rect 3230 1798 3238 1832
rect 3185 1786 3238 1798
<< mvpdiff >>
rect 2195 1570 2248 1588
rect 2195 1536 2203 1570
rect 2237 1536 2248 1570
rect 2195 1502 2248 1536
rect 2195 1468 2203 1502
rect 2237 1468 2248 1502
rect 2195 1434 2248 1468
rect 2195 1400 2203 1434
rect 2237 1400 2248 1434
rect 2195 1388 2248 1400
rect 2368 1502 2424 1588
rect 2368 1468 2379 1502
rect 2413 1468 2424 1502
rect 2368 1434 2424 1468
rect 2368 1400 2379 1434
rect 2413 1400 2424 1434
rect 2368 1388 2424 1400
rect 2544 1570 2597 1588
rect 2544 1536 2555 1570
rect 2589 1536 2597 1570
rect 2544 1502 2597 1536
rect 2544 1468 2555 1502
rect 2589 1468 2597 1502
rect 2544 1434 2597 1468
rect 2544 1400 2555 1434
rect 2589 1400 2597 1434
rect 2544 1388 2597 1400
rect 2660 1570 2713 1588
rect 2660 1536 2668 1570
rect 2702 1536 2713 1570
rect 2660 1502 2713 1536
rect 2660 1468 2668 1502
rect 2702 1468 2713 1502
rect 2660 1434 2713 1468
rect 2660 1400 2668 1434
rect 2702 1400 2713 1434
rect 2660 1388 2713 1400
rect 2833 1502 2889 1588
rect 2833 1468 2844 1502
rect 2878 1468 2889 1502
rect 2833 1434 2889 1468
rect 2833 1400 2844 1434
rect 2878 1400 2889 1434
rect 2833 1388 2889 1400
rect 3009 1570 3065 1588
rect 3009 1536 3020 1570
rect 3054 1536 3065 1570
rect 3009 1502 3065 1536
rect 3009 1468 3020 1502
rect 3054 1468 3065 1502
rect 3009 1434 3065 1468
rect 3009 1400 3020 1434
rect 3054 1400 3065 1434
rect 3009 1388 3065 1400
rect 3185 1570 3238 1588
rect 3185 1536 3196 1570
rect 3230 1536 3238 1570
rect 3185 1502 3238 1536
rect 3185 1468 3196 1502
rect 3230 1468 3238 1502
rect 3185 1434 3238 1468
rect 3185 1400 3196 1434
rect 3230 1400 3238 1434
rect 3185 1388 3238 1400
rect 2195 1308 2248 1320
rect 2195 1274 2203 1308
rect 2237 1274 2248 1308
rect 2195 1240 2248 1274
rect 2195 1206 2203 1240
rect 2237 1206 2248 1240
rect 2195 1172 2248 1206
rect 2195 1138 2203 1172
rect 2237 1138 2248 1172
rect 2195 1120 2248 1138
rect 2368 1308 2424 1320
rect 2368 1274 2379 1308
rect 2413 1274 2424 1308
rect 2368 1240 2424 1274
rect 2368 1206 2379 1240
rect 2413 1206 2424 1240
rect 2368 1172 2424 1206
rect 2368 1138 2379 1172
rect 2413 1138 2424 1172
rect 2368 1120 2424 1138
rect 2544 1308 2597 1320
rect 2544 1274 2555 1308
rect 2589 1274 2597 1308
rect 2544 1240 2597 1274
rect 2544 1206 2555 1240
rect 2589 1206 2597 1240
rect 2544 1172 2597 1206
rect 2544 1138 2555 1172
rect 2589 1138 2597 1172
rect 2544 1120 2597 1138
rect 2660 1308 2713 1320
rect 2660 1274 2668 1308
rect 2702 1274 2713 1308
rect 2660 1240 2713 1274
rect 2660 1206 2668 1240
rect 2702 1206 2713 1240
rect 2660 1172 2713 1206
rect 2660 1138 2668 1172
rect 2702 1138 2713 1172
rect 2660 1120 2713 1138
rect 2833 1308 2889 1320
rect 2833 1274 2844 1308
rect 2878 1274 2889 1308
rect 2833 1240 2889 1274
rect 2833 1206 2844 1240
rect 2878 1206 2889 1240
rect 2833 1172 2889 1206
rect 2833 1138 2844 1172
rect 2878 1138 2889 1172
rect 2833 1120 2889 1138
rect 3009 1308 3065 1320
rect 3009 1274 3020 1308
rect 3054 1274 3065 1308
rect 3009 1240 3065 1274
rect 3009 1206 3020 1240
rect 3054 1206 3065 1240
rect 3009 1172 3065 1206
rect 3009 1138 3020 1172
rect 3054 1138 3065 1172
rect 3009 1120 3065 1138
rect 3185 1308 3238 1320
rect 3185 1274 3196 1308
rect 3230 1274 3238 1308
rect 3185 1240 3238 1274
rect 3185 1206 3196 1240
rect 3230 1206 3238 1240
rect 3185 1172 3238 1206
rect 3185 1138 3196 1172
rect 3230 1138 3238 1172
rect 3185 1120 3238 1138
<< mvndiffc >>
rect 2203 1866 2237 1900
rect 2203 1798 2237 1832
rect 2379 1866 2413 1900
rect 2379 1798 2413 1832
rect 2555 1866 2589 1900
rect 2555 1798 2589 1832
rect 2668 1866 2702 1900
rect 2668 1798 2702 1832
rect 2844 1866 2878 1900
rect 2844 1798 2878 1832
rect 3020 1866 3054 1900
rect 3020 1798 3054 1832
rect 3196 1866 3230 1900
rect 3196 1798 3230 1832
<< mvpdiffc >>
rect 2203 1536 2237 1570
rect 2203 1468 2237 1502
rect 2203 1400 2237 1434
rect 2379 1468 2413 1502
rect 2379 1400 2413 1434
rect 2555 1536 2589 1570
rect 2555 1468 2589 1502
rect 2555 1400 2589 1434
rect 2668 1536 2702 1570
rect 2668 1468 2702 1502
rect 2668 1400 2702 1434
rect 2844 1468 2878 1502
rect 2844 1400 2878 1434
rect 3020 1536 3054 1570
rect 3020 1468 3054 1502
rect 3020 1400 3054 1434
rect 3196 1536 3230 1570
rect 3196 1468 3230 1502
rect 3196 1400 3230 1434
rect 2203 1274 2237 1308
rect 2203 1206 2237 1240
rect 2203 1138 2237 1172
rect 2379 1274 2413 1308
rect 2379 1206 2413 1240
rect 2379 1138 2413 1172
rect 2555 1274 2589 1308
rect 2555 1206 2589 1240
rect 2555 1138 2589 1172
rect 2668 1274 2702 1308
rect 2668 1206 2702 1240
rect 2668 1138 2702 1172
rect 2844 1274 2878 1308
rect 2844 1206 2878 1240
rect 2844 1138 2878 1172
rect 3020 1274 3054 1308
rect 3020 1206 3054 1240
rect 3020 1138 3054 1172
rect 3196 1274 3230 1308
rect 3196 1206 3230 1240
rect 3196 1138 3230 1172
<< mvpsubdiff >>
rect 2195 2000 2219 2034
rect 2253 2000 2288 2034
rect 2322 2000 2357 2034
rect 2391 2000 2426 2034
rect 2460 2000 2495 2034
rect 2529 2000 2564 2034
rect 2598 2000 2633 2034
rect 2667 2000 2702 2034
rect 2736 2000 2771 2034
rect 2805 2000 2840 2034
rect 2874 2000 2909 2034
rect 2943 2000 2978 2034
rect 3012 2000 3047 2034
rect 3081 2000 3116 2034
rect 3150 2000 3185 2034
rect 3219 2000 3254 2034
rect 3288 2000 3323 2034
rect 3357 2000 3392 2034
rect 3426 2000 3461 2034
rect 3495 2000 3530 2034
rect 3564 2000 3599 2034
rect 3633 2000 3668 2034
rect 3702 2000 3737 2034
rect 3771 2000 3806 2034
rect 3840 2000 3875 2034
rect 3909 2000 3944 2034
rect 3978 2000 4013 2034
rect 4047 2000 4082 2034
rect 4116 2000 4151 2034
rect 4185 2000 4220 2034
rect 4254 2000 4289 2034
rect 4323 2000 4358 2034
rect 4392 2000 4427 2034
rect 4461 2000 4496 2034
rect 4530 2000 4564 2034
rect 4598 2000 4632 2034
rect 4666 2000 4700 2034
rect 4734 2000 4768 2034
rect 4802 2000 4836 2034
rect 4870 2000 4904 2034
rect 4938 2000 4972 2034
rect 5006 2000 5040 2034
rect 5074 2000 5108 2034
rect 5142 2000 5176 2034
rect 5210 2000 5244 2034
rect 5278 2000 5312 2034
rect 5346 2000 5380 2034
rect 5414 2000 5448 2034
rect 5482 2000 5516 2034
rect 5550 2000 5584 2034
rect 5618 2000 5642 2034
rect 2195 23 2219 57
rect 2253 23 2288 57
rect 2322 23 2357 57
rect 2391 23 2426 57
rect 2460 23 2495 57
rect 2529 23 2564 57
rect 2598 23 2633 57
rect 2667 23 2702 57
rect 2736 23 2771 57
rect 2805 23 2840 57
rect 2874 23 2909 57
rect 2943 23 2978 57
rect 3012 23 3047 57
rect 3081 23 3116 57
rect 3150 23 3185 57
rect 3219 23 3254 57
rect 3288 23 3323 57
rect 3357 23 3391 57
rect 3425 23 3459 57
rect 3493 23 3527 57
rect 3561 23 3595 57
rect 3629 23 3663 57
rect 3697 23 3731 57
rect 3765 23 3799 57
rect 3833 23 3867 57
rect 3901 23 3935 57
rect 3969 23 4003 57
rect 4037 23 4071 57
rect 4105 23 4139 57
rect 4173 23 4207 57
rect 4241 23 4275 57
rect 4309 23 4343 57
rect 4377 23 4411 57
rect 4445 23 4479 57
rect 4513 23 4547 57
rect 4581 23 4615 57
rect 4649 23 4683 57
rect 4717 23 4751 57
rect 4785 23 4819 57
rect 4853 23 4887 57
rect 4921 23 4955 57
rect 4989 23 5023 57
rect 5057 23 5081 57
<< mvpsubdiffcont >>
rect 2219 2000 2253 2034
rect 2288 2000 2322 2034
rect 2357 2000 2391 2034
rect 2426 2000 2460 2034
rect 2495 2000 2529 2034
rect 2564 2000 2598 2034
rect 2633 2000 2667 2034
rect 2702 2000 2736 2034
rect 2771 2000 2805 2034
rect 2840 2000 2874 2034
rect 2909 2000 2943 2034
rect 2978 2000 3012 2034
rect 3047 2000 3081 2034
rect 3116 2000 3150 2034
rect 3185 2000 3219 2034
rect 3254 2000 3288 2034
rect 3323 2000 3357 2034
rect 3392 2000 3426 2034
rect 3461 2000 3495 2034
rect 3530 2000 3564 2034
rect 3599 2000 3633 2034
rect 3668 2000 3702 2034
rect 3737 2000 3771 2034
rect 3806 2000 3840 2034
rect 3875 2000 3909 2034
rect 3944 2000 3978 2034
rect 4013 2000 4047 2034
rect 4082 2000 4116 2034
rect 4151 2000 4185 2034
rect 4220 2000 4254 2034
rect 4289 2000 4323 2034
rect 4358 2000 4392 2034
rect 4427 2000 4461 2034
rect 4496 2000 4530 2034
rect 4564 2000 4598 2034
rect 4632 2000 4666 2034
rect 4700 2000 4734 2034
rect 4768 2000 4802 2034
rect 4836 2000 4870 2034
rect 4904 2000 4938 2034
rect 4972 2000 5006 2034
rect 5040 2000 5074 2034
rect 5108 2000 5142 2034
rect 5176 2000 5210 2034
rect 5244 2000 5278 2034
rect 5312 2000 5346 2034
rect 5380 2000 5414 2034
rect 5448 2000 5482 2034
rect 5516 2000 5550 2034
rect 5584 2000 5618 2034
rect 2219 23 2253 57
rect 2288 23 2322 57
rect 2357 23 2391 57
rect 2426 23 2460 57
rect 2495 23 2529 57
rect 2564 23 2598 57
rect 2633 23 2667 57
rect 2702 23 2736 57
rect 2771 23 2805 57
rect 2840 23 2874 57
rect 2909 23 2943 57
rect 2978 23 3012 57
rect 3047 23 3081 57
rect 3116 23 3150 57
rect 3185 23 3219 57
rect 3254 23 3288 57
rect 3323 23 3357 57
rect 3391 23 3425 57
rect 3459 23 3493 57
rect 3527 23 3561 57
rect 3595 23 3629 57
rect 3663 23 3697 57
rect 3731 23 3765 57
rect 3799 23 3833 57
rect 3867 23 3901 57
rect 3935 23 3969 57
rect 4003 23 4037 57
rect 4071 23 4105 57
rect 4139 23 4173 57
rect 4207 23 4241 57
rect 4275 23 4309 57
rect 4343 23 4377 57
rect 4411 23 4445 57
rect 4479 23 4513 57
rect 4547 23 4581 57
rect 4615 23 4649 57
rect 4683 23 4717 57
rect 4751 23 4785 57
rect 4819 23 4853 57
rect 4887 23 4921 57
rect 4955 23 4989 57
rect 5023 23 5057 57
<< poly >>
rect 2248 1926 2368 1952
rect 2424 1926 2544 1952
rect 2713 1926 2833 1952
rect 2889 1926 3009 1952
rect 3065 1926 3185 1952
rect 2248 1738 2368 1786
rect 2248 1704 2289 1738
rect 2323 1704 2368 1738
rect 2248 1670 2368 1704
rect 2248 1636 2289 1670
rect 2323 1636 2368 1670
rect 2248 1588 2368 1636
rect 2424 1738 2544 1786
rect 2424 1704 2467 1738
rect 2501 1704 2544 1738
rect 2424 1670 2544 1704
rect 2424 1636 2467 1670
rect 2501 1636 2544 1670
rect 2424 1588 2544 1636
rect 2713 1738 2833 1786
rect 2713 1704 2754 1738
rect 2788 1704 2833 1738
rect 2713 1670 2833 1704
rect 2713 1636 2754 1670
rect 2788 1636 2833 1670
rect 2713 1588 2833 1636
rect 2889 1738 3009 1786
rect 2889 1704 2932 1738
rect 2966 1704 3009 1738
rect 2889 1670 3009 1704
rect 2889 1636 2932 1670
rect 2966 1636 3009 1670
rect 2889 1588 3009 1636
rect 3065 1738 3185 1786
rect 3065 1704 3109 1738
rect 3143 1704 3185 1738
rect 3065 1670 3185 1704
rect 3065 1636 3109 1670
rect 3143 1636 3185 1670
rect 3065 1588 3185 1636
rect 2248 1320 2368 1388
rect 2424 1320 2544 1388
rect 2713 1320 2833 1388
rect 2889 1320 3009 1388
rect 3065 1320 3185 1388
rect 3351 1346 3471 1362
rect 3527 1346 3647 1362
rect 3703 1346 3823 1362
rect 2248 1094 2368 1120
rect 2424 1094 2544 1120
rect 2713 1094 2833 1120
rect 2889 1094 3009 1120
rect 3065 1094 3185 1120
<< polycont >>
rect 2289 1704 2323 1738
rect 2289 1636 2323 1670
rect 2467 1704 2501 1738
rect 2467 1636 2501 1670
rect 2754 1704 2788 1738
rect 2754 1636 2788 1670
rect 2932 1704 2966 1738
rect 2932 1636 2966 1670
rect 3109 1704 3143 1738
rect 3109 1636 3143 1670
<< locali >>
rect 2195 2000 2211 2034
rect 2253 2000 2284 2034
rect 2322 2000 2357 2034
rect 2391 2000 2426 2034
rect 2464 2000 2495 2034
rect 2537 2000 2564 2034
rect 2610 2000 2633 2034
rect 2683 2000 2702 2034
rect 2756 2000 2771 2034
rect 2829 2000 2840 2034
rect 2902 2000 2909 2034
rect 2975 2000 2978 2034
rect 3012 2000 3014 2034
rect 3081 2000 3087 2034
rect 3150 2000 3160 2034
rect 3219 2000 3233 2034
rect 3288 2000 3306 2034
rect 3357 2000 3378 2034
rect 3426 2000 3450 2034
rect 3495 2000 3522 2034
rect 3564 2000 3594 2034
rect 3633 2000 3666 2034
rect 3702 2000 3737 2034
rect 3772 2000 3806 2034
rect 3844 2000 3875 2034
rect 3916 2000 3944 2034
rect 3988 2000 4013 2034
rect 4060 2000 4082 2034
rect 4132 2000 4151 2034
rect 4204 2000 4220 2034
rect 4276 2000 4289 2034
rect 4348 2000 4358 2034
rect 4420 2000 4427 2034
rect 4492 2000 4496 2034
rect 4598 2000 4602 2034
rect 4666 2000 4674 2034
rect 4734 2000 4746 2034
rect 4802 2000 4818 2034
rect 4870 2000 4890 2034
rect 4938 2000 4962 2034
rect 5006 2000 5034 2034
rect 5074 2000 5106 2034
rect 5142 2000 5176 2034
rect 5212 2000 5244 2034
rect 5284 2000 5312 2034
rect 5356 2000 5380 2034
rect 5428 2000 5448 2034
rect 5500 2000 5516 2034
rect 5572 2000 5584 2034
rect 2203 1900 2237 1915
rect 2203 1832 2237 1843
rect 2203 1782 2237 1798
rect 2379 1900 2413 1916
rect 2379 1832 2413 1866
rect 2273 1704 2289 1738
rect 2323 1704 2339 1738
rect 2273 1670 2339 1704
rect 2273 1655 2289 1670
rect 2323 1655 2339 1670
rect 1460 1586 1494 1624
rect 2270 1636 2289 1655
rect 2270 1621 2308 1636
rect 2379 1586 2413 1798
rect 2555 1900 2589 1915
rect 2555 1832 2589 1843
rect 2555 1782 2589 1798
rect 2668 1900 2702 1915
rect 2668 1832 2702 1843
rect 2668 1782 2702 1798
rect 2844 1900 2878 1916
rect 2844 1832 2878 1866
rect 2451 1704 2467 1738
rect 2501 1729 2517 1738
rect 2451 1695 2472 1704
rect 2506 1695 2517 1729
rect 2738 1704 2754 1738
rect 2788 1704 2804 1738
rect 2738 1699 2804 1704
rect 2451 1670 2517 1695
rect 2451 1636 2467 1670
rect 2501 1657 2517 1670
rect 2733 1670 2771 1699
rect 2733 1665 2754 1670
rect 2506 1636 2517 1657
rect 2738 1636 2754 1665
rect 2788 1636 2804 1665
rect 2844 1586 2878 1798
rect 3020 1900 3054 1915
rect 3020 1832 3054 1843
rect 3020 1782 3054 1798
rect 3196 1900 3230 1916
rect 3196 1832 3230 1866
rect 2916 1704 2932 1738
rect 2966 1731 2982 1738
rect 2916 1697 2934 1704
rect 2968 1697 2982 1731
rect 2916 1670 2982 1697
rect 2916 1636 2932 1670
rect 2966 1659 2982 1670
rect 2968 1636 2982 1659
rect 3093 1704 3109 1738
rect 3143 1704 3159 1738
rect 3093 1670 3159 1704
rect 3093 1636 3109 1670
rect 3143 1636 3159 1670
rect 2203 1570 2413 1586
rect 2237 1552 2413 1570
rect 2555 1570 2589 1586
rect 2203 1502 2237 1536
rect 2203 1434 2237 1468
rect 2379 1502 2413 1518
rect 2379 1434 2413 1468
rect 2203 1376 2206 1400
rect 2203 1338 2240 1376
rect 2203 1308 2206 1338
rect 2379 1308 2413 1400
rect 2203 1240 2237 1274
rect 2203 1172 2237 1206
rect 2203 1092 2237 1138
rect 2379 1240 2413 1274
rect 2379 1172 2413 1206
rect 2379 1122 2413 1138
rect 2555 1502 2589 1536
rect 2555 1434 2589 1468
rect 2555 1308 2589 1400
rect 2555 1240 2589 1274
rect 2555 1198 2589 1206
rect 2555 1126 2589 1138
rect 2668 1570 2878 1586
rect 2702 1552 2878 1570
rect 3020 1570 3054 1586
rect 2668 1527 2702 1536
rect 2668 1455 2702 1468
rect 2668 1308 2702 1400
rect 2668 1240 2702 1274
rect 2668 1172 2702 1206
rect 2668 1092 2702 1138
rect 2844 1502 2878 1518
rect 2844 1434 2878 1468
rect 2844 1308 2878 1400
rect 2844 1240 2878 1274
rect 2844 1172 2878 1206
rect 2844 1122 2878 1138
rect 3020 1502 3054 1536
rect 3020 1434 3054 1468
rect 3093 1543 3159 1636
rect 3093 1509 3108 1543
rect 3142 1509 3159 1543
rect 3093 1471 3159 1509
rect 3093 1437 3108 1471
rect 3142 1437 3159 1471
rect 3093 1420 3159 1437
rect 3196 1731 3230 1798
rect 3196 1659 3230 1697
rect 3482 1659 3516 1697
rect 3196 1570 3230 1625
rect 3196 1502 3230 1536
rect 3196 1434 3230 1468
rect 3381 1562 3447 1639
rect 3381 1528 3397 1562
rect 3431 1528 3447 1562
rect 3381 1490 3447 1528
rect 3381 1456 3397 1490
rect 3431 1456 3447 1490
rect 3552 1562 3618 1674
rect 4216 1666 4250 1704
rect 3552 1528 3573 1562
rect 3607 1528 3618 1562
rect 3552 1490 3618 1528
rect 3552 1456 3573 1490
rect 3607 1456 3618 1490
rect 4016 1562 4082 1636
rect 4299 1666 4333 1704
rect 4565 1666 4599 1704
rect 4016 1528 4032 1562
rect 4066 1528 4082 1562
rect 4016 1490 4082 1528
rect 4016 1456 4032 1490
rect 4066 1456 4082 1490
rect 3381 1438 3447 1456
rect 4016 1434 4082 1456
rect 4368 1562 4434 1636
rect 5039 1706 5081 1740
rect 5115 1706 5157 1740
rect 5427 1706 5468 1740
rect 5502 1706 5542 1740
rect 4738 1666 4772 1704
rect 5161 1629 5212 1663
rect 5246 1629 5297 1663
rect 5331 1629 5381 1663
rect 5415 1629 5465 1663
rect 4368 1528 4384 1562
rect 4418 1528 4434 1562
rect 4368 1490 4434 1528
rect 4368 1456 4384 1490
rect 4418 1456 4434 1490
rect 4368 1434 4434 1456
rect 4827 1464 4861 1502
rect 3020 1308 3054 1400
rect 3020 1240 3054 1274
rect 3020 1198 3054 1206
rect 3020 1126 3054 1138
rect 3196 1308 3230 1400
rect 3196 1240 3230 1274
rect 3196 1172 3230 1206
rect 3196 1120 3230 1138
rect 5760 555 5779 589
rect 5813 555 5826 589
rect 5760 517 5826 555
rect 5760 483 5779 517
rect 5813 483 5826 517
rect 5760 422 5826 483
rect 5867 353 5901 391
rect 5960 350 5994 388
rect 2195 23 2219 57
rect 2253 23 2272 57
rect 2322 23 2345 57
rect 2391 23 2418 57
rect 2460 23 2491 57
rect 2529 23 2564 57
rect 2598 23 2633 57
rect 2671 23 2702 57
rect 2744 23 2771 57
rect 2817 23 2840 57
rect 2890 23 2909 57
rect 2962 23 2978 57
rect 3034 23 3047 57
rect 3106 23 3116 57
rect 3178 23 3185 57
rect 3250 23 3254 57
rect 3322 23 3323 57
rect 3357 23 3360 57
rect 3425 23 3432 57
rect 3493 23 3504 57
rect 3561 23 3576 57
rect 3629 23 3648 57
rect 3697 23 3720 57
rect 3765 23 3792 57
rect 3833 23 3864 57
rect 3901 23 3935 57
rect 3970 23 4003 57
rect 4042 23 4071 57
rect 4114 23 4139 57
rect 4186 23 4207 57
rect 4258 23 4275 57
rect 4330 23 4343 57
rect 4402 23 4411 57
rect 4474 23 4479 57
rect 4546 23 4547 57
rect 4581 23 4584 57
rect 4649 23 4656 57
rect 4717 23 4728 57
rect 4785 23 4800 57
rect 4853 23 4872 57
rect 4921 23 4944 57
rect 4989 23 5016 57
rect 5057 23 5081 57
<< viali >>
rect 2211 2000 2219 2034
rect 2219 2000 2245 2034
rect 2284 2000 2288 2034
rect 2288 2000 2318 2034
rect 2357 2000 2391 2034
rect 2430 2000 2460 2034
rect 2460 2000 2464 2034
rect 2503 2000 2529 2034
rect 2529 2000 2537 2034
rect 2576 2000 2598 2034
rect 2598 2000 2610 2034
rect 2649 2000 2667 2034
rect 2667 2000 2683 2034
rect 2722 2000 2736 2034
rect 2736 2000 2756 2034
rect 2795 2000 2805 2034
rect 2805 2000 2829 2034
rect 2868 2000 2874 2034
rect 2874 2000 2902 2034
rect 2941 2000 2943 2034
rect 2943 2000 2975 2034
rect 3014 2000 3047 2034
rect 3047 2000 3048 2034
rect 3087 2000 3116 2034
rect 3116 2000 3121 2034
rect 3160 2000 3185 2034
rect 3185 2000 3194 2034
rect 3233 2000 3254 2034
rect 3254 2000 3267 2034
rect 3306 2000 3323 2034
rect 3323 2000 3340 2034
rect 3378 2000 3392 2034
rect 3392 2000 3412 2034
rect 3450 2000 3461 2034
rect 3461 2000 3484 2034
rect 3522 2000 3530 2034
rect 3530 2000 3556 2034
rect 3594 2000 3599 2034
rect 3599 2000 3628 2034
rect 3666 2000 3668 2034
rect 3668 2000 3700 2034
rect 3738 2000 3771 2034
rect 3771 2000 3772 2034
rect 3810 2000 3840 2034
rect 3840 2000 3844 2034
rect 3882 2000 3909 2034
rect 3909 2000 3916 2034
rect 3954 2000 3978 2034
rect 3978 2000 3988 2034
rect 4026 2000 4047 2034
rect 4047 2000 4060 2034
rect 4098 2000 4116 2034
rect 4116 2000 4132 2034
rect 4170 2000 4185 2034
rect 4185 2000 4204 2034
rect 4242 2000 4254 2034
rect 4254 2000 4276 2034
rect 4314 2000 4323 2034
rect 4323 2000 4348 2034
rect 4386 2000 4392 2034
rect 4392 2000 4420 2034
rect 4458 2000 4461 2034
rect 4461 2000 4492 2034
rect 4530 2000 4564 2034
rect 4602 2000 4632 2034
rect 4632 2000 4636 2034
rect 4674 2000 4700 2034
rect 4700 2000 4708 2034
rect 4746 2000 4768 2034
rect 4768 2000 4780 2034
rect 4818 2000 4836 2034
rect 4836 2000 4852 2034
rect 4890 2000 4904 2034
rect 4904 2000 4924 2034
rect 4962 2000 4972 2034
rect 4972 2000 4996 2034
rect 5034 2000 5040 2034
rect 5040 2000 5068 2034
rect 5106 2000 5108 2034
rect 5108 2000 5140 2034
rect 5178 2000 5210 2034
rect 5210 2000 5212 2034
rect 5250 2000 5278 2034
rect 5278 2000 5284 2034
rect 5322 2000 5346 2034
rect 5346 2000 5356 2034
rect 5394 2000 5414 2034
rect 5414 2000 5428 2034
rect 5466 2000 5482 2034
rect 5482 2000 5500 2034
rect 5538 2000 5550 2034
rect 5550 2000 5572 2034
rect 5610 2000 5618 2034
rect 5618 2000 5644 2034
rect 2203 1915 2237 1949
rect 2203 1866 2237 1877
rect 2203 1843 2237 1866
rect 1460 1624 1494 1658
rect 2236 1621 2270 1655
rect 2308 1636 2323 1655
rect 2323 1636 2342 1655
rect 2308 1621 2342 1636
rect 2555 1915 2589 1949
rect 2555 1866 2589 1877
rect 2555 1843 2589 1866
rect 2668 1915 2702 1949
rect 2668 1866 2702 1877
rect 2668 1843 2702 1866
rect 2472 1704 2501 1729
rect 2501 1704 2506 1729
rect 2472 1695 2506 1704
rect 2699 1665 2733 1699
rect 2771 1670 2805 1699
rect 2771 1665 2788 1670
rect 2788 1665 2805 1670
rect 2472 1636 2501 1657
rect 2501 1636 2506 1657
rect 2472 1623 2506 1636
rect 3020 1915 3054 1949
rect 3020 1866 3054 1877
rect 3020 1843 3054 1866
rect 2934 1704 2966 1731
rect 2966 1704 2968 1731
rect 2934 1697 2968 1704
rect 2934 1636 2966 1659
rect 2966 1636 2968 1659
rect 2934 1625 2968 1636
rect 1460 1552 1494 1586
rect 2206 1400 2237 1410
rect 2237 1400 2240 1410
rect 2206 1376 2240 1400
rect 2206 1308 2240 1338
rect 2206 1304 2237 1308
rect 2237 1304 2240 1308
rect 2555 1172 2589 1198
rect 2555 1164 2589 1172
rect 2555 1092 2589 1126
rect 2668 1502 2702 1527
rect 2668 1493 2702 1502
rect 2668 1434 2702 1455
rect 2668 1421 2702 1434
rect 3108 1509 3142 1543
rect 3108 1437 3142 1471
rect 3196 1697 3230 1731
rect 3196 1625 3230 1659
rect 3482 1697 3516 1731
rect 4216 1704 4250 1738
rect 3482 1625 3516 1659
rect 3397 1528 3431 1562
rect 3397 1456 3431 1490
rect 3573 1528 3607 1562
rect 3573 1456 3607 1490
rect 4216 1632 4250 1666
rect 4299 1704 4333 1738
rect 4299 1632 4333 1666
rect 4565 1704 4599 1738
rect 4032 1528 4066 1562
rect 4032 1456 4066 1490
rect 4565 1632 4599 1666
rect 4738 1704 4772 1738
rect 5005 1706 5039 1740
rect 5081 1706 5115 1740
rect 5157 1706 5191 1740
rect 5393 1706 5427 1740
rect 5468 1706 5502 1740
rect 5542 1706 5576 1740
rect 4738 1632 4772 1666
rect 5127 1629 5161 1663
rect 5212 1629 5246 1663
rect 5297 1629 5331 1663
rect 5381 1629 5415 1663
rect 5465 1629 5499 1663
rect 4384 1528 4418 1562
rect 4384 1456 4418 1490
rect 4827 1502 4861 1536
rect 3020 1172 3054 1198
rect 3020 1164 3054 1172
rect 3020 1092 3054 1126
rect 4827 1430 4861 1464
rect 5779 555 5813 589
rect 5779 483 5813 517
rect 5867 391 5901 425
rect 5867 319 5901 353
rect 5960 388 5994 422
rect 5960 316 5994 350
rect 2272 23 2288 57
rect 2288 23 2306 57
rect 2345 23 2357 57
rect 2357 23 2379 57
rect 2418 23 2426 57
rect 2426 23 2452 57
rect 2491 23 2495 57
rect 2495 23 2525 57
rect 2564 23 2598 57
rect 2637 23 2667 57
rect 2667 23 2671 57
rect 2710 23 2736 57
rect 2736 23 2744 57
rect 2783 23 2805 57
rect 2805 23 2817 57
rect 2856 23 2874 57
rect 2874 23 2890 57
rect 2928 23 2943 57
rect 2943 23 2962 57
rect 3000 23 3012 57
rect 3012 23 3034 57
rect 3072 23 3081 57
rect 3081 23 3106 57
rect 3144 23 3150 57
rect 3150 23 3178 57
rect 3216 23 3219 57
rect 3219 23 3250 57
rect 3288 23 3322 57
rect 3360 23 3391 57
rect 3391 23 3394 57
rect 3432 23 3459 57
rect 3459 23 3466 57
rect 3504 23 3527 57
rect 3527 23 3538 57
rect 3576 23 3595 57
rect 3595 23 3610 57
rect 3648 23 3663 57
rect 3663 23 3682 57
rect 3720 23 3731 57
rect 3731 23 3754 57
rect 3792 23 3799 57
rect 3799 23 3826 57
rect 3864 23 3867 57
rect 3867 23 3898 57
rect 3936 23 3969 57
rect 3969 23 3970 57
rect 4008 23 4037 57
rect 4037 23 4042 57
rect 4080 23 4105 57
rect 4105 23 4114 57
rect 4152 23 4173 57
rect 4173 23 4186 57
rect 4224 23 4241 57
rect 4241 23 4258 57
rect 4296 23 4309 57
rect 4309 23 4330 57
rect 4368 23 4377 57
rect 4377 23 4402 57
rect 4440 23 4445 57
rect 4445 23 4474 57
rect 4512 23 4513 57
rect 4513 23 4546 57
rect 4584 23 4615 57
rect 4615 23 4618 57
rect 4656 23 4683 57
rect 4683 23 4690 57
rect 4728 23 4751 57
rect 4751 23 4762 57
rect 4800 23 4819 57
rect 4819 23 4834 57
rect 4872 23 4887 57
rect 4887 23 4906 57
rect 4944 23 4955 57
rect 4955 23 4978 57
rect 5016 23 5023 57
rect 5023 23 5050 57
<< metal1 >>
rect 2148 2046 2338 2050
rect 4216 2046 4416 2050
rect 2148 2044 5153 2046
rect 2148 1992 2149 2044
rect 2201 2034 2217 2044
rect 2269 2034 2285 2044
rect 2337 2034 4216 2044
rect 4268 2034 4290 2044
rect 4342 2034 4364 2044
rect 4416 2040 5153 2044
rect 4416 2034 5656 2040
rect 2201 2000 2211 2034
rect 2269 2000 2284 2034
rect 2337 2000 2357 2034
rect 2391 2000 2430 2034
rect 2464 2000 2503 2034
rect 2537 2000 2576 2034
rect 2610 2000 2649 2034
rect 2683 2000 2722 2034
rect 2756 2000 2795 2034
rect 2829 2000 2868 2034
rect 2902 2000 2941 2034
rect 2975 2000 3014 2034
rect 3048 2000 3087 2034
rect 3121 2000 3160 2034
rect 3194 2000 3233 2034
rect 3267 2000 3306 2034
rect 3340 2000 3378 2034
rect 3412 2000 3450 2034
rect 3484 2000 3522 2034
rect 3556 2000 3594 2034
rect 3628 2000 3666 2034
rect 3700 2000 3738 2034
rect 3772 2000 3810 2034
rect 3844 2000 3882 2034
rect 3916 2000 3954 2034
rect 3988 2000 4026 2034
rect 4060 2000 4098 2034
rect 4132 2000 4170 2034
rect 4204 2000 4216 2034
rect 4276 2000 4290 2034
rect 4348 2000 4364 2034
rect 4420 2000 4458 2034
rect 4492 2000 4530 2034
rect 4564 2000 4602 2034
rect 4636 2000 4674 2034
rect 4708 2000 4746 2034
rect 4780 2000 4818 2034
rect 4852 2000 4890 2034
rect 4924 2000 4962 2034
rect 4996 2000 5034 2034
rect 5068 2000 5106 2034
rect 5140 2000 5178 2034
rect 5212 2000 5250 2034
rect 5284 2000 5322 2034
rect 5356 2000 5394 2034
rect 5428 2000 5466 2034
rect 5500 2000 5538 2034
rect 5572 2000 5610 2034
rect 5644 2000 5656 2034
rect 2201 1992 2217 2000
rect 2269 1992 2285 2000
rect 2337 1992 4216 2000
rect 4268 1992 4290 2000
rect 4342 1992 4364 2000
rect 4416 1994 5656 2000
rect 4416 1992 5153 1994
rect 2148 1967 5153 1992
rect 2148 1915 2149 1967
rect 2201 1949 2217 1967
rect 2201 1915 2203 1949
rect 2269 1915 2285 1967
rect 2337 1949 4216 1967
rect 2337 1915 2555 1949
rect 2589 1915 2668 1949
rect 2702 1915 3020 1949
rect 3054 1915 4216 1949
rect 4268 1915 4290 1967
rect 4342 1915 4364 1967
rect 4416 1915 5153 1967
rect 2148 1889 5153 1915
rect 2148 1837 2149 1889
rect 2201 1877 2217 1889
rect 2201 1843 2203 1877
rect 2201 1837 2217 1843
rect 2269 1837 2285 1889
rect 2337 1877 4216 1889
rect 2337 1843 2555 1877
rect 2589 1843 2668 1877
rect 2702 1843 3020 1877
rect 3054 1843 4216 1877
rect 2337 1837 4216 1843
rect 4268 1837 4290 1889
rect 4342 1837 4364 1889
rect 4416 1837 5153 1889
rect 2148 1831 5153 1837
rect 4867 1830 4892 1831
rect 1673 1772 3531 1803
tri 1949 1670 2020 1741 se
rect 2020 1740 2512 1741
rect 2020 1734 2518 1740
rect 2020 1689 2466 1734
rect 2928 1731 3236 1743
rect 2020 1670 2023 1689
tri 2023 1670 2042 1689 nw
rect 1454 1618 1460 1670
rect 1512 1618 1524 1670
rect 1576 1618 1971 1670
tri 1971 1618 2023 1670 nw
rect 2466 1668 2518 1682
rect 1454 1586 1500 1618
tri 2094 1595 2160 1661 se
rect 2160 1655 2354 1661
rect 2160 1621 2236 1655
rect 2270 1621 2308 1655
rect 2342 1621 2354 1655
rect 2160 1615 2354 1621
tri 2588 1639 2654 1705 se
rect 2654 1699 2817 1705
rect 2654 1665 2699 1699
rect 2733 1665 2771 1699
rect 2805 1665 2817 1699
rect 2654 1659 2817 1665
rect 2928 1697 2934 1731
rect 2968 1697 3196 1731
rect 3230 1697 3236 1731
rect 2928 1659 3236 1697
tri 3292 1676 3388 1772 ne
rect 3388 1743 3531 1772
tri 3531 1743 3591 1803 sw
rect 3388 1737 3754 1743
rect 3388 1731 3702 1737
rect 3388 1697 3482 1731
rect 3516 1697 3702 1731
rect 3388 1685 3702 1697
tri 2654 1639 2674 1659 nw
tri 2160 1595 2180 1615 nw
rect 2466 1610 2518 1616
tri 2576 1627 2588 1639 se
rect 2588 1627 2622 1639
rect 1454 1552 1460 1586
rect 1494 1552 1500 1586
rect 1454 1540 1500 1552
tri 2041 1542 2094 1595 se
rect 2094 1542 2107 1595
tri 2107 1542 2160 1595 nw
tri 1787 1373 1821 1407 se
rect 1821 1373 1873 1452
tri 1873 1373 1907 1407 sw
rect 558 1371 776 1373
rect 558 1319 564 1371
rect 616 1319 641 1371
rect 693 1319 718 1371
rect 770 1319 776 1371
rect 558 1299 776 1319
rect 558 1247 564 1299
rect 616 1247 641 1299
rect 693 1247 718 1299
rect 770 1247 776 1299
rect 558 1227 776 1247
rect 558 1175 564 1227
rect 616 1175 641 1227
rect 693 1175 718 1227
rect 770 1175 776 1227
rect 558 1174 776 1175
rect 1826 1367 1983 1373
rect 1878 1315 1930 1367
rect 1982 1315 1983 1367
rect 1826 1300 1983 1315
rect 1878 1248 1930 1300
rect 1982 1248 1983 1300
rect 1826 1232 1983 1248
rect 1878 1180 1930 1232
rect 1982 1180 1983 1232
rect 1826 1174 1983 1180
rect 335 732 387 738
tri 301 658 335 692 ne
rect 1876 727 1983 777
rect 1887 725 1983 727
rect 335 668 387 680
rect 335 610 387 616
rect 1665 406 1793 536
rect 1872 420 1963 529
rect 1694 377 1983 378
rect 1694 325 1700 377
rect 1752 325 1812 377
rect 1864 325 1925 377
rect 1977 325 1983 377
rect 1694 303 1983 325
rect 1694 251 1700 303
rect 1752 251 1812 303
rect 1864 251 1925 303
rect 1977 251 1983 303
rect 1694 229 1983 251
rect 1694 177 1700 229
rect 1752 177 1812 229
rect 1864 177 1925 229
rect 1977 177 1983 229
rect 1694 176 1983 177
tri 1999 67 2041 109 se
rect 2041 87 2093 1542
tri 2093 1528 2107 1542 nw
rect 2200 1410 2246 1422
rect 2200 1376 2206 1410
rect 2240 1391 2246 1410
tri 2535 1391 2576 1432 se
rect 2576 1412 2622 1627
tri 2622 1607 2654 1639 nw
rect 2928 1625 2934 1659
rect 2968 1625 3196 1659
rect 3230 1625 3236 1659
rect 2928 1613 3236 1625
rect 3388 1673 3754 1685
rect 3388 1659 3702 1673
rect 3388 1625 3482 1659
rect 3516 1625 3702 1659
rect 3388 1621 3702 1625
rect 3388 1613 3754 1621
rect 4210 1738 4256 1750
rect 4210 1704 4216 1738
rect 4250 1704 4256 1738
rect 4210 1666 4256 1704
rect 4210 1632 4216 1666
rect 4250 1632 4256 1666
rect 4210 1620 4256 1632
rect 4293 1738 4778 1750
rect 4293 1704 4299 1738
rect 4333 1704 4565 1738
rect 4599 1704 4738 1738
rect 4772 1704 4778 1738
rect 4293 1666 4778 1704
tri 4891 1680 4957 1746 se
rect 4957 1740 5588 1746
rect 4957 1706 5005 1740
rect 5039 1706 5081 1740
rect 5115 1706 5157 1740
rect 5191 1706 5393 1740
rect 5427 1706 5468 1740
rect 5502 1706 5542 1740
rect 5576 1706 5588 1740
rect 4957 1700 5588 1706
tri 4957 1680 4977 1700 nw
rect 4293 1632 4299 1666
rect 4333 1632 4565 1666
rect 4599 1632 4738 1666
rect 4772 1632 4778 1666
rect 4293 1620 4778 1632
tri 4825 1614 4891 1680 se
tri 4891 1614 4957 1680 nw
rect 5115 1663 5511 1669
rect 5167 1629 5212 1663
rect 5246 1629 5297 1663
rect 5331 1629 5381 1663
rect 5415 1629 5465 1663
rect 5499 1629 5511 1663
tri 4821 1610 4825 1614 se
rect 4825 1610 4867 1614
rect 3391 1562 4424 1574
rect 3102 1554 3303 1555
rect 3102 1548 3354 1554
rect 3102 1543 3302 1548
rect 2576 1391 2601 1412
tri 2601 1391 2622 1412 nw
rect 2662 1527 2708 1539
rect 2662 1493 2668 1527
rect 2702 1493 2708 1527
rect 2662 1455 2708 1493
rect 2662 1421 2668 1455
rect 2702 1421 2708 1455
rect 3102 1509 3108 1543
rect 3142 1509 3302 1543
rect 3102 1496 3302 1509
rect 3102 1484 3354 1496
rect 3102 1471 3302 1484
rect 3102 1437 3108 1471
rect 3142 1437 3302 1471
rect 3102 1432 3302 1437
rect 3391 1528 3397 1562
rect 3431 1528 3573 1562
rect 3607 1528 4032 1562
rect 4066 1528 4384 1562
rect 4418 1528 4424 1562
rect 3391 1490 4424 1528
rect 3391 1456 3397 1490
rect 3431 1456 3573 1490
rect 3607 1456 4032 1490
rect 4066 1456 4384 1490
rect 4418 1456 4424 1490
rect 3391 1444 4424 1456
rect 4821 1536 4867 1610
tri 4867 1590 4891 1614 nw
rect 5167 1623 5511 1629
rect 5115 1599 5167 1611
rect 5115 1541 5167 1547
rect 4821 1502 4827 1536
rect 4861 1502 4867 1536
rect 4821 1464 4867 1502
rect 3102 1426 3354 1432
rect 4821 1430 4827 1464
rect 4861 1430 4867 1464
rect 3102 1425 3303 1426
rect 2662 1409 2708 1421
rect 4821 1416 4867 1430
rect 2240 1376 2555 1391
rect 2200 1345 2555 1376
tri 2555 1345 2601 1391 nw
tri 3490 1350 3556 1416 se
rect 3556 1383 4867 1416
rect 3556 1370 4854 1383
tri 4854 1370 4867 1383 nw
tri 3556 1350 3576 1370 nw
rect 2200 1338 2246 1345
rect 2200 1304 2206 1338
rect 2240 1304 2246 1338
tri 3453 1313 3490 1350 se
rect 3490 1313 3519 1350
tri 3519 1313 3556 1350 nw
rect 2200 1292 2246 1304
rect 2400 1261 2406 1313
rect 2458 1261 2470 1313
rect 2522 1267 3473 1313
tri 3473 1267 3519 1313 nw
rect 2522 1261 2528 1267
rect 3686 1266 3692 1318
rect 3744 1266 3756 1318
rect 3808 1266 5800 1318
rect 5852 1266 5864 1318
rect 5916 1266 5922 1318
rect 2191 1210 2601 1211
rect 2635 1210 3285 1211
rect 2191 1205 5329 1210
rect 2191 1198 2636 1205
rect 2191 1164 2555 1198
rect 2589 1164 2636 1198
rect 2191 1153 2636 1164
rect 2688 1153 2710 1205
rect 2762 1153 2784 1205
rect 2836 1198 5329 1205
rect 2836 1164 3020 1198
rect 3054 1164 5329 1198
rect 2836 1153 5329 1164
rect 2191 1133 5329 1153
rect 2191 1126 2636 1133
rect 2191 1092 2555 1126
rect 2589 1092 2636 1126
rect 2191 1081 2636 1092
rect 2688 1081 2710 1133
rect 2762 1081 2784 1133
rect 2836 1126 5329 1133
rect 2836 1092 3020 1126
rect 3054 1092 5329 1126
rect 2836 1081 5329 1092
rect 2191 1061 5329 1081
rect 2191 1009 2636 1061
rect 2688 1009 2710 1061
rect 2762 1009 2784 1061
rect 2836 1049 5329 1061
rect 2836 1009 6089 1049
rect 2191 1008 6089 1009
rect 2635 989 2837 1008
rect 2635 937 2636 989
rect 2688 937 2710 989
rect 2762 937 2784 989
rect 2836 937 2837 989
rect 2635 917 2837 937
rect 2635 865 2636 917
rect 2688 865 2710 917
rect 2762 865 2784 917
rect 2836 865 2837 917
rect 2635 859 2837 865
rect 4929 847 6089 1008
rect 5773 595 5825 601
rect 3302 565 5119 571
rect 3354 525 5119 565
rect 3302 501 3354 513
rect 3086 388 3143 459
tri 5089 495 5119 525 ne
tri 5119 495 5195 571 sw
rect 5825 544 5947 590
tri 5947 544 5993 590 sw
rect 5773 529 5825 543
tri 5927 517 5954 544 ne
rect 5954 537 5993 544
tri 5993 537 6000 544 sw
rect 3302 443 3354 449
tri 5119 419 5195 495 ne
tri 5195 437 5253 495 sw
rect 5773 471 5825 477
rect 5195 425 5907 437
rect 5195 419 5867 425
rect 3297 349 5045 401
rect 5097 349 5109 401
rect 5161 349 5167 401
tri 5195 380 5234 419 ne
rect 5234 391 5867 419
rect 5901 391 5907 425
rect 5234 353 5907 391
rect 5234 319 5867 353
rect 5901 319 5907 353
rect 5234 307 5907 319
rect 5954 422 6000 537
rect 5954 388 5960 422
rect 5994 388 6000 422
rect 5954 350 6000 388
rect 5954 316 5960 350
rect 5994 316 6000 350
rect 5954 304 6000 316
rect 2041 67 2069 87
rect 335 15 341 67
rect 393 15 405 67
rect 457 63 2069 67
tri 2069 63 2093 87 nw
rect 4216 221 4416 227
rect 4268 169 4290 221
rect 4342 169 4364 221
rect 4216 146 4416 169
rect 4268 94 4290 146
rect 4342 94 4364 146
rect 4216 70 4416 94
rect 457 15 2021 63
tri 2021 15 2069 63 nw
rect 2260 57 4216 63
rect 2260 23 2272 57
rect 2306 23 2345 57
rect 2379 23 2418 57
rect 2452 23 2491 57
rect 2525 23 2564 57
rect 2598 23 2637 57
rect 2671 23 2710 57
rect 2744 23 2783 57
rect 2817 23 2856 57
rect 2890 23 2928 57
rect 2962 23 3000 57
rect 3034 23 3072 57
rect 3106 23 3144 57
rect 3178 23 3216 57
rect 3250 23 3288 57
rect 3322 23 3360 57
rect 3394 23 3432 57
rect 3466 23 3504 57
rect 3538 23 3576 57
rect 3610 23 3648 57
rect 3682 23 3720 57
rect 3754 23 3792 57
rect 3826 23 3864 57
rect 3898 23 3936 57
rect 3970 23 4008 57
rect 4042 23 4080 57
rect 4114 23 4152 57
rect 4186 23 4216 57
rect 2260 18 4216 23
rect 4268 18 4290 70
rect 4342 18 4364 70
rect 4416 57 5062 63
rect 4416 23 4440 57
rect 4474 23 4512 57
rect 4546 23 4584 57
rect 4618 23 4656 57
rect 4690 23 4728 57
rect 4762 23 4800 57
rect 4834 23 4872 57
rect 4906 23 4944 57
rect 4978 23 5016 57
rect 5050 23 5062 57
rect 4416 18 5062 23
rect 2260 17 5062 18
rect 4216 12 4416 17
rect 5073 13 6037 227
<< via1 >>
rect 2149 1992 2201 2044
rect 2217 2034 2269 2044
rect 2285 2034 2337 2044
rect 4216 2034 4268 2044
rect 4290 2034 4342 2044
rect 4364 2034 4416 2044
rect 2217 2000 2245 2034
rect 2245 2000 2269 2034
rect 2285 2000 2318 2034
rect 2318 2000 2337 2034
rect 4216 2000 4242 2034
rect 4242 2000 4268 2034
rect 4290 2000 4314 2034
rect 4314 2000 4342 2034
rect 4364 2000 4386 2034
rect 4386 2000 4416 2034
rect 2217 1992 2269 2000
rect 2285 1992 2337 2000
rect 4216 1992 4268 2000
rect 4290 1992 4342 2000
rect 4364 1992 4416 2000
rect 2149 1915 2201 1967
rect 2217 1949 2269 1967
rect 2217 1915 2237 1949
rect 2237 1915 2269 1949
rect 2285 1915 2337 1967
rect 4216 1915 4268 1967
rect 4290 1915 4342 1967
rect 4364 1915 4416 1967
rect 2149 1837 2201 1889
rect 2217 1877 2269 1889
rect 2217 1843 2237 1877
rect 2237 1843 2269 1877
rect 2217 1837 2269 1843
rect 2285 1837 2337 1889
rect 4216 1837 4268 1889
rect 4290 1837 4342 1889
rect 4364 1837 4416 1889
rect 2466 1729 2518 1734
rect 2466 1695 2472 1729
rect 2472 1695 2506 1729
rect 2506 1695 2518 1729
rect 2466 1682 2518 1695
rect 1460 1658 1512 1670
rect 1460 1624 1494 1658
rect 1494 1624 1512 1658
rect 1460 1618 1512 1624
rect 1524 1618 1576 1670
rect 2466 1657 2518 1668
rect 2466 1623 2472 1657
rect 2472 1623 2506 1657
rect 2506 1623 2518 1657
rect 3702 1685 3754 1737
rect 2466 1616 2518 1623
rect 564 1319 616 1371
rect 641 1319 693 1371
rect 718 1319 770 1371
rect 564 1247 616 1299
rect 641 1247 693 1299
rect 718 1247 770 1299
rect 564 1175 616 1227
rect 641 1175 693 1227
rect 718 1175 770 1227
rect 1826 1315 1878 1367
rect 1930 1315 1982 1367
rect 1826 1248 1878 1300
rect 1930 1248 1982 1300
rect 1826 1180 1878 1232
rect 1930 1180 1982 1232
rect 335 680 387 732
rect 335 616 387 668
rect 1700 325 1752 377
rect 1812 325 1864 377
rect 1925 325 1977 377
rect 1700 251 1752 303
rect 1812 251 1864 303
rect 1925 251 1977 303
rect 1700 177 1752 229
rect 1812 177 1864 229
rect 1925 177 1977 229
rect 3702 1621 3754 1673
rect 5115 1629 5127 1663
rect 5127 1629 5161 1663
rect 5161 1629 5167 1663
rect 3302 1496 3354 1548
rect 3302 1432 3354 1484
rect 5115 1611 5167 1629
rect 5115 1547 5167 1599
rect 2406 1261 2458 1313
rect 2470 1261 2522 1313
rect 3692 1266 3744 1318
rect 3756 1266 3808 1318
rect 5800 1266 5852 1318
rect 5864 1266 5916 1318
rect 2636 1153 2688 1205
rect 2710 1153 2762 1205
rect 2784 1153 2836 1205
rect 2636 1081 2688 1133
rect 2710 1081 2762 1133
rect 2784 1081 2836 1133
rect 2636 1009 2688 1061
rect 2710 1009 2762 1061
rect 2784 1009 2836 1061
rect 2636 937 2688 989
rect 2710 937 2762 989
rect 2784 937 2836 989
rect 2636 865 2688 917
rect 2710 865 2762 917
rect 2784 865 2836 917
rect 5773 589 5825 595
rect 3302 513 3354 565
rect 3302 449 3354 501
rect 5773 555 5779 589
rect 5779 555 5813 589
rect 5813 555 5825 589
rect 5773 543 5825 555
rect 5773 517 5825 529
rect 5773 483 5779 517
rect 5779 483 5813 517
rect 5813 483 5825 517
rect 5773 477 5825 483
rect 5045 349 5097 401
rect 5109 349 5161 401
rect 341 15 393 67
rect 405 15 457 67
rect 4216 169 4268 221
rect 4290 169 4342 221
rect 4364 169 4416 221
rect 4216 94 4268 146
rect 4290 94 4342 146
rect 4364 94 4416 146
rect 4216 57 4268 70
rect 4216 23 4224 57
rect 4224 23 4258 57
rect 4258 23 4268 57
rect 4216 18 4268 23
rect 4290 57 4342 70
rect 4290 23 4296 57
rect 4296 23 4330 57
rect 4330 23 4342 57
rect 4290 18 4342 23
rect 4364 57 4416 70
rect 4364 23 4368 57
rect 4368 23 4402 57
rect 4402 23 4416 57
rect 4364 18 4416 23
<< metal2 >>
rect 2148 2044 2339 2050
rect 2148 1992 2149 2044
rect 2201 1992 2217 2044
rect 2269 1992 2285 2044
rect 2337 1992 2339 2044
rect 2148 1967 2339 1992
rect 2148 1915 2149 1967
rect 2201 1915 2217 1967
rect 2269 1915 2285 1967
rect 2337 1915 2339 1967
rect 2148 1889 2339 1915
rect 2148 1837 2149 1889
rect 2201 1837 2217 1889
rect 2269 1837 2285 1889
rect 2337 1837 2339 1889
rect 1454 1618 1460 1670
rect 1512 1618 1524 1670
rect 1576 1618 1582 1670
tri 2114 1373 2148 1407 se
rect 2148 1373 2339 1837
rect 2466 1734 2518 1740
rect 2466 1668 2518 1682
rect 558 1371 776 1372
rect 558 1319 564 1371
rect 616 1319 641 1371
rect 693 1319 718 1371
rect 770 1319 776 1371
rect 558 1299 776 1319
rect 558 1247 564 1299
rect 616 1247 641 1299
rect 693 1247 718 1299
rect 770 1247 776 1299
rect 558 1227 776 1247
rect 558 1175 564 1227
rect 616 1175 641 1227
rect 693 1175 718 1227
rect 770 1175 776 1227
rect 558 1174 776 1175
rect 1826 1367 2339 1373
rect 1878 1315 1930 1367
rect 1982 1315 2339 1367
rect 1826 1300 2339 1315
rect 1878 1248 1930 1300
rect 1982 1248 2339 1300
tri 2400 1313 2466 1379 se
rect 2466 1313 2518 1616
tri 2518 1313 2528 1323 sw
rect 2400 1261 2406 1313
rect 2458 1261 2470 1313
rect 2522 1261 2528 1313
rect 1826 1232 2339 1248
rect 1878 1180 1930 1232
rect 1982 1180 2339 1232
rect 1826 1174 2339 1180
rect 2635 1205 2837 2077
rect 4216 2044 4416 2050
rect 4268 1992 4290 2044
rect 4342 1992 4364 2044
rect 4216 1967 4416 1992
rect 4268 1915 4290 1967
rect 4342 1915 4364 1967
rect 4216 1889 4416 1915
rect 4268 1837 4290 1889
rect 4342 1837 4364 1889
rect 3702 1737 3754 1743
rect 3702 1673 3754 1685
rect 2635 1153 2636 1205
rect 2688 1153 2710 1205
rect 2762 1153 2784 1205
rect 2836 1153 2837 1205
rect 2635 1133 2837 1153
rect 2635 1081 2636 1133
rect 2688 1081 2710 1133
rect 2762 1081 2784 1133
rect 2836 1081 2837 1133
rect 2635 1061 2837 1081
rect 2635 1009 2636 1061
rect 2688 1009 2710 1061
rect 2762 1009 2784 1061
rect 2836 1009 2837 1061
rect 2635 989 2837 1009
rect 2635 937 2636 989
rect 2688 937 2710 989
rect 2762 937 2784 989
rect 2836 937 2837 989
rect 2635 917 2837 937
rect 2635 865 2636 917
rect 2688 865 2710 917
rect 2762 865 2784 917
rect 2836 865 2837 917
rect 335 732 387 738
rect 335 668 387 680
rect 335 67 387 616
tri 2427 378 2635 586 se
rect 2635 378 2837 865
rect 3302 1548 3354 1554
rect 3302 1484 3354 1496
rect 3302 565 3354 1432
rect 3702 1318 3754 1621
rect 3686 1266 3692 1318
rect 3744 1266 3756 1318
rect 3808 1266 3814 1318
rect 3302 501 3354 513
rect 3302 443 3354 449
rect 1694 377 2837 378
rect 1694 325 1700 377
rect 1752 325 1812 377
rect 1864 325 1925 377
rect 1977 325 2837 377
rect 1694 303 2837 325
rect 1694 251 1700 303
rect 1752 251 1812 303
rect 1864 251 1925 303
rect 1977 294 2837 303
rect 1977 251 2719 294
rect 1694 229 2719 251
rect 1694 177 1700 229
rect 1752 177 1812 229
rect 1864 177 1925 229
rect 1977 177 2719 229
rect 1694 176 2719 177
tri 2719 176 2837 294 nw
rect 4216 221 4416 1837
rect 5115 1663 5167 1669
rect 5115 1599 5167 1611
tri 5039 401 5115 477 se
rect 5115 401 5167 1547
rect 5794 1266 5800 1318
rect 5852 1266 5864 1318
rect 5916 1266 5922 1318
tri 5773 964 5819 1010 se
rect 5819 988 5871 1266
rect 5819 964 5825 988
rect 5773 595 5825 964
tri 5825 942 5871 988 nw
rect 5773 529 5825 543
rect 5773 471 5825 477
rect 5039 349 5045 401
rect 5097 349 5109 401
rect 5161 349 5167 401
rect 4268 169 4290 221
rect 4342 169 4364 221
rect 4216 146 4416 169
tri 387 67 421 101 sw
rect 4268 94 4290 146
rect 4342 94 4364 146
rect 4216 70 4416 94
rect 335 15 341 67
rect 393 15 405 67
rect 457 15 463 67
rect 4268 18 4290 70
rect 4342 18 4364 70
rect 4216 12 4416 18
use sky130_fd_io__enh_nand2_1_i2c_fix  sky130_fd_io__enh_nand2_1_i2c_fix_0
timestamp 1676037725
transform 1 0 3232 0 -1 2070
box -42 24 710 1116
use sky130_fd_io__enh_nand2_1_sp  sky130_fd_io__enh_nand2_1_sp_0
timestamp 1676037725
transform -1 0 4583 0 -1 2069
box -42 24 710 1116
use sky130_fd_io__enh_nor2_x1  sky130_fd_io__enh_nor2_x1_0
timestamp 1676037725
transform 1 0 5611 0 1 -12
box 0 24 534 1116
use sky130_fd_io__enh_nor2_x1  sky130_fd_io__enh_nor2_x1_1
timestamp 1676037725
transform 1 0 4401 0 -1 2069
box 0 24 534 1116
use sky130_fd_io__gpio_ovtv2_ctl_ls_i2c_fix_1  sky130_fd_io__gpio_ovtv2_ctl_ls_i2c_fix_1_0
timestamp 1676037725
transform 1 0 -94 0 1 52
box -71 10 2077 2019
use sky130_fd_io__hvsbt_inv_x1  sky130_fd_io__hvsbt_inv_x1_0
timestamp 1676037725
transform 1 0 2946 0 -1 2070
box 107 226 240 873
use sky130_fd_io__hvsbt_nor  sky130_fd_io__hvsbt_nor_0
timestamp 1676037725
transform -1 0 3128 0 -1 2070
box 107 226 460 873
use sky130_fd_io__hvsbt_nor  sky130_fd_io__hvsbt_nor_1
timestamp 1676037725
transform -1 0 2663 0 -1 2070
box 107 226 460 873
use sky130_fd_io__nand2_2_enhpath  sky130_fd_io__nand2_2_enhpath_0
timestamp 1676037725
transform 1 0 4863 0 -1 2069
box 0 24 886 1116
use sky130_fd_io__nor2_4_enhpath  sky130_fd_io__nor2_4_enhpath_0
timestamp 1676037725
transform -1 0 8072 0 1 -1097
box 2931 1109 5929 2209
<< labels >>
flabel metal1 s 4182 1495 4271 1550 3 FreeSans 520 0 0 0 ENABLE_H
port 2 nsew
flabel metal1 s 4218 1664 4245 1709 3 FreeSans 520 0 0 0 HLD_H_N
port 3 nsew
flabel metal1 s 1876 727 1919 777 3 FreeSans 520 0 0 0 HLD_OVR
port 4 nsew
flabel metal1 s 3219 1051 3357 1148 3 FreeSans 520 0 0 0 VCC_IO
port 5 nsew
flabel metal1 s 2941 1886 3057 2029 3 FreeSans 520 0 0 0 VGND
port 6 nsew
flabel metal1 s 1872 420 1963 529 3 FreeSans 520 0 0 0 VPWR
port 7 nsew
flabel metal1 s 2665 1430 2703 1491 3 FreeSans 520 0 0 0 HLD_I_OVR_H
port 8 nsew
flabel metal1 s 3205 1469 3260 1521 3 FreeSans 520 0 0 0 OD_I_H_N
port 9 nsew
flabel metal1 s 3086 388 3143 459 3 FreeSans 520 180 0 0 HLD_I_H_N
port 10 nsew
flabel metal2 s 4268 1610 4366 1714 0 FreeSans 200 0 0 0 VGND
port 6 nsew
flabel metal2 s 2702 1610 2800 1714 0 FreeSans 200 0 0 0 VCC_IO
port 5 nsew
<< properties >>
string GDS_END 31922076
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 31887442
<< end >>
