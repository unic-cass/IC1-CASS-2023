magic
tech sky130B
magscale 1 2
timestamp 1676037725
<< nwell >>
rect -36 679 404 1471
<< locali >>
rect 0 1397 368 1431
rect 64 658 98 724
rect 179 674 213 708
rect 0 -17 368 17
use pinv_3  pinv_3_0
timestamp 1676037725
transform 1 0 0 0 1 0
box -36 -17 404 1471
<< labels >>
rlabel locali s 196 691 196 691 4 Z
port 2 nsew
rlabel locali s 81 691 81 691 4 A
port 1 nsew
rlabel locali s 184 1414 184 1414 4 vdd
port 3 nsew
rlabel locali s 184 0 184 0 4 gnd
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 368 1414
string GDS_END 3593902
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sram_1rw1r_32_256_8_sky130.gds
string GDS_START 3593064
<< end >>
