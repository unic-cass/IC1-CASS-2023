magic
tech sky130A
magscale 1 2
timestamp 1676037725
<< nwell >>
rect -38 261 2062 582
<< pwell >>
rect 1 21 2023 203
rect 29 -17 63 21
<< scnmos >>
rect 79 47 109 177
rect 163 47 193 177
rect 247 47 277 177
rect 331 47 361 177
rect 545 47 575 177
rect 629 47 659 177
rect 713 47 743 177
rect 797 47 827 177
rect 881 47 911 177
rect 965 47 995 177
rect 1049 47 1079 177
rect 1133 47 1163 177
rect 1321 47 1351 177
rect 1405 47 1435 177
rect 1489 47 1519 177
rect 1573 47 1603 177
rect 1657 47 1687 177
rect 1741 47 1771 177
rect 1825 47 1855 177
rect 1909 47 1939 177
<< scpmoshvt >>
rect 79 297 109 497
rect 163 297 193 497
rect 247 297 277 497
rect 331 297 361 497
rect 477 297 507 497
rect 629 297 659 497
rect 713 297 743 497
rect 797 297 827 497
rect 900 297 930 497
rect 984 297 1014 497
rect 1068 297 1098 497
rect 1233 297 1263 497
rect 1321 297 1351 497
rect 1405 297 1435 497
rect 1489 297 1519 497
rect 1573 297 1603 497
rect 1657 297 1687 497
rect 1741 297 1771 497
rect 1825 297 1855 497
rect 1909 297 1939 497
<< ndiff >>
rect 27 93 79 177
rect 27 59 35 93
rect 69 59 79 93
rect 27 47 79 59
rect 109 101 163 177
rect 109 67 119 101
rect 153 67 163 101
rect 109 47 163 67
rect 193 93 247 177
rect 193 59 203 93
rect 237 59 247 93
rect 193 47 247 59
rect 277 109 331 177
rect 277 75 287 109
rect 321 75 331 109
rect 277 47 331 75
rect 361 93 413 177
rect 361 59 371 93
rect 405 59 413 93
rect 361 47 413 59
rect 493 93 545 177
rect 493 59 501 93
rect 535 59 545 93
rect 493 47 545 59
rect 575 161 629 177
rect 575 127 585 161
rect 619 127 629 161
rect 575 47 629 127
rect 659 93 713 177
rect 659 59 669 93
rect 703 59 713 93
rect 659 47 713 59
rect 743 161 797 177
rect 743 127 753 161
rect 787 127 797 161
rect 743 47 797 127
rect 827 93 881 177
rect 827 59 837 93
rect 871 59 881 93
rect 827 47 881 59
rect 911 161 965 177
rect 911 127 921 161
rect 955 127 965 161
rect 911 47 965 127
rect 995 93 1049 177
rect 995 59 1005 93
rect 1039 59 1049 93
rect 995 47 1049 59
rect 1079 161 1133 177
rect 1079 127 1089 161
rect 1123 127 1133 161
rect 1079 47 1133 127
rect 1163 93 1215 177
rect 1163 59 1173 93
rect 1207 59 1215 93
rect 1163 47 1215 59
rect 1269 93 1321 177
rect 1269 59 1277 93
rect 1311 59 1321 93
rect 1269 47 1321 59
rect 1351 161 1405 177
rect 1351 127 1361 161
rect 1395 127 1405 161
rect 1351 47 1405 127
rect 1435 93 1489 177
rect 1435 59 1445 93
rect 1479 59 1489 93
rect 1435 47 1489 59
rect 1519 161 1573 177
rect 1519 127 1529 161
rect 1563 127 1573 161
rect 1519 47 1573 127
rect 1603 101 1657 177
rect 1603 67 1613 101
rect 1647 67 1657 101
rect 1603 47 1657 67
rect 1687 93 1741 177
rect 1687 59 1697 93
rect 1731 59 1741 93
rect 1687 47 1741 59
rect 1771 101 1825 177
rect 1771 67 1781 101
rect 1815 67 1825 101
rect 1771 47 1825 67
rect 1855 93 1909 177
rect 1855 59 1865 93
rect 1899 59 1909 93
rect 1855 47 1909 59
rect 1939 101 1997 177
rect 1939 67 1949 101
rect 1983 67 1997 101
rect 1939 47 1997 67
<< pdiff >>
rect 27 485 79 497
rect 27 451 35 485
rect 69 451 79 485
rect 27 297 79 451
rect 109 417 163 497
rect 109 383 119 417
rect 153 383 163 417
rect 109 349 163 383
rect 109 315 119 349
rect 153 315 163 349
rect 109 297 163 315
rect 193 485 247 497
rect 193 451 203 485
rect 237 451 247 485
rect 193 297 247 451
rect 277 417 331 497
rect 277 383 287 417
rect 321 383 331 417
rect 277 349 331 383
rect 277 315 287 349
rect 321 315 331 349
rect 277 297 331 315
rect 361 477 477 497
rect 361 443 433 477
rect 467 443 477 477
rect 361 297 477 443
rect 507 485 629 497
rect 507 451 517 485
rect 551 451 585 485
rect 619 451 629 485
rect 507 297 629 451
rect 659 477 713 497
rect 659 443 669 477
rect 703 443 713 477
rect 659 297 713 443
rect 743 485 797 497
rect 743 451 753 485
rect 787 451 797 485
rect 743 417 797 451
rect 743 383 753 417
rect 787 383 797 417
rect 743 297 797 383
rect 827 469 900 497
rect 827 435 837 469
rect 871 435 900 469
rect 827 297 900 435
rect 930 485 984 497
rect 930 451 940 485
rect 974 451 984 485
rect 930 417 984 451
rect 930 383 940 417
rect 974 383 984 417
rect 930 297 984 383
rect 1014 477 1068 497
rect 1014 443 1024 477
rect 1058 443 1068 477
rect 1014 409 1068 443
rect 1014 375 1024 409
rect 1058 375 1068 409
rect 1014 297 1068 375
rect 1098 485 1233 497
rect 1098 383 1115 485
rect 1217 383 1233 485
rect 1098 297 1233 383
rect 1263 477 1321 497
rect 1263 443 1277 477
rect 1311 443 1321 477
rect 1263 409 1321 443
rect 1263 375 1277 409
rect 1311 375 1321 409
rect 1263 297 1321 375
rect 1351 485 1405 497
rect 1351 451 1361 485
rect 1395 451 1405 485
rect 1351 417 1405 451
rect 1351 383 1361 417
rect 1395 383 1405 417
rect 1351 297 1405 383
rect 1435 477 1489 497
rect 1435 443 1445 477
rect 1479 443 1489 477
rect 1435 409 1489 443
rect 1435 375 1445 409
rect 1479 375 1489 409
rect 1435 297 1489 375
rect 1519 485 1573 497
rect 1519 451 1529 485
rect 1563 451 1573 485
rect 1519 297 1573 451
rect 1603 477 1657 497
rect 1603 443 1613 477
rect 1647 443 1657 477
rect 1603 409 1657 443
rect 1603 375 1613 409
rect 1647 375 1657 409
rect 1603 297 1657 375
rect 1687 485 1741 497
rect 1687 451 1697 485
rect 1731 451 1741 485
rect 1687 417 1741 451
rect 1687 383 1697 417
rect 1731 383 1741 417
rect 1687 297 1741 383
rect 1771 477 1825 497
rect 1771 443 1781 477
rect 1815 443 1825 477
rect 1771 409 1825 443
rect 1771 375 1781 409
rect 1815 375 1825 409
rect 1771 297 1825 375
rect 1855 485 1909 497
rect 1855 451 1865 485
rect 1899 451 1909 485
rect 1855 417 1909 451
rect 1855 383 1865 417
rect 1899 383 1909 417
rect 1855 297 1909 383
rect 1939 477 1997 497
rect 1939 443 1955 477
rect 1989 443 1997 477
rect 1939 409 1997 443
rect 1939 375 1955 409
rect 1989 375 1997 409
rect 1939 297 1997 375
<< ndiffc >>
rect 35 59 69 93
rect 119 67 153 101
rect 203 59 237 93
rect 287 75 321 109
rect 371 59 405 93
rect 501 59 535 93
rect 585 127 619 161
rect 669 59 703 93
rect 753 127 787 161
rect 837 59 871 93
rect 921 127 955 161
rect 1005 59 1039 93
rect 1089 127 1123 161
rect 1173 59 1207 93
rect 1277 59 1311 93
rect 1361 127 1395 161
rect 1445 59 1479 93
rect 1529 127 1563 161
rect 1613 67 1647 101
rect 1697 59 1731 93
rect 1781 67 1815 101
rect 1865 59 1899 93
rect 1949 67 1983 101
<< pdiffc >>
rect 35 451 69 485
rect 119 383 153 417
rect 119 315 153 349
rect 203 451 237 485
rect 287 383 321 417
rect 287 315 321 349
rect 433 443 467 477
rect 517 451 551 485
rect 585 451 619 485
rect 669 443 703 477
rect 753 451 787 485
rect 753 383 787 417
rect 837 435 871 469
rect 940 451 974 485
rect 940 383 974 417
rect 1024 443 1058 477
rect 1024 375 1058 409
rect 1115 383 1217 485
rect 1277 443 1311 477
rect 1277 375 1311 409
rect 1361 451 1395 485
rect 1361 383 1395 417
rect 1445 443 1479 477
rect 1445 375 1479 409
rect 1529 451 1563 485
rect 1613 443 1647 477
rect 1613 375 1647 409
rect 1697 451 1731 485
rect 1697 383 1731 417
rect 1781 443 1815 477
rect 1781 375 1815 409
rect 1865 451 1899 485
rect 1865 383 1899 417
rect 1955 443 1989 477
rect 1955 375 1989 409
<< poly >>
rect 79 497 109 523
rect 163 497 193 523
rect 247 497 277 523
rect 331 497 361 523
rect 477 497 507 523
rect 629 497 659 523
rect 713 497 743 523
rect 797 497 827 523
rect 900 497 930 523
rect 984 497 1014 523
rect 1068 497 1098 523
rect 1233 497 1263 523
rect 1321 497 1351 523
rect 1405 497 1435 523
rect 1489 497 1519 523
rect 1573 497 1603 523
rect 1657 497 1687 523
rect 1741 497 1771 523
rect 1825 497 1855 523
rect 1909 497 1939 523
rect 79 265 109 297
rect 163 265 193 297
rect 247 265 277 297
rect 331 265 361 297
rect 79 261 361 265
rect 21 249 361 261
rect 21 215 37 249
rect 71 215 105 249
rect 139 215 173 249
rect 207 215 241 249
rect 275 215 361 249
rect 21 203 361 215
rect 79 199 361 203
rect 477 265 507 297
rect 629 265 659 297
rect 713 265 743 297
rect 797 265 827 297
rect 900 269 930 297
rect 984 269 1014 297
rect 1068 269 1098 297
rect 1233 269 1263 297
rect 477 249 827 265
rect 477 215 511 249
rect 545 215 579 249
rect 613 215 647 249
rect 681 215 715 249
rect 749 215 783 249
rect 817 215 827 249
rect 477 199 827 215
rect 79 177 109 199
rect 163 177 193 199
rect 247 177 277 199
rect 331 177 361 199
rect 545 177 575 199
rect 629 177 659 199
rect 713 177 743 199
rect 797 177 827 199
rect 881 249 1263 269
rect 881 215 941 249
rect 975 215 1009 249
rect 1043 215 1077 249
rect 1111 215 1145 249
rect 1179 215 1213 249
rect 1247 215 1263 249
rect 881 202 1263 215
rect 1321 269 1351 297
rect 1405 269 1435 297
rect 1489 269 1519 297
rect 1573 269 1603 297
rect 1321 249 1603 269
rect 1321 215 1337 249
rect 1371 215 1405 249
rect 1439 215 1473 249
rect 1507 215 1541 249
rect 1575 215 1603 249
rect 1321 202 1603 215
rect 881 199 1079 202
rect 881 177 911 199
rect 965 177 995 199
rect 1049 177 1079 199
rect 1133 177 1163 202
rect 1321 199 1519 202
rect 1321 177 1351 199
rect 1405 177 1435 199
rect 1489 177 1519 199
rect 1573 177 1603 202
rect 1657 265 1687 297
rect 1741 265 1771 297
rect 1825 265 1855 297
rect 1909 265 1939 297
rect 1657 261 1939 265
rect 1657 249 1995 261
rect 1657 215 1673 249
rect 1707 215 1741 249
rect 1775 215 1809 249
rect 1843 215 1877 249
rect 1911 215 1945 249
rect 1979 215 1995 249
rect 1657 203 1995 215
rect 1657 199 1939 203
rect 1657 177 1687 199
rect 1741 177 1771 199
rect 1825 177 1855 199
rect 1909 177 1939 199
rect 79 21 109 47
rect 163 21 193 47
rect 247 21 277 47
rect 331 21 361 47
rect 545 21 575 47
rect 629 21 659 47
rect 713 21 743 47
rect 797 21 827 47
rect 881 21 911 47
rect 965 21 995 47
rect 1049 21 1079 47
rect 1133 21 1163 47
rect 1321 21 1351 47
rect 1405 21 1435 47
rect 1489 21 1519 47
rect 1573 21 1603 47
rect 1657 21 1687 47
rect 1741 21 1771 47
rect 1825 21 1855 47
rect 1909 21 1939 47
<< polycont >>
rect 37 215 71 249
rect 105 215 139 249
rect 173 215 207 249
rect 241 215 275 249
rect 511 215 545 249
rect 579 215 613 249
rect 647 215 681 249
rect 715 215 749 249
rect 783 215 817 249
rect 941 215 975 249
rect 1009 215 1043 249
rect 1077 215 1111 249
rect 1145 215 1179 249
rect 1213 215 1247 249
rect 1337 215 1371 249
rect 1405 215 1439 249
rect 1473 215 1507 249
rect 1541 215 1575 249
rect 1673 215 1707 249
rect 1741 215 1775 249
rect 1809 215 1843 249
rect 1877 215 1911 249
rect 1945 215 1979 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2024 561
rect 433 485 467 493
rect 18 451 35 485
rect 69 451 203 485
rect 237 477 467 485
rect 237 451 433 477
rect 501 485 635 527
rect 501 451 517 485
rect 551 451 585 485
rect 619 451 635 485
rect 669 477 703 493
rect 21 261 65 393
rect 103 383 119 417
rect 153 383 169 417
rect 103 349 169 383
rect 270 383 287 417
rect 321 383 337 417
rect 270 349 337 383
rect 433 415 467 443
rect 669 415 703 443
rect 433 381 703 415
rect 737 485 803 527
rect 924 485 990 527
rect 737 451 753 485
rect 787 451 803 485
rect 737 417 803 451
rect 737 383 753 417
rect 787 383 803 417
rect 837 469 871 485
rect 103 315 119 349
rect 153 315 287 349
rect 321 337 337 349
rect 669 349 703 381
rect 837 349 871 435
rect 924 451 940 485
rect 974 451 990 485
rect 924 417 990 451
rect 924 383 940 417
rect 974 383 990 417
rect 1024 477 1058 493
rect 1024 409 1058 443
rect 1099 485 1233 527
rect 1099 383 1115 485
rect 1217 383 1233 485
rect 1277 477 1311 493
rect 1277 409 1311 443
rect 1024 349 1058 375
rect 1345 485 1411 527
rect 1345 451 1361 485
rect 1395 451 1411 485
rect 1345 417 1411 451
rect 1345 383 1361 417
rect 1395 383 1411 417
rect 1445 477 1479 493
rect 1445 409 1479 443
rect 1277 349 1311 375
rect 1513 485 1579 527
rect 1513 451 1529 485
rect 1563 451 1579 485
rect 1513 383 1579 451
rect 1613 477 1647 493
rect 1613 409 1647 443
rect 1445 349 1479 375
rect 1681 485 1747 527
rect 1681 451 1697 485
rect 1731 451 1747 485
rect 1681 417 1747 451
rect 1681 383 1697 417
rect 1731 383 1747 417
rect 1781 477 1815 493
rect 1781 409 1815 443
rect 1613 349 1647 375
rect 1849 485 1915 527
rect 1849 451 1865 485
rect 1899 451 1915 485
rect 1849 417 1915 451
rect 1849 383 1865 417
rect 1899 383 1915 417
rect 1955 477 1989 493
rect 1955 409 1989 443
rect 1781 349 1815 375
rect 1955 349 1989 375
rect 321 315 431 337
rect 669 315 1989 349
rect 270 299 431 315
rect 21 249 349 261
rect 21 215 37 249
rect 71 215 105 249
rect 139 215 173 249
rect 207 215 241 249
rect 275 215 349 249
rect 387 161 431 299
rect 477 249 841 265
rect 477 215 511 249
rect 545 215 579 249
rect 613 215 647 249
rect 681 215 715 249
rect 749 215 783 249
rect 817 215 841 249
rect 881 249 1263 257
rect 881 215 941 249
rect 975 215 1009 249
rect 1043 215 1077 249
rect 1111 215 1145 249
rect 1179 215 1213 249
rect 1247 215 1263 249
rect 1312 249 1591 260
rect 1312 215 1337 249
rect 1371 215 1405 249
rect 1439 215 1473 249
rect 1507 215 1541 249
rect 1575 215 1591 249
rect 1657 249 1995 256
rect 1657 215 1673 249
rect 1707 215 1741 249
rect 1775 215 1809 249
rect 1843 215 1877 249
rect 1911 215 1945 249
rect 1979 215 1995 249
rect 477 199 841 215
rect 119 127 585 161
rect 619 127 753 161
rect 787 127 803 161
rect 905 127 921 161
rect 955 127 1089 161
rect 1123 127 1361 161
rect 1395 127 1529 161
rect 1563 127 1579 161
rect 1613 127 1983 161
rect 119 101 153 127
rect 18 59 35 93
rect 69 59 85 93
rect 18 17 85 59
rect 287 109 321 127
rect 119 51 153 67
rect 187 59 203 93
rect 237 59 253 93
rect 187 17 253 59
rect 1613 101 1647 127
rect 287 51 321 75
rect 355 59 371 93
rect 405 59 421 93
rect 485 59 501 93
rect 535 59 669 93
rect 703 59 837 93
rect 871 59 1005 93
rect 1039 59 1173 93
rect 1207 59 1223 93
rect 1261 59 1277 93
rect 1311 59 1445 93
rect 1479 67 1613 93
rect 1781 101 1815 127
rect 1479 59 1647 67
rect 355 17 421 59
rect 1613 51 1647 59
rect 1681 59 1697 93
rect 1731 59 1747 93
rect 1681 17 1747 59
rect 1949 101 1983 127
rect 1781 51 1815 67
rect 1849 59 1865 93
rect 1899 59 1915 93
rect 1849 17 1915 59
rect 1949 51 1983 67
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2024 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
<< metal1 >>
rect 0 561 2024 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2024 561
rect 0 496 2024 527
rect 0 17 2024 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2024 17
rect 0 -48 2024 -17
<< labels >>
flabel locali s 305 221 339 255 0 FreeSans 200 0 0 0 B1
port 5 nsew signal input
flabel locali s 1128 221 1162 255 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 576 221 610 255 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel locali s 668 221 702 255 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel locali s 1868 221 1902 255 0 FreeSans 200 0 0 0 A4
port 4 nsew signal input
flabel locali s 1776 221 1810 255 0 FreeSans 200 0 0 0 A4
port 4 nsew signal input
flabel locali s 1684 221 1718 255 0 FreeSans 200 0 0 0 A4
port 4 nsew signal input
flabel locali s 1408 221 1442 255 0 FreeSans 200 0 0 0 A3
port 3 nsew signal input
flabel locali s 1316 221 1350 255 0 FreeSans 200 0 0 0 A3
port 3 nsew signal input
flabel locali s 1960 221 1994 255 0 FreeSans 200 0 0 0 A4
port 4 nsew signal input
flabel locali s 1036 221 1070 255 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 944 221 978 255 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 1500 221 1534 255 0 FreeSans 200 0 0 0 A3
port 3 nsew signal input
flabel locali s 760 221 794 255 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel locali s 1220 221 1254 255 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 397 221 431 255 0 FreeSans 200 0 0 0 Y
port 10 nsew signal output
flabel locali s 397 289 431 323 0 FreeSans 200 0 0 0 Y
port 10 nsew signal output
flabel locali s 484 221 518 255 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel locali s 213 221 247 255 0 FreeSans 200 0 0 0 B1
port 5 nsew signal input
flabel locali s 29 221 63 255 0 FreeSans 200 0 0 0 B1
port 5 nsew signal input
flabel locali s 29 289 63 323 0 FreeSans 200 0 0 0 B1
port 5 nsew signal input
flabel locali s 29 357 63 391 0 FreeSans 200 0 0 0 B1
port 5 nsew signal input
flabel locali s 121 221 155 255 0 FreeSans 200 0 0 0 B1
port 5 nsew signal input
flabel locali s 397 153 431 187 0 FreeSans 200 0 0 0 Y
port 10 nsew signal output
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel pwell s 46 0 46 0 0 FreeSans 200 0 0 0 VNB
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
flabel nwell s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 6 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 9 nsew power bidirectional abutment
flabel metal1 s 46 544 46 544 0 FreeSans 200 0 0 0 VPWR
flabel metal1 s 46 0 46 0 0 FreeSans 200 0 0 0 VGND
rlabel comment s 0 0 0 0 4 a41oi_4
rlabel metal1 s 0 -48 2024 48 1 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 496 2024 592 1 VPWR
port 9 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 2024 544
string GDS_END 3658588
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3642030
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
