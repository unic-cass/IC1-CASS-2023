VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO egd_top_wrapper
  CLASS BLOCK ;
  FOREIGN egd_top_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 265.795 BY 276.515 ;
  PIN la_data_in_58_43[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.070 0.000 121.350 4.000 ;
    END
  END la_data_in_58_43[0]
  PIN la_data_in_58_43[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.270 0.000 199.550 4.000 ;
    END
  END la_data_in_58_43[10]
  PIN la_data_in_58_43[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.090 0.000 207.370 4.000 ;
    END
  END la_data_in_58_43[11]
  PIN la_data_in_58_43[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.910 0.000 215.190 4.000 ;
    END
  END la_data_in_58_43[12]
  PIN la_data_in_58_43[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.730 0.000 223.010 4.000 ;
    END
  END la_data_in_58_43[13]
  PIN la_data_in_58_43[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.550 0.000 230.830 4.000 ;
    END
  END la_data_in_58_43[14]
  PIN la_data_in_58_43[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.370 0.000 238.650 4.000 ;
    END
  END la_data_in_58_43[15]
  PIN la_data_in_58_43[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 0.000 129.170 4.000 ;
    END
  END la_data_in_58_43[1]
  PIN la_data_in_58_43[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.710 0.000 136.990 4.000 ;
    END
  END la_data_in_58_43[2]
  PIN la_data_in_58_43[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.530 0.000 144.810 4.000 ;
    END
  END la_data_in_58_43[3]
  PIN la_data_in_58_43[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.350 0.000 152.630 4.000 ;
    END
  END la_data_in_58_43[4]
  PIN la_data_in_58_43[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.170 0.000 160.450 4.000 ;
    END
  END la_data_in_58_43[5]
  PIN la_data_in_58_43[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.990 0.000 168.270 4.000 ;
    END
  END la_data_in_58_43[6]
  PIN la_data_in_58_43[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.810 0.000 176.090 4.000 ;
    END
  END la_data_in_58_43[7]
  PIN la_data_in_58_43[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 0.000 183.910 4.000 ;
    END
  END la_data_in_58_43[8]
  PIN la_data_in_58_43[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.450 0.000 191.730 4.000 ;
    END
  END la_data_in_58_43[9]
  PIN la_data_in_60_59[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.190 0.000 246.470 4.000 ;
    END
  END la_data_in_60_59[0]
  PIN la_data_in_60_59[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.010 0.000 254.290 4.000 ;
    END
  END la_data_in_60_59[1]
  PIN la_data_in_65
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.830 0.000 262.110 4.000 ;
    END
  END la_data_in_65
  PIN la_data_out_23_16[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.770 0.000 4.050 4.000 ;
    END
  END la_data_out_23_16[0]
  PIN la_data_out_23_16[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 0.000 11.870 4.000 ;
    END
  END la_data_out_23_16[1]
  PIN la_data_out_23_16[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END la_data_out_23_16[2]
  PIN la_data_out_23_16[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.230 0.000 27.510 4.000 ;
    END
  END la_data_out_23_16[3]
  PIN la_data_out_23_16[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.050 0.000 35.330 4.000 ;
    END
  END la_data_out_23_16[4]
  PIN la_data_out_23_16[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.870 0.000 43.150 4.000 ;
    END
  END la_data_out_23_16[5]
  PIN la_data_out_23_16[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.690 0.000 50.970 4.000 ;
    END
  END la_data_out_23_16[6]
  PIN la_data_out_23_16[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.510 0.000 58.790 4.000 ;
    END
  END la_data_out_23_16[7]
  PIN la_data_out_26_24[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.330 0.000 66.610 4.000 ;
    END
  END la_data_out_26_24[0]
  PIN la_data_out_26_24[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 4.000 ;
    END
  END la_data_out_26_24[1]
  PIN la_data_out_26_24[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.970 0.000 82.250 4.000 ;
    END
  END la_data_out_26_24[2]
  PIN la_data_out_30_27[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.790 0.000 90.070 4.000 ;
    END
  END la_data_out_30_27[0]
  PIN la_data_out_30_27[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.610 0.000 97.890 4.000 ;
    END
  END la_data_out_30_27[1]
  PIN la_data_out_30_27[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.430 0.000 105.710 4.000 ;
    END
  END la_data_out_30_27[2]
  PIN la_data_out_30_27[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.250 0.000 113.530 4.000 ;
    END
  END la_data_out_30_27[3]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 264.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 264.080 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 264.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 264.080 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 137.400 4.000 138.000 ;
    END
  END wb_clk_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 259.900 263.925 ;
      LAYER met1 ;
        RECT 2.830 0.380 265.350 264.080 ;
      LAYER met2 ;
        RECT 2.860 4.280 265.720 264.025 ;
        RECT 2.860 0.350 3.490 4.280 ;
        RECT 4.330 0.350 11.310 4.280 ;
        RECT 12.150 0.350 19.130 4.280 ;
        RECT 19.970 0.350 26.950 4.280 ;
        RECT 27.790 0.350 34.770 4.280 ;
        RECT 35.610 0.350 42.590 4.280 ;
        RECT 43.430 0.350 50.410 4.280 ;
        RECT 51.250 0.350 58.230 4.280 ;
        RECT 59.070 0.350 66.050 4.280 ;
        RECT 66.890 0.350 73.870 4.280 ;
        RECT 74.710 0.350 81.690 4.280 ;
        RECT 82.530 0.350 89.510 4.280 ;
        RECT 90.350 0.350 97.330 4.280 ;
        RECT 98.170 0.350 105.150 4.280 ;
        RECT 105.990 0.350 112.970 4.280 ;
        RECT 113.810 0.350 120.790 4.280 ;
        RECT 121.630 0.350 128.610 4.280 ;
        RECT 129.450 0.350 136.430 4.280 ;
        RECT 137.270 0.350 144.250 4.280 ;
        RECT 145.090 0.350 152.070 4.280 ;
        RECT 152.910 0.350 159.890 4.280 ;
        RECT 160.730 0.350 167.710 4.280 ;
        RECT 168.550 0.350 175.530 4.280 ;
        RECT 176.370 0.350 183.350 4.280 ;
        RECT 184.190 0.350 191.170 4.280 ;
        RECT 192.010 0.350 198.990 4.280 ;
        RECT 199.830 0.350 206.810 4.280 ;
        RECT 207.650 0.350 214.630 4.280 ;
        RECT 215.470 0.350 222.450 4.280 ;
        RECT 223.290 0.350 230.270 4.280 ;
        RECT 231.110 0.350 238.090 4.280 ;
        RECT 238.930 0.350 245.910 4.280 ;
        RECT 246.750 0.350 253.730 4.280 ;
        RECT 254.570 0.350 261.550 4.280 ;
        RECT 262.390 0.350 265.720 4.280 ;
      LAYER met3 ;
        RECT 3.745 138.400 265.355 264.005 ;
        RECT 4.400 137.000 265.355 138.400 ;
        RECT 3.745 4.255 265.355 137.000 ;
      LAYER met4 ;
        RECT 4.895 10.240 20.640 237.825 ;
        RECT 23.040 10.240 97.440 237.825 ;
        RECT 99.840 10.240 174.240 237.825 ;
        RECT 176.640 10.240 251.040 237.825 ;
        RECT 253.440 10.240 261.905 237.825 ;
        RECT 4.895 4.255 261.905 10.240 ;
  END
END egd_top_wrapper
END LIBRARY

