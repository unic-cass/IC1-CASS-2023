magic
tech sky130B
magscale 1 2
timestamp 1676037725
<< metal1 >>
tri 4773 8766 4810 8803 sw
tri 846 8565 1026 8745 nw
tri 4697 8711 4731 8745 ne
tri 4833 8630 4867 8664 nw
rect 1602 8543 4514 8595
tri 1210 8514 1239 8543 nw
tri 4437 8512 4468 8543 ne
tri 6246 8505 6405 8664 ne
tri 6655 8505 6814 8664 nw
tri 8156 8630 8190 8664 ne
tri 8607 8622 8641 8656 nw
tri 13133 8622 13167 8656 ne
tri 4321 8269 4324 8272 se
tri 4370 8269 4373 8272 sw
tri 584 8198 618 8232 ne
tri 497 8129 522 8154 ne
tri 4321 8138 4324 8141 ne
tri 4370 8138 4373 8141 nw
tri 408 8055 433 8080 ne
tri 159 7426 193 7460 ne
tri 1210 7389 1284 7463 sw
rect 1201 7275 4220 7389
tri 4220 7275 4334 7389 sw
tri 13579 7356 13582 7359 ne
tri 4434 7275 4468 7309 se
rect 1266 7223 4514 7275
tri 846 7090 920 7164 sw
tri 4697 7090 4731 7124 se
rect 4266 7039 4737 7044
tri 687 6937 788 7038 se
rect 788 6937 976 7038
tri 83 6873 147 6937 se
rect 147 6891 976 6937
tri 976 6891 1123 7038 nw
rect 2187 6940 3802 6992
tri 3780 6918 3802 6940 ne
tri 3802 6930 3864 6992 sw
rect 3802 6918 3864 6930
tri 3802 6908 3812 6918 ne
rect 147 6873 149 6891
tri 149 6873 167 6891 nw
tri 49 6797 83 6831 se
rect 83 6797 129 6873
tri 129 6853 149 6873 nw
tri 245 6806 279 6840 sw
rect -74 6669 129 6797
tri 245 6720 279 6754 nw
tri 129 6669 177 6717 sw
tri -809 6593 -803 6599 nw
tri 83 6575 177 6669 ne
tri 177 6663 183 6669 sw
tri 240 6663 296 6719 se
rect 296 6716 304 6719
tri 870 6716 873 6719 sw
rect 296 6663 2180 6716
rect 177 6630 2180 6663
tri 3401 6652 3475 6726 se
rect 3475 6674 3633 6726
tri 3475 6652 3497 6674 nw
rect 177 6575 890 6630
tri 177 6547 205 6575 ne
rect 205 6547 890 6575
tri 890 6547 973 6630 nw
tri 3365 6616 3401 6652 se
rect 3401 6616 3417 6652
rect 1181 6360 1336 6385
tri 1336 6360 1361 6385 sw
rect 1181 6255 2292 6360
tri 1282 6230 1307 6255 ne
rect 1307 6230 2292 6255
tri 756 6178 790 6212 sw
tri 944 6178 956 6190 se
rect 756 6150 956 6178
tri 944 6138 956 6150 ne
tri 2771 5841 2805 5875 ne
rect 2122 5704 2160 5756
tri 2160 5704 2212 5756 sw
tri 1585 5599 1619 5633 ne
tri 2138 5630 2212 5704 ne
tri 2212 5630 2286 5704 sw
tri 2515 5635 2549 5669 ne
tri 1492 5537 1526 5571 ne
tri 2212 5556 2286 5630 ne
tri 2286 5556 2360 5630 sw
tri 2286 5482 2360 5556 ne
tri 2360 5482 2434 5556 sw
tri 2360 5408 2434 5482 ne
tri 2434 5414 2502 5482 sw
rect 2434 5408 2502 5414
tri -449 5357 -415 5391 se
tri 71 5377 97 5403 nw
tri 2434 5392 2450 5408 ne
tri -369 5357 -351 5375 sw
tri -457 5277 -423 5311 ne
tri -383 5279 -351 5311 nw
tri 844 5203 849 5208 nw
tri 2376 5157 2450 5231 se
rect 2450 5209 2502 5408
tri 2450 5157 2502 5209 nw
tri 2510 5157 2549 5196 se
rect 2549 5174 2601 5707
rect 3365 5549 3417 6616
tri 3417 6594 3475 6652 nw
tri 3678 6332 3712 6366 se
rect 3448 6280 3712 6332
rect 3448 5743 3500 6280
tri 3500 6230 3550 6280 nw
tri 3681 6249 3712 6280 ne
rect 3812 5708 3864 6918
tri 4266 6629 4676 7039 ne
rect 4676 6629 4737 7039
tri 7907 6797 7941 6831 se
tri 8800 6769 8834 6803 sw
tri 11321 6769 11404 6852 se
rect 4046 6568 4549 6629
tri 4549 6568 4610 6629 sw
tri 4676 6568 4737 6629 ne
rect 4046 6475 4610 6568
tri 4610 6475 4703 6568 sw
tri 4833 6542 4867 6576 sw
tri 8156 6542 8190 6576 se
tri 8607 6542 8641 6576 sw
tri 11563 6542 11597 6576 se
tri 11699 6542 11733 6576 sw
rect 4046 6455 4703 6475
tri 4493 6377 4571 6455 ne
rect 3895 5984 3947 6197
tri 3947 6163 3981 6197 nw
tri 3947 5984 3969 6006 sw
rect 4046 6005 4351 6179
tri 3895 5910 3969 5984 ne
tri 3969 5961 3992 5984 sw
rect 3969 5910 4036 5961
tri 4295 5949 4351 6005 ne
tri 4351 5989 4541 6179 sw
rect 4351 5949 4541 5989
tri 3969 5843 4036 5910 ne
tri 4351 5891 4409 5949 ne
tri 3812 5656 3864 5708 ne
tri 3864 5705 3889 5730 sw
rect 3864 5656 3889 5705
tri 3864 5631 3889 5656 ne
tri 3889 5631 3963 5705 sw
tri 3417 5549 3451 5583 sw
tri 3889 5557 3963 5631 ne
tri 3963 5557 4037 5631 sw
tri 2930 5534 2938 5542 se
tri 2971 5534 2976 5539 sw
rect 3365 5497 3535 5549
tri 3963 5483 4037 5557 ne
tri 4037 5483 4111 5557 sw
rect 4409 5507 4541 5949
rect 4571 5894 4703 6455
tri 4833 6406 4867 6440 nw
tri 8156 6406 8190 6440 ne
tri 8607 6406 8641 6440 nw
tri 11563 6406 11597 6440 ne
tri 11699 6406 11733 6440 nw
tri 7907 6151 7941 6185 ne
tri 11370 6179 11404 6213 ne
tri 2976 5438 3010 5472 sw
tri 3289 5442 3323 5476 sw
tri 3687 5442 3721 5476 se
tri 3289 5413 3291 5415 nw
tri 4037 5409 4111 5483 ne
tri 4111 5409 4185 5483 sw
tri 4612 5409 4742 5539 se
tri 2758 5381 2760 5383 ne
tri 2812 5349 2846 5383 nw
tri 3197 5351 3231 5385 sw
rect 3613 5309 3696 5351
tri 3696 5309 3738 5351 sw
tri 4111 5335 4185 5409 ne
tri 4185 5335 4259 5409 sw
tri 3189 5271 3223 5305 nw
rect 3613 5299 3738 5309
tri 3647 5260 3686 5299 ne
rect 2549 5157 2564 5174
tri 2333 5114 2376 5157 se
rect 2376 5114 2407 5157
tri 2407 5114 2450 5157 nw
tri 2490 5137 2510 5157 se
rect 2510 5137 2564 5157
tri 2564 5137 2601 5174 nw
tri 2467 5114 2490 5137 se
tri -9 5040 25 5074 se
tri 71 5040 105 5074 sw
rect 2282 5062 2355 5114
tri 2355 5062 2407 5114 nw
tri 2416 5063 2467 5114 se
rect 2467 5063 2490 5114
tri 2490 5063 2564 5137 nw
tri 2913 5127 2917 5131 ne
tri 2415 5062 2416 5063 se
tri 2342 4989 2415 5062 se
rect 2415 4989 2416 5062
tri 2416 4989 2490 5063 nw
tri 2623 5020 2657 5054 se
tri 2703 5020 2737 5054 sw
tri 3189 5020 3223 5054 sw
tri 2268 4915 2342 4989 se
tri 2342 4915 2416 4989 nw
tri 2246 4893 2268 4915 se
rect 2081 4841 2268 4893
tri 2268 4841 2342 4915 nw
tri 3426 4813 3451 4838 se
tri 3427 4705 3451 4729 ne
tri 3652 4376 3686 4410 se
rect 3686 4376 3738 5299
tri 3824 5212 3906 5294 nw
tri 4185 5261 4259 5335 ne
tri 4259 5261 4333 5335 sw
tri 4259 5239 4281 5261 ne
tri 3932 5123 3936 5127 ne
rect 3971 5122 3975 5127
tri 3971 5118 3975 5122 ne
tri 3975 5118 3984 5127 nw
tri 3852 5024 3856 5028 ne
tri 3895 5019 3904 5028 nw
tri 4127 4702 4152 4727 nw
tri 4011 4616 4024 4629 ne
tri 4050 4616 4063 4629 nw
rect 4281 4617 4333 5261
tri 4456 5253 4612 5409 se
rect 4612 5253 4742 5409
rect 4456 4685 4742 5253
tri 4456 4410 4731 4685 ne
rect 4731 4410 4742 4685
tri 5115 4647 5118 4650 ne
tri 8751 4647 8754 4650 ne
tri 8800 4647 8803 4650 nw
tri 5032 4581 5066 4615 sw
tri 7907 4581 7941 4615 se
tri 8800 4553 8834 4587 sw
rect 3441 4324 3738 4376
tri -651 3936 -617 3970 nw
tri 2768 3936 2802 3970 ne
tri -215 3811 -181 3845 ne
tri 266 3826 272 3832 ne
tri 620 3794 643 3817 se
tri 695 3794 729 3828 sw
tri 2332 3811 2366 3845 nw
tri -767 3595 -722 3640 se
rect -662 3561 -659 3627
tri -659 3561 -593 3627 sw
tri -508 3562 -488 3582 se
tri -442 3562 -422 3582 sw
rect -615 3240 -614 3264
rect -658 3236 -614 3240
tri -614 3236 -586 3264 nw
tri -511 3236 -488 3259 ne
rect -488 3236 -483 3259
rect -443 3236 -442 3258
tri -442 3236 -420 3258 nw
tri -767 3177 -721 3223 ne
rect -721 3187 -711 3223
tri -658 3192 -614 3236 nw
tri 1260 3231 1410 3381 nw
tri 1749 3347 1783 3381 ne
tri 1829 3347 1863 3381 nw
tri 2455 3347 2489 3381 ne
tri 2535 3347 2569 3381 nw
tri 2740 3353 2768 3381 ne
tri 2814 3347 2848 3381 nw
tri 1485 3338 1487 3340 se
rect 1487 3338 1493 3340
tri 1857 3324 1870 3337 se
rect 1870 3324 2243 3337
rect 1857 3305 2243 3324
rect 1857 3299 1907 3305
tri 1518 3260 1552 3294 nw
tri 1907 3274 1938 3305 nw
tri 2151 3265 2191 3305 ne
rect 2191 3299 2243 3305
tri -721 3177 -711 3187 nw
tri 1023 3142 1104 3223 ne
tri 1672 3194 1679 3201 sw
tri 3407 3196 3441 3230 se
rect 3441 3170 3493 4324
tri 3493 4290 3527 4324 nw
tri 4833 4318 4867 4352 sw
tri 8156 4318 8190 4352 se
tri 8607 4326 8641 4360 sw
tri 13739 4341 13741 4343 ne
tri 14871 4326 14905 4360 se
tri 15012 4326 15023 4337 sw
tri 13165 4292 13199 4326 ne
tri 13245 4292 13279 4326 nw
tri 14943 4292 14977 4326 ne
tri 3744 4243 3778 4277 se
tri 6665 4242 6668 4245 ne
tri 6714 4242 6717 4245 nw
tri 6991 4242 6994 4245 ne
tri 7040 4242 7043 4245 nw
tri 7317 4242 7320 4245 ne
tri 7366 4242 7369 4245 nw
tri 11024 4242 11027 4245 ne
tri 11073 4242 11076 4245 nw
tri 3583 4163 3617 4197 nw
tri 4209 4188 4243 4222 sw
tri 11904 4196 11977 4269 se
rect 11977 4217 12942 4269
rect 13674 4223 14669 4269
tri 13674 4217 13680 4223 nw
rect 11977 4196 11978 4217
tri 11978 4196 11999 4217 nw
tri 14649 4203 14669 4223 ne
tri 14669 4205 14733 4269 sw
rect 14669 4203 14733 4205
rect 10440 4144 11926 4196
tri 11926 4144 11978 4196 nw
tri 14669 4185 14687 4203 ne
tri 13480 4106 13514 4140 nw
tri 14667 4109 14687 4129 se
rect 14687 4109 14733 4203
tri 14655 4097 14667 4109 se
rect 14667 4097 14675 4109
tri 4209 4051 4243 4085 sw
rect 14538 4051 14675 4097
tri 14675 4051 14733 4109 nw
tri 4209 3994 4238 4023 nw
tri 10125 3970 10159 4004 ne
tri 10709 3967 10743 4001 ne
tri 10797 3999 10827 4029 sw
tri 13686 4017 13720 4051 ne
tri 13772 4017 13806 4051 nw
tri 13428 4004 13431 4007 ne
tri 13477 4004 13480 4007 nw
tri 13881 3980 13924 4023 se
rect 13924 3980 14606 4023
tri 14606 3980 14649 4023 sw
tri 4430 3914 4464 3948 sw
tri 13829 3928 13881 3980 se
rect 13881 3928 13920 3980
tri 13920 3945 13955 3980 nw
tri 5614 3892 5619 3897 ne
rect 5619 3892 5623 3897
tri 10743 3871 10777 3905 ne
tri 7543 3812 7577 3846 ne
tri 4228 3722 4262 3756 nw
tri 7993 3711 8017 3735 se
tri 4447 3649 4481 3683 nw
tri 8327 3653 8456 3782 se
rect 8456 3655 9400 3782
rect 8456 3653 8464 3655
rect 11452 3604 11880 3862
rect 11952 3755 12380 3862
tri 11952 3700 12007 3755 ne
rect 12007 3709 12380 3755
tri 12380 3709 12485 3814 sw
tri 13549 3797 13552 3800 ne
tri 13598 3797 13601 3800 nw
tri 13669 3725 13711 3767 se
rect 13711 3747 13757 3829
rect 14195 3810 14574 3952
tri 14589 3951 14618 3980 ne
rect 14618 3967 14649 3980
tri 14649 3967 14662 3980 sw
rect 13711 3725 13735 3747
tri 13735 3725 13757 3747 nw
rect 12007 3700 13014 3709
tri 11880 3604 11976 3700 sw
tri 12007 3657 12050 3700 ne
rect 12050 3657 13014 3700
tri 13603 3659 13669 3725 se
tri 13669 3659 13735 3725 nw
tri 13954 3661 13980 3687 se
rect 13980 3667 14026 3758
tri 14026 3749 14035 3758 nw
rect 14195 3733 14418 3779
tri 14452 3734 14528 3810 ne
rect 13980 3661 14000 3667
tri 13557 3613 13603 3659 se
rect 11452 3552 13052 3604
tri 4228 3412 4262 3446 sw
tri 5416 3417 5450 3451 se
tri 5710 3433 5744 3467 sw
rect 5708 3399 5710 3408
tri 5710 3399 5719 3408 nw
tri 4228 3331 4262 3365 nw
tri 6494 3354 6511 3371 se
tri 6563 3354 6586 3377 sw
tri 6494 3290 6512 3308 ne
tri 6563 3274 6597 3308 nw
tri 6745 3277 6779 3311 se
tri 6825 3277 6859 3311 sw
tri 3407 3110 3441 3144 ne
rect 12450 3131 12468 3292
tri 6592 3107 6616 3131 nw
tri -215 2973 -181 3007 se
tri 620 3000 644 3024 ne
tri 695 2990 729 3024 nw
tri 270 2986 273 2989 se
tri 1260 2961 1374 3075 sw
tri 2691 3068 2725 3102 sw
tri 12025 3062 12094 3131 ne
tri 12399 3062 12468 3131 ne
rect 12468 3062 12486 3131
tri 2691 3034 2697 3040 nw
tri 270 2937 273 2940 ne
tri -651 2848 -617 2882 sw
tri 8956 2829 9018 2891 ne
rect 3186 2675 3238 2766
tri 3238 2721 3272 2755 sw
tri 3345 2721 3379 2755 se
tri 2741 2643 2773 2675 se
tri 4229 2655 4263 2689 nw
tri 13053 2492 13113 2552 se
rect 13113 2492 13165 3392
rect 13557 3376 13603 3613
tri 13603 3593 13669 3659 nw
tri 13742 3550 13824 3632 ne
tri 13921 3374 13954 3407 se
rect 13954 3374 14000 3661
tri 14000 3641 14026 3667 nw
tri 14047 3628 14063 3644 se
rect 14063 3628 14115 3707
tri 14195 3699 14229 3733 nw
tri 14338 3699 14372 3733 ne
rect 14372 3690 14418 3733
rect 14047 3622 14115 3628
tri 14000 3374 14038 3412 sw
rect 14047 3408 14099 3622
tri 14099 3606 14115 3622 nw
tri 14135 3529 14256 3650 se
rect 14135 3440 14256 3529
tri 14047 3364 14091 3408 ne
rect 14091 3374 14099 3408
tri 14099 3374 14161 3436 sw
tri 14468 3421 14528 3481 se
rect 14528 3461 14574 3810
rect 14528 3421 14534 3461
tri 14534 3421 14574 3461 nw
rect 13847 3232 14251 3302
rect 13448 3155 13797 3201
tri 13813 3198 13847 3232 ne
tri 13565 3149 13571 3155 nw
tri 13813 3124 13847 3158 se
rect 13847 3124 13953 3232
tri 13953 3198 13987 3232 nw
tri 13953 3124 13987 3158 sw
rect 13847 3054 14251 3124
rect 14468 3106 14514 3421
tri 14514 3401 14534 3421 nw
tri 14550 3345 14618 3413 se
rect 14618 3383 14662 3967
rect 14618 3345 14624 3383
tri 14624 3345 14662 3383 nw
rect 14550 3290 14596 3345
tri 14596 3317 14624 3345 nw
rect 13557 2957 13603 2979
tri 13245 2883 13279 2917 sw
tri 13557 2911 13603 2957 ne
tri 13603 2945 13635 2977 sw
tri 14440 2945 14468 2973 se
rect 14468 2953 14514 2976
rect 14468 2945 14472 2953
rect 13603 2911 14472 2945
tri 14472 2911 14514 2953 nw
tri 14943 2883 14977 2917 se
tri 13245 2803 13279 2837 nw
tri 14943 2803 14977 2837 ne
rect 12881 2378 13165 2492
tri 2748 2358 2754 2364 se
rect 2754 2358 2755 2364
rect 12881 2330 13117 2378
tri 13117 2330 13165 2378 nw
tri 13281 2732 13349 2800 se
rect 13349 2748 14030 2800
rect 13349 2732 13355 2748
tri 13355 2732 13371 2748 nw
tri 8854 2192 8880 2218 se
tri 4278 2018 4381 2121 se
rect 4381 2028 5267 2121
tri 9002 2119 9090 2207 se
rect 9090 2119 9280 2293
tri 9817 2119 9823 2125 sw
rect 4381 2018 4394 2028
tri 4394 2018 4404 2028 nw
tri 1495 1935 1502 1942 ne
rect 1502 1935 1507 1942
rect 4215 1890 4266 2018
tri 4266 1890 4394 2018 nw
tri 5155 1916 5267 2028 ne
rect 9110 1916 9280 2119
tri 2087 1402 2098 1413 se
tri 2090 1367 2098 1375 ne
rect 2098 1367 2108 1375
tri -977 1224 -943 1258 sw
rect -317 1125 217 1224
tri -311 1066 -252 1125 nw
tri 3682 860 3715 893 se
rect 3715 871 3767 1890
tri 8552 1876 8558 1882 se
rect 8558 1876 8562 1882
tri 8686 1875 8693 1882 sw
tri 5854 1836 5878 1860 nw
tri 6982 1770 7016 1804 ne
tri 7607 1802 7641 1836 sw
tri 5628 1736 5662 1770 nw
tri 5729 1736 5763 1770 ne
tri 5809 1736 5843 1770 nw
tri 6600 1742 6618 1760 se
tri 7382 1737 7395 1750 se
tri 7607 1722 7641 1756 nw
tri 5976 1680 6010 1714 nw
tri 7041 1692 7062 1713 sw
tri 6612 1670 6620 1678 se
rect 5587 1583 5588 1589
tri 5588 1583 5594 1589 sw
tri 5992 1583 6026 1617 se
rect 6026 1583 6072 1657
tri 7361 1651 7395 1685 ne
tri 8086 1648 8120 1682 nw
tri 6072 1597 6106 1631 nw
tri 6250 1597 6284 1631 ne
tri 6418 1590 6452 1624 nw
rect 5588 1537 6072 1583
tri 6566 1570 6620 1624 ne
tri 8672 1592 8706 1626 ne
tri 7149 1506 7183 1540 nw
tri 8444 1536 8478 1570 ne
tri 8290 1450 8324 1484 se
tri 8359 1451 8367 1459 se
rect 8359 1450 8367 1451
tri 8367 1450 8376 1459 sw
tri 8966 1434 8967 1435 se
tri 9013 1434 9047 1468 sw
tri 6618 1352 6652 1386 sw
tri 7524 1370 7558 1404 sw
tri 8477 1370 8511 1404 se
tri 9646 1296 9689 1339 se
rect 9689 1296 9716 1339
tri 12467 1259 12501 1293 ne
tri 6393 990 6418 1015 nw
tri 11175 980 11209 1014 ne
tri 12976 992 13021 1037 se
rect 13021 1015 13073 1246
rect 13281 1245 13333 2732
tri 13333 2710 13355 2732 nw
tri 13479 2618 13513 2652 nw
rect 13672 2519 13990 2622
tri 13990 2519 14093 2622 sw
tri 14121 2618 14155 2652 ne
rect 13672 2423 14093 2519
rect 13021 992 13050 1015
tri 13050 992 13073 1015 nw
tri 6241 935 6266 960 sw
tri 6602 937 6636 971 se
tri 6664 924 6698 958 nw
tri 11101 924 11135 958 ne
rect 11304 940 12998 992
tri 12998 940 13050 992 nw
rect 6233 908 6241 912
tri 6241 908 6245 912 nw
rect 3715 860 3734 871
tri 3628 723 3682 777 se
rect 3682 723 3734 860
tri 3734 838 3767 871 nw
tri 6659 862 6693 896 se
rect 6719 844 6721 869
tri 6721 844 6746 869 nw
tri 6924 844 6948 868 ne
rect 6948 844 6949 868
tri 3776 795 3804 823 se
tri 6744 810 6773 839 se
rect 6773 810 6785 839
rect 974 721 3734 723
rect 974 671 3684 721
tri 3684 671 3734 721 nw
tri 3896 686 3930 720 sw
tri 7688 686 7694 692 sw
tri 8595 642 8601 648 nw
rect 11304 627 11356 940
tri 11356 906 11390 940 nw
tri 6994 612 7007 625 se
tri 6996 573 7007 584 ne
tri 7142 543 7162 563 se
tri 7155 511 7162 518 ne
tri 5267 423 5301 457 ne
tri 7627 448 7661 482 nw
rect 9667 456 9670 462
tri 9670 456 9676 462 nw
tri 7670 446 7674 450 se
tri 10959 448 10993 482 ne
tri 4121 389 4145 413 se
rect 7670 402 7674 446
tri 4283 281 4307 305 ne
tri 4614 300 4648 334 sw
tri 8063 323 8097 357 ne
tri 8521 338 8527 344 ne
tri 10102 338 10108 344 nw
tri 10523 323 10557 357 nw
tri 9595 306 9598 309 se
tri 11237 293 11261 317 sw
tri 13479 314 13513 348 sw
tri 14121 314 14155 348 se
rect 14155 314 14701 2652
tri 3715 263 3729 277 se
rect 3729 263 3739 277
tri 3714 225 3729 240 ne
rect 3729 225 3748 240
tri 5917 230 5951 264 ne
tri 9595 257 9598 260 ne
tri 5997 220 6031 254 nw
tri 5490 207 5496 213 se
rect 3680 186 3687 207
tri 3687 186 3708 207 sw
tri 3927 186 3948 207 se
rect 3948 186 3955 207
tri 3635 159 3655 179 ne
rect 3655 159 3657 179
rect 3976 159 3978 179
tri 3978 159 3998 179 nw
tri 5462 143 5496 177 ne
tri 11311 107 11499 295 se
rect 13433 118 14745 314
rect 11109 104 11499 107
rect 11109 -107 11683 104
tri 11683 -107 11894 104 nw
tri 13245 30 13279 64 sw
tri 14943 30 14977 64 se
tri -797 -472 -763 -438 nw
<< metal2 >>
tri 7818 8907 7993 9082 se
rect 7993 8982 8231 9829
rect 7993 8907 8156 8982
tri 8156 8907 8231 8982 nw
rect 1185 8724 1794 8878
tri 1794 8724 1948 8878 sw
tri 1730 8506 1948 8724 ne
tri 1948 8507 2165 8724 sw
tri 3798 8569 4136 8907 se
rect 4136 8669 7918 8907
tri 7918 8669 8156 8907 nw
rect 4136 8628 4195 8669
tri 4195 8628 4236 8669 nw
tri 9037 8628 9212 8803 se
rect 9212 8703 9450 9825
rect 9212 8628 9237 8703
tri 4136 8569 4195 8628 nw
tri 3736 8507 3798 8569 se
rect 3798 8507 4045 8569
rect 1948 8506 4045 8507
tri 1948 8412 2042 8506 ne
rect 2042 8478 4045 8506
tri 4045 8478 4136 8569 nw
tri 4222 8564 4286 8628 se
rect 4286 8564 9237 8628
tri 4136 8478 4222 8564 se
rect 4222 8490 9237 8564
tri 9237 8490 9450 8703 nw
tri 11756 8513 11807 8564 se
rect 11807 8513 14064 8564
tri 14064 8513 14115 8564 sw
tri 11733 8490 11756 8513 se
rect 11756 8512 14115 8513
rect 11756 8490 11807 8512
tri 11807 8490 11829 8512 nw
rect 4222 8478 9137 8490
rect 2042 8472 4039 8478
tri 4039 8472 4045 8478 nw
tri 4130 8472 4136 8478 se
rect 4136 8472 9137 8478
rect 2042 8381 3948 8472
tri 3948 8381 4039 8472 nw
tri 4039 8381 4130 8472 se
rect 4130 8390 9137 8472
tri 9137 8390 9237 8490 nw
tri 11659 8416 11733 8490 se
tri 11733 8416 11807 8490 nw
tri 14006 8455 14063 8512 ne
rect 4130 8381 4265 8390
rect 2042 8290 3857 8381
tri 3857 8290 3948 8381 nw
tri 3948 8290 4039 8381 se
rect 4039 8290 4265 8381
rect 2042 8269 3836 8290
tri 3836 8269 3857 8290 nw
tri 3927 8269 3948 8290 se
rect 3948 8269 4265 8290
tri 4265 8269 4386 8390 nw
tri 11585 8342 11659 8416 se
tri 11659 8342 11733 8416 nw
tri 11575 8332 11585 8342 se
rect 11585 8332 11649 8342
tri 11649 8332 11659 8342 nw
rect 2042 8117 2803 8269
tri 2803 8117 2955 8269 nw
tri 3610 7952 3927 8269 se
rect 3927 8248 4244 8269
tri 4244 8248 4265 8269 nw
tri 4286 8248 4307 8269 se
rect 4307 8248 4373 8269
rect 3927 8206 4202 8248
tri 4202 8206 4244 8248 nw
tri 4244 8206 4286 8248 se
rect 4286 8206 4373 8248
rect 3927 8183 4179 8206
tri 4179 8183 4202 8206 nw
tri 4221 8183 4244 8206 se
rect 4244 8183 4373 8206
rect 3927 8141 4137 8183
tri 4137 8141 4179 8183 nw
tri 4179 8141 4221 8183 se
rect 4221 8145 4373 8183
rect 4221 8141 4370 8145
tri 4370 8142 4373 8145 nw
rect 3927 8109 4105 8141
tri 4105 8109 4137 8141 nw
tri 4147 8109 4179 8141 se
rect 3927 8067 4063 8109
tri 4063 8067 4105 8109 nw
tri 4105 8067 4147 8109 se
rect 4147 8067 4179 8109
tri 4179 8067 4253 8141 nw
tri 11453 8136 11649 8332 nw
rect 3927 8035 4031 8067
tri 4031 8035 4063 8067 nw
tri 4073 8035 4105 8067 se
rect 3927 7993 3989 8035
tri 3989 7993 4031 8035 nw
tri 4031 7993 4073 8035 se
rect 4073 7993 4105 8035
tri 4105 7993 4179 8067 nw
rect 3927 7952 3948 7993
tri 3948 7952 3989 7993 nw
tri 3990 7952 4031 7993 se
tri 3525 7867 3610 7952 se
rect 3610 7910 3906 7952
tri 3906 7910 3948 7952 nw
tri 3957 7919 3990 7952 se
rect 3990 7919 4031 7952
tri 4031 7919 4105 7993 nw
tri 3948 7910 3957 7919 se
rect 3610 7909 3905 7910
tri 3905 7909 3906 7910 nw
tri 3947 7909 3948 7910 se
rect 3948 7909 3957 7910
rect 3610 7867 3863 7909
tri 3863 7867 3905 7909 nw
tri 3905 7867 3947 7909 se
rect 3947 7867 3957 7909
rect 2042 7825 3821 7867
tri 3821 7825 3863 7867 nw
tri 3883 7845 3905 7867 se
rect 3905 7845 3957 7867
tri 3957 7845 4031 7919 nw
tri 3863 7825 3883 7845 se
rect 2042 7813 3809 7825
tri 3809 7813 3821 7825 nw
tri 3851 7813 3863 7825 se
rect 3863 7813 3883 7825
rect 2042 7771 3767 7813
tri 3767 7771 3809 7813 nw
tri 3809 7771 3851 7813 se
rect 3851 7771 3883 7813
tri 3883 7771 3957 7845 nw
tri 6913 7838 6985 7910 se
rect 2042 7739 3735 7771
tri 3735 7739 3767 7771 nw
tri 3777 7739 3809 7771 se
rect 2042 7697 3693 7739
tri 3693 7697 3735 7739 nw
tri 3735 7697 3777 7739 se
rect 3777 7697 3809 7739
tri 3809 7697 3883 7771 nw
tri 1842 7493 2042 7693 se
rect 2042 7665 3661 7697
tri 3661 7665 3693 7697 nw
tri 3703 7665 3735 7697 se
rect 2042 7623 3619 7665
tri 3619 7623 3661 7665 nw
tri 3661 7623 3703 7665 se
rect 3703 7623 3735 7665
tri 3735 7623 3809 7697 nw
tri 4760 7631 4791 7662 se
rect 4791 7631 6136 7662
rect 2042 7591 3587 7623
tri 3587 7591 3619 7623 nw
tri 3629 7591 3661 7623 se
rect 2042 7549 3545 7591
tri 3545 7549 3587 7591 nw
tri 3587 7549 3629 7591 se
rect 3629 7549 3661 7591
tri 3661 7549 3735 7623 nw
rect 2042 7535 3531 7549
tri 3531 7535 3545 7549 nw
tri 3573 7535 3587 7549 se
rect 2042 7493 3489 7535
tri 3489 7493 3531 7535 nw
tri 3531 7493 3573 7535 se
rect 3573 7493 3587 7535
tri 1754 7405 1842 7493 se
rect 1842 7405 1908 7493
tri 1690 7079 1754 7143 se
rect 1754 7079 1908 7405
tri 1908 7341 2060 7493 nw
tri 3513 7475 3531 7493 se
rect 3531 7475 3587 7493
tri 3587 7475 3661 7549 nw
tri 3479 7441 3513 7475 se
rect 3513 7441 3553 7475
tri 3553 7441 3587 7475 nw
tri 2187 7367 2261 7441 se
rect 2261 7389 3501 7441
tri 3501 7389 3553 7441 nw
tri 2261 7367 2283 7389 nw
tri 2113 7293 2187 7367 se
tri 2187 7293 2261 7367 nw
tri 4490 7361 4760 7631 se
rect 4760 7498 6136 7631
tri 6136 7498 6300 7662 sw
tri 9707 7498 9779 7570 nw
rect 4760 7470 6300 7498
tri 4760 7361 4869 7470 nw
tri 4447 7318 4490 7361 se
rect 4490 7318 4525 7361
tri 1665 7054 1690 7079 se
rect 1690 7054 1729 7079
rect 1059 6900 1729 7054
tri 1729 6900 1908 7079 nw
tri 2092 7272 2113 7293 se
rect 2113 7272 2144 7293
tri 2059 6992 2092 7025 se
rect 2092 6992 2144 7272
tri 2144 7250 2187 7293 nw
tri 2434 7048 2704 7318 se
rect 2704 7126 4525 7318
tri 4525 7126 4760 7361 nw
tri 4903 7169 5164 7430 se
rect 5164 7169 5408 7430
tri 5721 7283 5760 7322 se
tri 6058 7283 6245 7470 ne
rect 6245 7361 6300 7470
tri 6300 7361 6437 7498 sw
rect 6245 7283 9284 7361
tri 6245 7169 6359 7283 ne
rect 6359 7169 9284 7283
tri 2704 7048 2782 7126 nw
tri 4824 7090 4903 7169 se
rect 4903 7090 5408 7169
tri 2144 6992 2178 7026 sw
tri 2274 6888 2434 7048 se
rect 2434 6888 2466 7048
tri -758 6727 -688 6797 se
rect -688 6727 -74 6797
rect -803 6669 -74 6727
rect -803 6599 -704 6669
tri -704 6599 -634 6669 nw
rect 2274 6588 2466 6888
tri 2466 6810 2704 7048 nw
tri 2873 6856 3107 7090 se
rect 3107 6923 5408 7090
tri 5811 6942 5812 6943 ne
tri 3107 6856 3174 6923 nw
tri 2728 6711 2873 6856 se
rect 2873 6711 2894 6856
tri 2625 6360 2728 6463 se
rect 2728 6360 2894 6711
tri 2894 6643 3107 6856 nw
rect 3465 6834 4731 6892
rect 2484 6301 2894 6360
rect 2484 6230 2823 6301
tri 2823 6230 2894 6301 nw
tri 956 6086 1008 6138 ne
rect 1008 6043 1084 6138
tri 1008 5967 1084 6043 ne
tri 1084 5978 1147 6041 sw
rect 1084 5967 1147 5978
tri 1084 5904 1147 5967 ne
tri 1147 5904 1221 5978 sw
rect 3465 5976 3523 6834
tri 3523 6800 3557 6834 nw
tri 13115 6675 13389 6949 se
rect 13389 6675 13822 7374
tri 3619 6601 3659 6641 se
rect 3659 6601 4731 6641
rect 3619 6589 4731 6601
tri 3523 5976 3547 6000 sw
tri 1147 5830 1221 5904 ne
tri 1221 5830 1295 5904 sw
tri 3465 5894 3547 5976 ne
tri 3547 5936 3587 5976 sw
rect 3619 5946 3671 6589
tri 3671 6535 3725 6589 nw
tri 3764 6332 3798 6366 sw
tri 4242 6332 4303 6393 se
rect 4303 6341 4731 6393
rect 8847 6376 13822 6675
rect 4303 6332 4316 6341
tri 4316 6332 4325 6341 nw
rect 3764 6280 4264 6332
tri 4264 6280 4316 6332 nw
tri 3764 6249 3795 6280 nw
tri 4344 6249 4403 6308 se
rect 4403 6256 4731 6308
rect 4403 6249 4418 6256
tri 4418 6249 4425 6256 nw
rect 4023 6197 4366 6249
tri 4366 6197 4418 6249 nw
tri 3773 6169 3797 6193 sw
tri 4426 6169 4485 6228 se
rect 4485 6176 4731 6228
rect 4485 6169 4500 6176
tri 4500 6169 4507 6176 nw
rect 3773 6117 4448 6169
tri 4448 6117 4500 6169 nw
tri 4509 6117 4540 6148 se
rect 4540 6117 4731 6148
tri 3773 6075 3815 6117 nw
tri 4458 6066 4509 6117 se
rect 4509 6090 4731 6117
rect 4509 6066 4540 6090
tri 4540 6066 4564 6090 nw
tri 13089 6076 13389 6376 ne
tri 4451 6059 4458 6066 se
rect 4458 6059 4475 6066
rect 3894 6001 4475 6059
tri 4475 6001 4540 6066 nw
tri 3671 5946 3693 5968 sw
tri 3619 5936 3629 5946 ne
rect 3629 5936 3693 5946
rect 3547 5894 3587 5936
tri 3587 5894 3629 5936 sw
tri 3629 5894 3671 5936 ne
rect 3671 5894 3693 5936
tri 2857 5853 2881 5877 sw
tri 3547 5853 3588 5894 ne
rect 3588 5872 3629 5894
tri 3629 5872 3651 5894 sw
tri 3671 5872 3693 5894 ne
tri 3693 5872 3767 5946 sw
rect 3588 5854 3651 5872
tri 3651 5854 3669 5872 sw
tri 3693 5854 3711 5872 ne
rect 3711 5854 3767 5872
rect 3588 5853 3669 5854
tri 1221 5756 1295 5830 ne
tri 1295 5756 1369 5830 sw
rect 2857 5811 3532 5853
tri 3532 5811 3574 5853 sw
tri 3588 5811 3630 5853 ne
rect 3630 5812 3669 5853
tri 3669 5812 3711 5854 sw
tri 3711 5812 3753 5854 ne
rect 3753 5812 3767 5854
rect 3630 5811 3711 5812
rect 2857 5801 3574 5811
tri 2857 5767 2891 5801 nw
tri 405 5685 439 5719 sw
tri 1295 5704 1347 5756 ne
rect 1347 5704 1994 5756
tri 3510 5743 3568 5801 ne
rect 3568 5755 3574 5801
tri 3574 5755 3630 5811 sw
tri 3630 5755 3686 5811 ne
rect 3686 5798 3711 5811
tri 3711 5798 3725 5812 sw
tri 3753 5798 3767 5812 ne
tri 3767 5798 3841 5872 sw
rect 3686 5772 3725 5798
tri 3725 5772 3751 5798 sw
tri 3767 5772 3793 5798 ne
rect 3793 5772 3841 5798
rect 3686 5755 3751 5772
rect 3568 5743 3630 5755
tri 3426 5721 3448 5743 se
tri 3568 5681 3630 5743 ne
tri 3630 5730 3655 5755 sw
tri 3686 5730 3711 5755 ne
rect 3711 5730 3751 5755
tri 3751 5730 3793 5772 sw
tri 3793 5730 3835 5772 ne
rect 3835 5766 3841 5772
tri 3841 5766 3873 5798 sw
rect 3894 5787 3946 6001
tri 3946 5967 3980 6001 nw
tri 3946 5787 3968 5809 sw
tri 3894 5766 3915 5787 ne
rect 3915 5768 3968 5787
tri 3968 5768 3987 5787 sw
rect 4036 5768 4088 5943
rect 4571 5839 4703 5883
tri 4088 5768 4103 5783 sw
rect 3915 5766 3987 5768
rect 3835 5730 3873 5766
rect 3630 5681 3655 5730
tri 3655 5681 3704 5730 sw
tri 3711 5681 3760 5730 ne
rect 3760 5724 3793 5730
tri 3793 5724 3799 5730 sw
tri 3835 5724 3841 5730 ne
rect 3841 5724 3873 5730
tri 3873 5724 3915 5766 sw
tri 3915 5724 3957 5766 ne
rect 3957 5761 3987 5766
tri 3987 5761 3994 5768 sw
rect 4036 5761 4103 5768
rect 3957 5724 3994 5761
rect 3760 5690 3799 5724
tri 3799 5690 3833 5724 sw
tri 3841 5690 3875 5724 ne
rect 3875 5692 3915 5724
tri 3915 5692 3947 5724 sw
tri 3957 5692 3989 5724 ne
rect 3989 5719 3994 5724
tri 3994 5719 4036 5761 sw
tri 4036 5719 4078 5761 ne
rect 4078 5719 4103 5761
rect 3989 5694 4036 5719
tri 4036 5694 4061 5719 sw
tri 4078 5694 4103 5719 ne
tri 4103 5694 4177 5768 sw
tri 4571 5707 4703 5839 ne
tri 4703 5774 4783 5854 sw
rect 4703 5707 4783 5774
rect 3989 5692 4061 5694
rect 3875 5690 3947 5692
rect 3760 5681 3833 5690
tri 3383 5615 3448 5680 ne
rect 3448 5615 3451 5680
tri 3630 5607 3704 5681 ne
tri 3704 5648 3737 5681 sw
tri 3760 5648 3793 5681 ne
rect 3793 5648 3833 5681
tri 3833 5648 3875 5690 sw
tri 3875 5650 3915 5690 ne
rect 3915 5650 3947 5690
tri 3947 5650 3989 5692 sw
tri 3989 5650 4031 5692 ne
rect 4031 5652 4061 5692
tri 4061 5652 4103 5694 sw
tri 4103 5652 4145 5694 ne
rect 4145 5652 4177 5694
rect 4031 5650 4103 5652
rect 3704 5607 3737 5648
tri 3737 5607 3778 5648 sw
tri 3793 5607 3834 5648 ne
rect 3834 5608 3875 5648
tri 3875 5608 3915 5648 sw
tri 3915 5608 3957 5650 ne
rect 3957 5618 3989 5650
tri 3989 5618 4021 5650 sw
tri 4031 5618 4063 5650 ne
rect 4063 5620 4103 5650
tri 4103 5620 4135 5652 sw
tri 4145 5620 4177 5652 ne
tri 4177 5620 4251 5694 sw
rect 4541 5627 4688 5633
tri 4688 5627 4694 5633 sw
tri 4703 5627 4783 5707 ne
tri 4783 5627 4930 5774 sw
rect 4063 5618 4135 5620
rect 3957 5608 4021 5618
rect 3834 5607 3915 5608
tri 2897 5599 2904 5606 se
tri 3058 5599 3065 5606 sw
tri 3704 5533 3778 5607 ne
tri 3778 5566 3819 5607 sw
tri 3834 5566 3875 5607 ne
rect 3875 5566 3915 5607
tri 3915 5566 3957 5608 sw
tri 3957 5576 3989 5608 ne
rect 3989 5576 4021 5608
tri 4021 5576 4063 5618 sw
tri 4063 5576 4105 5618 ne
rect 4105 5578 4135 5618
tri 4135 5578 4177 5620 sw
tri 4177 5578 4219 5620 ne
rect 4219 5578 4251 5620
rect 4105 5576 4177 5578
tri 3989 5566 3999 5576 ne
rect 3999 5566 4063 5576
rect 3778 5533 3819 5566
tri 3819 5533 3852 5566 sw
tri 3875 5533 3908 5566 ne
rect 3908 5533 3957 5566
tri 1259 5435 1293 5469 sw
tri 3613 5463 3647 5497 nw
rect 3778 5479 3852 5533
tri 3852 5479 3906 5533 sw
tri 3908 5484 3957 5533 ne
tri 3957 5526 3997 5566 sw
tri 3999 5526 4039 5566 ne
rect 4039 5544 4063 5566
tri 4063 5544 4095 5576 sw
tri 4105 5544 4137 5576 ne
rect 4137 5546 4177 5576
tri 4177 5546 4209 5578 sw
tri 4219 5546 4251 5578 ne
tri 4251 5546 4325 5620 sw
rect 4541 5608 4694 5627
tri 4694 5608 4713 5627 sw
rect 4137 5544 4209 5546
rect 4039 5526 4095 5544
rect 3957 5484 3997 5526
tri 3997 5484 4039 5526 sw
tri 4039 5502 4063 5526 ne
rect 4063 5502 4095 5526
tri 4095 5502 4137 5544 sw
tri 4137 5502 4179 5544 ne
rect 4179 5504 4209 5544
tri 4209 5504 4251 5546 sw
tri 4251 5504 4293 5546 ne
rect 4293 5504 4325 5546
rect 4179 5502 4251 5504
tri 4063 5484 4081 5502 ne
rect 4081 5484 4137 5502
tri 3501 5351 3535 5385 se
tri 1426 5337 1439 5350 se
rect 3778 5346 3906 5479
tri 3957 5402 4039 5484 ne
tri 4039 5444 4079 5484 sw
tri 4081 5444 4121 5484 ne
rect 4121 5470 4137 5484
tri 4137 5470 4169 5502 sw
tri 4179 5470 4211 5502 ne
rect 4211 5472 4251 5502
tri 4251 5472 4283 5504 sw
tri 4293 5472 4325 5504 ne
tri 4325 5472 4399 5546 sw
rect 4541 5538 4713 5608
tri 4713 5538 4783 5608 sw
tri 4783 5538 4872 5627 ne
rect 4872 5538 4930 5627
rect 4541 5503 4783 5538
rect 4211 5470 4283 5472
rect 4121 5444 4169 5470
rect 4039 5402 4079 5444
tri 4079 5402 4121 5444 sw
tri 4121 5428 4137 5444 ne
rect 4137 5428 4169 5444
tri 4169 5428 4211 5470 sw
tri 4211 5428 4253 5470 ne
rect 4253 5430 4283 5470
tri 4283 5430 4325 5472 sw
tri 4325 5430 4367 5472 ne
rect 4367 5430 4399 5472
rect 4253 5428 4325 5430
tri 4137 5402 4163 5428 ne
rect 4163 5402 4211 5428
tri 4039 5320 4121 5402 ne
tri 4121 5362 4161 5402 sw
tri 4163 5362 4203 5402 ne
rect 4203 5396 4211 5402
tri 4211 5396 4243 5428 sw
tri 4253 5396 4285 5428 ne
rect 4285 5398 4325 5428
tri 4325 5398 4357 5430 sw
tri 4367 5398 4399 5430 ne
tri 4399 5398 4473 5472 sw
tri 4634 5431 4706 5503 ne
rect 4706 5480 4783 5503
tri 4783 5480 4841 5538 sw
tri 4872 5480 4930 5538 ne
tri 4930 5480 5077 5627 sw
tri 5473 5480 5592 5599 se
rect 5592 5480 5646 5660
rect 4706 5431 4841 5480
tri 4841 5431 4890 5480 sw
rect 4285 5396 4357 5398
rect 4203 5362 4243 5396
rect 4121 5320 4161 5362
tri 4161 5320 4203 5362 sw
tri 4203 5354 4211 5362 ne
rect 4211 5354 4243 5362
tri 4243 5354 4285 5396 sw
tri 4285 5354 4327 5396 ne
rect 4327 5356 4357 5396
tri 4357 5356 4399 5398 sw
tri 4399 5356 4441 5398 ne
rect 4441 5356 4473 5398
rect 4327 5354 4399 5356
tri 4211 5320 4245 5354 ne
rect 4245 5322 4285 5354
tri 4285 5322 4317 5354 sw
tri 4327 5322 4359 5354 ne
rect 4359 5324 4399 5354
tri 4399 5324 4431 5356 sw
tri 4441 5324 4473 5356 ne
tri 4473 5324 4547 5398 sw
rect 4359 5322 4431 5324
rect 4245 5320 4317 5322
tri 1426 5298 1439 5311 ne
rect 1439 5298 1440 5311
tri 1456 5264 1490 5298 ne
tri 1518 5264 1552 5298 nw
tri 3929 5252 3932 5255 se
tri 4121 5238 4203 5320 ne
tri 4203 5280 4243 5320 sw
tri 4245 5280 4285 5320 ne
rect 4285 5280 4317 5320
tri 4317 5280 4359 5322 sw
tri 4359 5280 4401 5322 ne
rect 4401 5282 4431 5322
tri 4431 5282 4473 5324 sw
tri 4473 5282 4515 5324 ne
rect 4515 5282 4547 5324
rect 4401 5280 4473 5282
rect 4203 5238 4243 5280
tri 4243 5238 4285 5280 sw
tri 4285 5238 4327 5280 ne
rect 4327 5248 4359 5280
tri 4359 5248 4391 5280 sw
tri 4401 5248 4433 5280 ne
rect 4433 5250 4473 5280
tri 4473 5250 4505 5282 sw
tri 4515 5250 4547 5282 ne
tri 4547 5250 4621 5324 sw
rect 4433 5248 4505 5250
rect 4327 5238 4391 5248
tri -744 5165 -710 5199 nw
tri 3907 5175 3932 5200 ne
tri 3043 5156 3044 5157 sw
tri 4203 5156 4285 5238 ne
tri 4285 5199 4324 5238 sw
tri 4327 5199 4366 5238 ne
rect 4366 5206 4391 5238
tri 4391 5206 4433 5248 sw
tri 4433 5206 4475 5248 ne
rect 4475 5208 4505 5248
tri 4505 5208 4547 5250 sw
tri 4547 5208 4589 5250 ne
rect 4589 5208 4621 5250
rect 4475 5206 4547 5208
rect 4366 5199 4433 5206
rect 4285 5157 4324 5199
tri 4324 5157 4366 5199 sw
tri 4366 5157 4408 5199 ne
rect 4408 5174 4433 5199
tri 4433 5174 4465 5206 sw
tri 4475 5174 4507 5206 ne
rect 4507 5176 4547 5206
tri 4547 5176 4579 5208 sw
tri 4589 5176 4621 5208 ne
tri 4621 5176 4695 5250 sw
tri 4706 5247 4890 5431 ne
tri 4890 5391 4930 5431 sw
tri 4930 5391 5019 5480 ne
rect 5019 5469 5646 5480
tri 5646 5469 5837 5660 nw
tri 9172 5653 9422 5903 se
rect 9422 5653 10200 5903
tri 6172 5615 6210 5653 se
rect 6210 5615 10200 5653
tri 6026 5469 6172 5615 se
rect 6172 5523 10200 5615
rect 13389 5608 13822 6376
rect 6172 5469 6210 5523
tri 6210 5469 6264 5523 nw
rect 5019 5391 5527 5469
rect 4890 5350 4930 5391
tri 4930 5350 4971 5391 sw
tri 5019 5350 5060 5391 ne
rect 5060 5350 5527 5391
tri 5527 5350 5646 5469 nw
rect 4890 5247 4971 5350
tri 4971 5247 5074 5350 sw
tri 5842 5285 6026 5469 se
tri 6026 5285 6210 5469 nw
tri 5804 5247 5842 5285 se
rect 5842 5247 5858 5285
rect 4507 5174 4579 5176
rect 4408 5157 4465 5174
rect 4285 5156 4366 5157
tri 1207 5131 1221 5145 ne
tri 1249 5135 1259 5145 nw
tri 1407 5118 1410 5121 ne
tri 1433 5095 1459 5121 nw
tri 1685 5040 1759 5114 se
rect 1759 5062 2154 5114
tri 3818 5071 3852 5105 ne
tri 4285 5075 4366 5156 ne
tri 4366 5132 4391 5157 sw
tri 4408 5132 4433 5157 ne
rect 4433 5132 4465 5157
tri 4465 5132 4507 5174 sw
tri 4507 5132 4549 5174 ne
rect 4549 5134 4579 5174
tri 4579 5134 4621 5176 sw
tri 4621 5134 4663 5176 ne
rect 4663 5134 4695 5176
rect 4549 5132 4621 5134
rect 4366 5099 4391 5132
tri 4391 5099 4424 5132 sw
tri 4433 5102 4463 5132 ne
rect 4463 5131 4507 5132
tri 4507 5131 4508 5132 sw
tri 1759 5040 1781 5062 nw
tri 1651 5006 1685 5040 se
rect 1685 5006 1703 5040
tri -227 4654 -225 4656 se
tri -458 4612 -438 4632 ne
tri -412 4626 -406 4632 nw
tri -334 4601 -306 4629 nw
tri -660 4417 -631 4446 nw
tri 328 3878 362 3912 se
tri 272 3794 304 3826 ne
tri 356 3792 390 3826 nw
rect 1651 3708 1703 5006
tri 1703 4984 1759 5040 nw
tri 1953 4821 1973 4841 ne
tri 1703 3708 1725 3730 sw
tri 1651 3634 1725 3708 ne
tri 1725 3634 1799 3708 sw
tri 1725 3560 1799 3634 ne
tri 1799 3560 1873 3634 sw
tri 1799 3502 1857 3560 ne
rect 1857 3524 1873 3560
tri 1873 3524 1909 3560 sw
tri 1466 3339 1490 3363 se
rect 1857 3301 1909 3524
rect 1973 3266 2025 4841
tri 2025 4785 2081 4841 nw
tri 4083 4838 4100 4855 se
tri 4074 4760 4100 4786 ne
tri 2649 4640 2683 4674 ne
tri 3977 4671 4011 4705 ne
tri 4281 4468 4302 4489 ne
tri 4123 4188 4157 4222 se
tri 2812 4075 2846 4109 sw
tri 4123 4075 4157 4109 se
tri 4128 3994 4157 4023 ne
tri 2649 3915 2683 3949 se
tri 2711 3915 2745 3949 sw
rect 4302 3948 4334 4617
rect 4366 4288 4424 5099
tri 4334 3948 4368 3982 sw
tri 4123 3877 4157 3911 se
tri 4438 3864 4463 3889 se
rect 4463 3864 4508 5131
tri 4549 5102 4579 5132 ne
rect 4579 5102 4621 5132
tri 4621 5102 4653 5134 sw
tri 4663 5102 4695 5134 ne
tri 4695 5102 4769 5176 sw
tri 4890 5117 5020 5247 ne
rect 5020 5117 5858 5247
tri 5858 5117 6026 5285 nw
tri 4579 5053 4628 5102 ne
rect 4628 5075 4653 5102
tri 4653 5075 4680 5102 sw
tri 4695 5080 4717 5102 ne
tri 4140 3836 4157 3853 ne
rect 4157 3836 4160 3853
rect 4264 3815 4508 3864
tri 4163 3719 4176 3732 se
tri 4142 3657 4176 3691 ne
tri 2116 3567 2190 3641 se
rect 2190 3611 3939 3641
tri 3939 3611 3969 3641 sw
rect 2190 3589 3969 3611
tri 2190 3567 2212 3589 nw
tri 2092 3543 2116 3567 se
rect 2116 3543 2144 3567
tri 273 2989 304 3020 se
tri 356 2989 390 3023 sw
tri -655 2955 -621 2989 sw
tri -655 2869 -621 2903 nw
tri 2078 2671 2092 2685 se
rect 2092 2671 2144 3543
tri 2144 3521 2190 3567 nw
tri 3917 3537 3969 3589 ne
tri 3969 3537 4043 3611 sw
tri 4221 3537 4264 3580 se
rect 4264 3537 4316 3815
tri 4316 3781 4350 3815 nw
tri 4395 3571 4407 3583 ne
tri 4434 3570 4447 3583 nw
tri 2241 3495 2282 3536 se
rect 2282 3495 3861 3536
tri 3861 3495 3902 3536 sw
tri 2191 3445 2241 3495 se
rect 2241 3485 3902 3495
tri 3902 3485 3912 3495 sw
tri 3969 3485 4021 3537 ne
rect 4021 3515 4316 3537
rect 4021 3485 4286 3515
tri 4286 3485 4316 3515 nw
tri 4482 3527 4537 3582 se
rect 4537 3560 4589 4416
rect 4537 3527 4556 3560
tri 4556 3527 4589 3560 nw
rect 2241 3484 3912 3485
rect 2241 3445 2243 3484
rect 2191 3301 2243 3445
tri 2243 3423 2304 3484 nw
tri 3839 3421 3902 3484 ne
rect 3902 3421 3912 3484
tri 3912 3421 3976 3485 sw
tri 4151 3421 4176 3446 se
tri 3902 3369 3954 3421 ne
rect 3954 3372 4176 3421
rect 3954 3369 4177 3372
tri 4125 3318 4176 3369 ne
rect 4176 3318 4177 3369
tri 3493 3094 3527 3128 sw
tri 4142 3094 4176 3128 se
tri 4134 3000 4176 3042 ne
tri 3431 2914 3458 2941 sw
tri 4143 2914 4176 2947 se
tri 3186 2894 3190 2898 se
tri 3234 2894 3238 2898 sw
tri 3287 2829 3306 2848 ne
tri 3333 2842 3339 2848 nw
tri 3431 2828 3465 2862 nw
tri 4133 2819 4176 2862 ne
rect 1627 2618 1679 2671
tri 1627 2566 1679 2618 ne
tri 1679 2600 1719 2640 sw
tri 2007 2600 2078 2671 se
rect 2078 2663 2144 2671
rect 2078 2600 2081 2663
tri 2081 2600 2144 2663 nw
rect 1679 2566 2029 2600
tri 1679 2548 1697 2566 ne
rect 1697 2548 2029 2566
tri 2029 2548 2081 2600 nw
tri 4095 2394 4176 2475 se
rect 2882 2313 3052 2364
tri 3052 2313 3103 2364 sw
tri 4157 2347 4176 2366 ne
rect 2882 2312 4265 2313
tri 3030 2261 3081 2312 ne
rect 3081 2261 4265 2312
tri 1512 1987 1546 2021 se
tri 1598 1987 1630 2019 sw
rect 4482 1957 4534 3527
tri 4534 3505 4556 3527 nw
tri 4562 3404 4628 3470 se
rect 4628 3448 4680 5075
rect 4628 3404 4636 3448
tri 4636 3404 4680 3448 nw
tri 3264 1847 3275 1858 ne
rect 3275 1847 3277 1858
rect 3426 1847 3435 1858
tri 3435 1847 3446 1858 nw
tri 705 1466 739 1500 ne
tri 767 1475 792 1500 nw
tri 2388 1351 2398 1361 ne
tri 2436 1327 2470 1361 nw
tri 2864 1340 2888 1364 ne
tri 2915 1330 2949 1364 nw
tri 549 1150 562 1163 se
tri 613 1150 647 1184 sw
tri -267 1006 -233 1040 sw
tri -217 556 -174 599 se
tri -124 556 -89 591 sw
tri -399 489 -389 499 se
tri -361 489 -347 503 sw
tri -188 470 -154 504 ne
rect -128 473 -124 504
tri -128 469 -124 473 ne
tri -124 469 -89 504 nw
tri 4211 413 4245 447 se
rect 4562 392 4614 3404
tri 4614 3382 4636 3404 nw
rect 4717 2947 4769 5102
rect 11453 4703 11985 4989
tri 11985 4703 12271 4989 sw
rect 11453 4661 13156 4703
tri 13156 4661 13198 4703 sw
rect 11453 4650 13833 4661
tri 13135 4609 13176 4650 ne
rect 13176 4648 13833 4650
tri 13833 4648 13846 4661 sw
rect 13176 4609 13846 4648
tri 13811 4574 13846 4609 ne
tri 13846 4574 13920 4648 sw
tri 5513 4558 5516 4561 se
rect 5516 4558 13553 4561
tri 13553 4558 13556 4561 sw
tri 5476 4521 5513 4558 se
rect 5513 4533 13556 4558
rect 5513 4521 5516 4533
tri 5516 4521 5528 4533 nw
tri 5436 4481 5476 4521 se
tri 5476 4481 5516 4521 nw
tri 5516 4481 5540 4505 se
rect 5540 4481 12584 4505
tri 5396 4441 5436 4481 se
tri 5436 4441 5476 4481 nw
tri 5500 4465 5516 4481 se
rect 5516 4477 12584 4481
rect 5516 4465 5524 4477
tri 5476 4441 5500 4465 se
rect 5500 4449 5524 4465
tri 5524 4449 5552 4477 nw
tri 12558 4451 12584 4477 ne
tri 12584 4470 12619 4505 sw
tri 13527 4504 13556 4533 ne
tri 13556 4504 13610 4558 sw
tri 13846 4552 13868 4574 ne
rect 12584 4451 12619 4470
tri 5394 4439 5396 4441 se
rect 5396 4439 5422 4441
tri 5087 4324 5121 4358 ne
rect 5121 3891 5173 4387
tri 5173 4328 5203 4358 nw
tri 5276 3920 5310 3954 ne
tri 5173 3891 5192 3910 sw
rect 5121 3888 5192 3891
tri 5121 3817 5192 3888 ne
tri 5192 3817 5266 3891 sw
tri 5192 3795 5214 3817 ne
tri 5138 2313 5214 2389 se
rect 5214 2313 5266 3817
rect 5394 1372 5422 4439
tri 5422 4427 5436 4441 nw
tri 5450 4415 5476 4441 se
rect 5476 4425 5500 4441
tri 5500 4425 5524 4449 nw
rect 5476 4415 5478 4425
rect 5450 3365 5478 4415
tri 5478 4403 5500 4425 nw
tri 6433 4410 6472 4449 se
rect 6472 4419 11174 4449
tri 11174 4419 11204 4449 sw
tri 12584 4444 12591 4451 ne
rect 6472 4411 11204 4419
rect 6472 4410 6480 4411
rect 5780 4383 6480 4410
tri 6480 4383 6508 4411 nw
rect 5780 4358 6455 4383
tri 6455 4358 6480 4383 nw
tri 6543 4333 6593 4383 se
rect 6593 4370 10277 4383
tri 10277 4370 10290 4383 sw
rect 6593 4347 10290 4370
tri 6593 4333 6607 4347 nw
tri 6493 4283 6543 4333 se
tri 6543 4283 6593 4333 nw
tri 10239 4296 10290 4347 ne
tri 10290 4296 10364 4370 sw
tri 11158 4365 11204 4411 ne
tri 11204 4365 11258 4419 sw
tri 11204 4349 11220 4365 ne
tri 6443 4233 6493 4283 se
tri 6493 4233 6543 4283 nw
tri 10290 4274 10312 4296 ne
tri 6398 4188 6443 4233 se
rect 6443 4188 6448 4233
tri 6448 4188 6493 4233 nw
rect 10312 4196 10364 4296
tri 10364 4196 10398 4230 sw
tri 6106 4138 6156 4188 se
rect 6156 4160 6420 4188
tri 6420 4160 6448 4188 nw
rect 11220 4185 11258 4365
tri 6156 4138 6178 4160 nw
tri 11220 4147 11258 4185 ne
tri 11258 4156 11303 4201 sw
rect 11258 4147 11303 4156
tri 6070 4102 6106 4138 se
rect 6106 4102 6120 4138
tri 6120 4102 6156 4138 nw
tri 6877 4106 6911 4140 nw
tri 9816 4110 9850 4144 ne
tri 9895 4125 9914 4144 nw
tri 11258 4102 11303 4147 ne
tri 11303 4102 11357 4156 sw
tri 5546 4028 5620 4102 se
rect 5620 4066 6084 4102
tri 6084 4066 6120 4102 nw
tri 5620 4028 5658 4066 nw
tri 11303 4048 11357 4102 ne
tri 11357 4048 11411 4102 sw
tri 5536 4018 5546 4028 se
rect 5546 4018 5588 4028
tri 5478 3493 5502 3517 sw
tri 5462 3088 5536 3162 se
rect 5536 3140 5588 4018
tri 5588 3996 5620 4028 nw
tri 7023 3970 7057 4004 ne
tri 7073 3969 7108 4004 nw
tri 9443 3975 9477 4009 se
tri 9505 3975 9539 4009 sw
tri 11357 3994 11411 4048 ne
tri 11411 3994 11465 4048 sw
tri 9816 3940 9850 3974 se
tri 9898 3940 9932 3974 sw
tri 9977 3939 10002 3964 se
tri 10054 3939 10088 3973 sw
tri 10200 3921 10234 3955 sw
tri 10874 3921 10908 3955 se
tri 11411 3940 11465 3994 ne
tri 11465 3940 11519 3994 sw
tri 5619 3856 5655 3892 ne
tri 5692 3837 5747 3892 nw
tri 11465 3886 11519 3940 ne
tri 11519 3886 11573 3940 sw
tri 11519 3832 11573 3886 ne
tri 11573 3832 11627 3886 sw
tri 11573 3778 11627 3832 ne
tri 11627 3778 11681 3832 sw
tri 11627 3724 11681 3778 ne
tri 11681 3724 11735 3778 sw
tri 8050 3649 8084 3683 ne
tri 8111 3649 8145 3683 nw
rect 10712 3554 11373 3678
tri 11373 3554 11497 3678 sw
tri 11681 3670 11735 3724 ne
tri 11735 3670 11789 3724 sw
tri 11735 3616 11789 3670 ne
tri 11789 3616 11843 3670 sw
tri 11789 3562 11843 3616 ne
tri 11843 3562 11897 3616 sw
tri 5826 3428 5860 3462 nw
tri 11259 3316 11497 3554 ne
tri 11497 3316 11735 3554 sw
tri 11843 3546 11859 3562 ne
tri 11497 3261 11552 3316 ne
rect 11552 3305 11735 3316
tri 11735 3305 11746 3316 sw
tri 6464 3159 6512 3207 se
tri 6555 3159 6592 3196 sw
tri 5536 3088 5588 3140 nw
rect 5462 1589 5514 3088
tri 5514 3066 5536 3088 nw
tri 5640 2865 5653 2878 se
tri 6402 2863 6436 2897 sw
tri 8815 2863 8849 2897 se
tri 8899 2863 8921 2885 sw
tri 5684 2794 5703 2813 nw
tri 6423 2718 6457 2752 ne
tri 8912 2456 8946 2490 ne
tri 8974 2456 9008 2490 nw
tri 9222 2379 9246 2403 sw
rect 11552 2376 11746 3305
rect 11859 2519 11897 3562
rect 12591 3508 12619 4451
tri 13556 4450 13610 4504 ne
tri 13610 4450 13664 4504 sw
tri 13610 4396 13664 4450 ne
tri 13664 4396 13718 4450 sw
tri 13664 4342 13718 4396 ne
tri 13718 4342 13772 4396 sw
tri 13718 4340 13720 4342 ne
rect 13720 4097 13772 4342
rect 13061 3928 13220 3951
tri 13220 3928 13243 3951 sw
rect 13868 3928 13920 4574
rect 14063 3950 14115 8512
rect 13061 3899 13549 3928
tri 13162 3800 13261 3899 ne
rect 13261 3800 13549 3899
rect 13061 3684 13227 3709
tri 13227 3684 13252 3709 sw
rect 13061 3657 13742 3684
tri 13205 3632 13230 3657 ne
rect 13230 3632 13742 3657
tri 14069 3621 14143 3695 se
tri 14143 3621 14173 3651 nw
tri 14052 3604 14069 3621 se
rect 14069 3604 14076 3621
rect 13052 3554 14076 3604
tri 14076 3554 14143 3621 nw
rect 13052 3552 14074 3554
tri 14074 3552 14076 3554 nw
tri 12591 3480 12619 3508 ne
tri 12619 3480 12668 3529 sw
tri 14101 3520 14135 3554 se
tri 12619 3431 12668 3480 ne
tri 12668 3431 12717 3480 sw
rect 13165 3468 14135 3520
tri 13165 3434 13199 3468 nw
tri 14108 3441 14135 3468 ne
tri 12668 3403 12696 3431 ne
rect 12696 3403 12940 3431
tri 12910 3373 12940 3403 ne
tri 12940 3375 12996 3431 sw
rect 12940 3373 12996 3375
tri 12940 3317 12996 3373 ne
tri 12996 3317 13054 3375 sw
rect 12064 3101 12888 3294
tri 12888 3292 12890 3294 sw
tri 12913 3259 12946 3292 sw
tri 12996 3259 13054 3317 ne
tri 13054 3259 13112 3317 sw
tri 14133 3302 14167 3336 ne
rect 12913 3201 12946 3259
tri 12946 3201 13004 3259 sw
tri 13054 3201 13112 3259 ne
tri 13112 3201 13170 3259 sw
rect 12913 3101 13004 3201
tri 13004 3101 13104 3201 sw
tri 13112 3149 13164 3201 ne
rect 13164 3149 13474 3201
tri 13700 3124 13850 3274 se
tri 13637 3101 13660 3124 se
rect 13660 3101 13953 3124
rect 12064 3017 13953 3101
tri 13984 3077 14011 3104 se
rect 14011 3077 14056 3152
tri 14056 3118 14090 3152 nw
rect 13984 3069 14056 3077
rect 12064 2995 13681 3017
tri 13681 2995 13703 3017 nw
tri 11859 2481 11897 2519 ne
tri 11897 2497 11935 2535 sw
rect 12064 2497 12888 2995
tri 12888 2826 13057 2995 nw
tri 13902 2800 13984 2882 se
rect 13984 2800 14030 3069
tri 14030 3043 14056 3069 nw
tri 14133 3025 14167 3059 se
rect 13114 2700 13579 2756
tri 13493 2614 13579 2700 ne
tri 13579 2622 13713 2756 sw
rect 13579 2614 13716 2622
tri 13579 2570 13623 2614 ne
rect 13623 2570 13716 2614
rect 11897 2481 11935 2497
tri 11897 2452 11926 2481 ne
rect 11926 2452 11935 2481
tri 11935 2452 11980 2497 sw
tri 11926 2398 11980 2452 ne
tri 11980 2398 12034 2452 sw
rect 13105 2398 13463 2463
tri 9393 2284 9432 2323 se
rect 9432 2284 9645 2323
tri 9662 2317 9696 2351 ne
tri 11980 2344 12034 2398 ne
tri 12034 2344 12088 2398 sw
tri 12034 2306 12072 2344 ne
rect 12072 2306 13337 2344
tri 13321 2290 13337 2306 ne
tri 13337 2300 13381 2344 sw
tri 13402 2337 13463 2398 ne
tri 13463 2382 13544 2463 sw
rect 13463 2337 13544 2382
rect 13337 2290 13381 2300
tri 8899 2218 8946 2265 se
tri 8974 2218 9008 2252 sw
rect 9311 2128 9645 2284
tri 13337 2246 13381 2290 ne
tri 13381 2246 13435 2300 sw
tri 13463 2256 13544 2337 ne
tri 13544 2256 13670 2382 sw
tri 13381 2192 13435 2246 ne
tri 13435 2192 13489 2246 sw
tri 5703 2041 5737 2075 sw
rect 9311 2051 9435 2128
tri 9090 2045 9094 2049 ne
rect 9094 2045 9096 2049
rect 9302 2046 9435 2051
tri 9435 2046 9517 2128 nw
tri 9689 2125 9697 2133 se
tri 9724 2125 9758 2159 sw
tri 13435 2138 13489 2192 ne
tri 13489 2138 13543 2192 sw
tri 13489 2084 13543 2138 ne
tri 13543 2137 13544 2138 sw
tri 13544 2137 13663 2256 ne
rect 13663 2137 13670 2256
rect 13543 2084 13544 2137
tri 13544 2084 13597 2137 sw
tri 13663 2130 13670 2137 ne
tri 13670 2130 13796 2256 sw
tri 13670 2094 13706 2130 ne
tri 13543 2082 13545 2084 ne
rect 13545 2052 13597 2084
rect 9302 2045 9311 2046
tri 9311 2045 9312 2046 nw
tri 5872 1955 5906 1989 ne
tri 5726 1810 5752 1836 ne
tri 5802 1802 5836 1836 nw
tri 8600 1796 8634 1830 ne
tri 7744 1755 7778 1789 ne
rect 12709 1687 12764 1702
rect 12709 1681 12768 1687
tri 12722 1635 12768 1681 ne
tri 5514 1589 5543 1618 sw
tri 5422 1502 5446 1526 sw
tri 7830 1492 7864 1526 sw
tri 8686 1471 8720 1505 sw
tri 8769 1471 8797 1499 se
tri 8763 1385 8797 1419 ne
tri 10792 1339 10950 1497 se
rect 10950 1348 12172 1497
rect 10950 1339 10973 1348
rect 9771 1159 10973 1339
tri 10973 1159 11162 1348 nw
tri 12089 1265 12172 1348 ne
tri 12172 1339 12330 1497 sw
rect 12172 1265 12717 1339
tri 5872 1053 5906 1087 se
tri 12172 1082 12355 1265 ne
rect 12355 1082 12717 1265
tri 12734 1047 12768 1081 se
tri 5872 967 5906 1001 ne
tri 6974 810 7008 844 nw
tri 6810 753 6844 787 ne
tri 6865 751 6901 787 nw
tri 6587 713 6621 747 ne
tri 7150 685 7170 705 sw
tri 7554 686 7560 692 se
tri 7547 640 7560 653 ne
tri 7132 576 7154 598 nw
rect 13706 521 13796 2130
tri 9974 390 10012 428 se
tri 10036 390 10102 456 sw
tri 10846 421 10880 455 sw
tri 8515 378 8527 390 se
rect 8527 378 8528 390
tri -399 351 -389 361 ne
tri -361 347 -347 361 nw
tri 4373 333 4407 367 se
tri 8513 338 8527 352 ne
tri 11089 334 11123 368 se
tri 3766 277 3800 311 se
tri 3823 277 3857 311 sw
tri 7636 266 7660 290 ne
rect 7660 266 7662 290
tri 10636 230 10670 264 ne
tri 10722 217 10756 251 sw
tri 11196 -154 11304 -46 se
rect 11304 -102 11356 499
tri 11304 -154 11356 -102 nw
tri 11189 -161 11196 -154 se
rect 11196 -161 11245 -154
tri 8864 -235 8938 -161 se
rect 8938 -213 11245 -161
tri 11245 -213 11304 -154 nw
tri 8938 -235 8960 -213 nw
tri 8861 -238 8864 -235 se
rect 8864 -238 8913 -235
tri 426 -413 436 -403 se
tri 464 -413 478 -399 sw
rect 8861 -406 8913 -238
tri 8913 -260 8938 -235 nw
tri 8913 -406 8935 -384 sw
tri -176 -448 -154 -426 se
tri 8861 -480 8935 -406 ne
tri 8935 -480 9009 -406 sw
tri 8935 -502 8957 -480 ne
tri 8883 -2183 8957 -2109 se
rect 8957 -2131 9009 -480
tri 8957 -2183 9009 -2131 nw
tri 8809 -2257 8883 -2183 se
tri 8883 -2257 8957 -2183 nw
tri 8711 -2355 8809 -2257 se
rect 8809 -2355 8839 -2257
tri 8839 -2301 8883 -2257 nw
rect 8711 -2381 8839 -2355
<< metal3 >>
tri 908 3636 998 3726 se
rect 998 3636 1064 6904
tri 1054 2462 1124 2532 se
rect 1124 2462 1190 8728
tri 6285 6779 6474 6968 se
rect 6474 6783 6951 7493
tri 6951 7318 7126 7493 nw
rect 6474 6779 6754 6783
tri 1190 2462 1195 2467 sw
rect 6285 360 6754 6779
tri 6754 6586 6951 6783 nw
tri 9271 4912 9426 5067 ne
rect 9426 -592 9895 5067
tri 9895 4893 10069 5067 nw
tri 12570 4104 13014 4548 se
rect 13014 4396 13308 5783
rect 13014 4104 13016 4396
tri 13016 4104 13308 4396 nw
tri 10341 -7548 10347 -7542 se
rect 10347 -8480 10711 3059
rect 12068 1047 12884 4104
tri 12884 3972 13016 4104 nw
use sky130_fd_io__amux_switch_1v2b  sky130_fd_io__amux_switch_1v2b_0
timestamp 1676037725
transform 1 0 4755 0 -1 8802
box -50 -73 10379 2429
use sky130_fd_io__amux_switch_1v2b  sky130_fd_io__amux_switch_1v2b_1
timestamp 1676037725
transform 1 0 4755 0 1 4180
box -50 -73 10379 2429
use sky130_fd_io__gpiov2_amux_ctl_logic  sky130_fd_io__gpiov2_amux_ctl_logic_0
timestamp 1676037725
transform 1 0 -26998 0 1 6306
box 26021 -16454 41918 1960
use sky130_fd_io__res75only_small  sky130_fd_io__res75only_small_0
timestamp 1676037725
transform 1 0 3419 0 -1 6879
box 0 0 882 404
use sky130_fd_io__res75only_small  sky130_fd_io__res75only_small_1
timestamp 1676037725
transform 1 0 2619 0 -1 6379
box 0 0 882 404
use sky130_fd_io__res75only_small  sky130_fd_io__res75only_small_2
timestamp 1676037725
transform 1 0 2619 0 -1 6879
box 0 0 882 404
use sky130_fd_io__res75only_small  sky130_fd_io__res75only_small_3
timestamp 1676037725
transform 1 0 3419 0 -1 6379
box 0 0 882 404
use sky130_fd_io__res75only_small  sky130_fd_io__res75only_small_4
timestamp 1676037725
transform -1 0 8708 0 1 9409
box 0 0 882 404
use sky130_fd_io__res75only_small  sky130_fd_io__res75only_small_5
timestamp 1676037725
transform 1 0 8626 0 1 9409
box 0 0 882 404
use sky130_fd_io__res75only_small  sky130_fd_io__res75only_small_6
timestamp 1676037725
transform 0 1 12464 1 0 3136
box 0 0 882 404
use sky130_fd_io__res75only_small  sky130_fd_io__res75only_small_7
timestamp 1676037725
transform 0 -1 12368 1 0 3136
box 0 0 882 404
use sky130_fd_io__res75only_small  sky130_fd_io__res75only_small_8
timestamp 1676037725
transform 0 1 12464 -1 0 3218
box 0 0 882 404
use sky130_fd_io__res75only_small  sky130_fd_io__res75only_small_9
timestamp 1676037725
transform 0 -1 11869 1 0 3136
box 0 0 882 404
use sky130_fd_io__res75only_small  sky130_fd_io__res75only_small_10
timestamp 1676037725
transform -1 0 1901 0 -1 6879
box 0 0 882 404
use sky130_fd_io__res75only_small  sky130_fd_io__res75only_small_11
timestamp 1676037725
transform -1 0 2701 0 -1 6879
box 0 0 882 404
use sky130_fd_io__res75only_small  sky130_fd_io__res75only_small_12
timestamp 1676037725
transform -1 0 2701 0 -1 6379
box 0 0 882 404
use sky130_fd_io__res75only_small  sky130_fd_io__res75only_small_13
timestamp 1676037725
transform -1 0 1901 0 -1 6379
box 0 0 882 404
use sky130_fd_pr__nfet_01v8__example_55959141808592  sky130_fd_pr__nfet_01v8__example_55959141808592_0
timestamp 1676037725
transform 1 0 14424 0 1 3035
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808592  sky130_fd_pr__nfet_01v8__example_55959141808592_1
timestamp 1676037725
transform 1 0 13880 0 1 3035
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808592  sky130_fd_pr__nfet_01v8__example_55959141808592_2
timestamp 1676037725
transform 1 0 13608 0 1 3035
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808592  sky130_fd_pr__nfet_01v8__example_55959141808592_3
timestamp 1676037725
transform 1 0 14152 0 1 3035
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808592  sky130_fd_pr__nfet_01v8__example_55959141808592_4
timestamp 1676037725
transform 1 0 13608 0 -1 3321
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808592  sky130_fd_pr__nfet_01v8__example_55959141808592_5
timestamp 1676037725
transform 1 0 14152 0 -1 3321
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808592  sky130_fd_pr__nfet_01v8__example_55959141808592_6
timestamp 1676037725
transform 1 0 14424 0 -1 3321
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808592  sky130_fd_pr__nfet_01v8__example_55959141808592_7
timestamp 1676037725
transform 1 0 13880 0 -1 3321
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808593  sky130_fd_pr__nfet_01v8__example_55959141808593_0
timestamp 1676037725
transform 1 0 13603 0 1 3415
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808593  sky130_fd_pr__nfet_01v8__example_55959141808593_1
timestamp 1676037725
transform 1 0 14151 0 1 3415
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808593  sky130_fd_pr__nfet_01v8__example_55959141808593_2
timestamp 1676037725
transform 1 0 14423 0 1 3415
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808593  sky130_fd_pr__nfet_01v8__example_55959141808593_3
timestamp 1676037725
transform 1 0 13875 0 1 3415
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808594  sky130_fd_pr__nfet_01v8__example_55959141808594_0
timestamp 1676037725
transform 0 -1 14630 -1 0 2528
box -1 0 2129 1
use sky130_fd_pr__pfet_01v8__example_55959141808591  sky130_fd_pr__pfet_01v8__example_55959141808591_0
timestamp 1676037725
transform 0 1 1282 -1 0 8427
box -1 0 1037 1
<< properties >>
string GDS_END 44785602
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 44268844
<< end >>
