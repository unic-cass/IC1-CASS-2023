magic
tech sky130A
magscale 1 2
timestamp 1676037725
<< locali >>
rect 0 1397 846 1431
rect 430 724 464 1167
rect 430 690 559 724
rect 657 690 691 724
rect 345 485 379 551
rect 212 361 246 427
rect 79 237 113 303
rect 0 -17 846 17
use pdriver_3  pdriver_3_0
timestamp 1676037725
transform 1 0 478 0 1 0
box -36 -17 404 1471
use pnand3  pnand3_0
timestamp 1676037725
transform 1 0 0 0 1 0
box -36 -17 514 1471
<< labels >>
rlabel locali s 674 707 674 707 4 Z
port 4 nsew
rlabel locali s 423 1414 423 1414 4 vdd
port 5 nsew
rlabel locali s 423 0 423 0 4 gnd
port 6 nsew
rlabel locali s 96 270 96 270 4 A
port 1 nsew
rlabel locali s 362 518 362 518 4 C
port 3 nsew
rlabel locali s 229 394 229 394 4 B
port 2 nsew
<< properties >>
string FIXED_BBOX 0 0 846 1414
string GDS_END 5257658
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sram_1rw1r_32_256_8_sky130.gds
string GDS_START 5256418
<< end >>
