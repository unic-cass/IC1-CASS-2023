VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO R4_butter
  CLASS BLOCK ;
  FOREIGN R4_butter ;
  ORIGIN 0.000 0.000 ;
  SIZE 182.000 BY 194.000 ;
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.030 0.000 179.310 4.000 ;
    END
  END CLK
  PIN RST
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.000 168.680 182.000 169.280 ;
    END
  END RST
  PIN Xio[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.830 0.000 124.110 4.000 ;
    END
  END Xio[0]
  PIN Xio[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.190 0.000 131.470 4.000 ;
    END
  END Xio[1]
  PIN Xio[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 0.000 138.830 4.000 ;
    END
  END Xio[2]
  PIN Xio[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.910 0.000 146.190 4.000 ;
    END
  END Xio[3]
  PIN Xro[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.150 0.000 120.430 4.000 ;
    END
  END Xro[0]
  PIN Xro[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.510 0.000 127.790 4.000 ;
    END
  END Xro[1]
  PIN Xro[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.870 0.000 135.150 4.000 ;
    END
  END Xro[2]
  PIN Xro[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.230 0.000 142.510 4.000 ;
    END
  END Xro[3]
  PIN c1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.000 23.840 182.000 24.440 ;
    END
  END c1
  PIN c2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.000 72.120 182.000 72.720 ;
    END
  END c2
  PIN c3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.000 120.400 182.000 121.000 ;
    END
  END c3
  PIN la_oenb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.590 0.000 149.870 4.000 ;
    END
  END la_oenb[0]
  PIN la_oenb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.270 0.000 153.550 4.000 ;
    END
  END la_oenb[1]
  PIN la_oenb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.950 0.000 157.230 4.000 ;
    END
  END la_oenb[2]
  PIN la_oenb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.630 0.000 160.910 4.000 ;
    END
  END la_oenb[3]
  PIN la_oenb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 0.000 164.590 4.000 ;
    END
  END la_oenb[4]
  PIN la_oenb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.990 0.000 168.270 4.000 ;
    END
  END la_oenb[5]
  PIN la_oenb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.670 0.000 171.950 4.000 ;
    END
  END la_oenb[6]
  PIN la_oenb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.350 0.000 175.630 4.000 ;
    END
  END la_oenb[7]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 182.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 182.480 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 182.480 ;
    END
  END vssd1
  PIN xi0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.070 0.000 6.350 4.000 ;
    END
  END xi0[0]
  PIN xi0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 4.000 ;
    END
  END xi0[1]
  PIN xi0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.950 0.000 65.230 4.000 ;
    END
  END xi0[2]
  PIN xi0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.390 0.000 94.670 4.000 ;
    END
  END xi0[3]
  PIN xi1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.430 0.000 13.710 4.000 ;
    END
  END xi1[0]
  PIN xi1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.870 0.000 43.150 4.000 ;
    END
  END xi1[1]
  PIN xi1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.310 0.000 72.590 4.000 ;
    END
  END xi1[2]
  PIN xi1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.750 0.000 102.030 4.000 ;
    END
  END xi1[3]
  PIN xi2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 0.000 21.070 4.000 ;
    END
  END xi2[0]
  PIN xi2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.230 0.000 50.510 4.000 ;
    END
  END xi2[1]
  PIN xi2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.670 0.000 79.950 4.000 ;
    END
  END xi2[2]
  PIN xi2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.110 0.000 109.390 4.000 ;
    END
  END xi2[3]
  PIN xi3[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.150 0.000 28.430 4.000 ;
    END
  END xi3[0]
  PIN xi3[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.590 0.000 57.870 4.000 ;
    END
  END xi3[1]
  PIN xi3[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 4.000 ;
    END
  END xi3[2]
  PIN xi3[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.470 0.000 116.750 4.000 ;
    END
  END xi3[3]
  PIN xr0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.390 0.000 2.670 4.000 ;
    END
  END xr0[0]
  PIN xr0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.830 0.000 32.110 4.000 ;
    END
  END xr0[1]
  PIN xr0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 4.000 ;
    END
  END xr0[2]
  PIN xr0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.710 0.000 90.990 4.000 ;
    END
  END xr0[3]
  PIN xr1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 0.000 10.030 4.000 ;
    END
  END xr1[0]
  PIN xr1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.190 0.000 39.470 4.000 ;
    END
  END xr1[1]
  PIN xr1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.630 0.000 68.910 4.000 ;
    END
  END xr1[2]
  PIN xr1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.070 0.000 98.350 4.000 ;
    END
  END xr1[3]
  PIN xr2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.110 0.000 17.390 4.000 ;
    END
  END xr2[0]
  PIN xr2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.550 0.000 46.830 4.000 ;
    END
  END xr2[1]
  PIN xr2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.990 0.000 76.270 4.000 ;
    END
  END xr2[2]
  PIN xr2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.430 0.000 105.710 4.000 ;
    END
  END xr2[3]
  PIN xr3[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.470 0.000 24.750 4.000 ;
    END
  END xr3[0]
  PIN xr3[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.910 0.000 54.190 4.000 ;
    END
  END xr3[1]
  PIN xr3[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.350 0.000 83.630 4.000 ;
    END
  END xr3[2]
  PIN xr3[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 0.000 113.070 4.000 ;
    END
  END xr3[3]
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 176.180 182.325 ;
      LAYER met1 ;
        RECT 2.370 4.460 179.330 182.480 ;
      LAYER met2 ;
        RECT 2.400 4.280 179.300 182.425 ;
        RECT 2.950 3.670 5.790 4.280 ;
        RECT 6.630 3.670 9.470 4.280 ;
        RECT 10.310 3.670 13.150 4.280 ;
        RECT 13.990 3.670 16.830 4.280 ;
        RECT 17.670 3.670 20.510 4.280 ;
        RECT 21.350 3.670 24.190 4.280 ;
        RECT 25.030 3.670 27.870 4.280 ;
        RECT 28.710 3.670 31.550 4.280 ;
        RECT 32.390 3.670 35.230 4.280 ;
        RECT 36.070 3.670 38.910 4.280 ;
        RECT 39.750 3.670 42.590 4.280 ;
        RECT 43.430 3.670 46.270 4.280 ;
        RECT 47.110 3.670 49.950 4.280 ;
        RECT 50.790 3.670 53.630 4.280 ;
        RECT 54.470 3.670 57.310 4.280 ;
        RECT 58.150 3.670 60.990 4.280 ;
        RECT 61.830 3.670 64.670 4.280 ;
        RECT 65.510 3.670 68.350 4.280 ;
        RECT 69.190 3.670 72.030 4.280 ;
        RECT 72.870 3.670 75.710 4.280 ;
        RECT 76.550 3.670 79.390 4.280 ;
        RECT 80.230 3.670 83.070 4.280 ;
        RECT 83.910 3.670 86.750 4.280 ;
        RECT 87.590 3.670 90.430 4.280 ;
        RECT 91.270 3.670 94.110 4.280 ;
        RECT 94.950 3.670 97.790 4.280 ;
        RECT 98.630 3.670 101.470 4.280 ;
        RECT 102.310 3.670 105.150 4.280 ;
        RECT 105.990 3.670 108.830 4.280 ;
        RECT 109.670 3.670 112.510 4.280 ;
        RECT 113.350 3.670 116.190 4.280 ;
        RECT 117.030 3.670 119.870 4.280 ;
        RECT 120.710 3.670 123.550 4.280 ;
        RECT 124.390 3.670 127.230 4.280 ;
        RECT 128.070 3.670 130.910 4.280 ;
        RECT 131.750 3.670 134.590 4.280 ;
        RECT 135.430 3.670 138.270 4.280 ;
        RECT 139.110 3.670 141.950 4.280 ;
        RECT 142.790 3.670 145.630 4.280 ;
        RECT 146.470 3.670 149.310 4.280 ;
        RECT 150.150 3.670 152.990 4.280 ;
        RECT 153.830 3.670 156.670 4.280 ;
        RECT 157.510 3.670 160.350 4.280 ;
        RECT 161.190 3.670 164.030 4.280 ;
        RECT 164.870 3.670 167.710 4.280 ;
        RECT 168.550 3.670 171.390 4.280 ;
        RECT 172.230 3.670 175.070 4.280 ;
        RECT 175.910 3.670 178.750 4.280 ;
      LAYER met3 ;
        RECT 21.050 169.680 178.000 182.405 ;
        RECT 21.050 168.280 177.600 169.680 ;
        RECT 21.050 121.400 178.000 168.280 ;
        RECT 21.050 120.000 177.600 121.400 ;
        RECT 21.050 73.120 178.000 120.000 ;
        RECT 21.050 71.720 177.600 73.120 ;
        RECT 21.050 24.840 178.000 71.720 ;
        RECT 21.050 23.440 177.600 24.840 ;
        RECT 21.050 10.715 178.000 23.440 ;
  END
END R4_butter
END LIBRARY

