magic
tech sky130A
magscale 1 2
timestamp 1676037725
<< locali >>
rect 0 1397 3114 1431
rect 430 724 464 1167
rect 430 690 559 724
rect 1741 690 1775 724
rect 345 485 379 551
rect 212 361 246 427
rect 79 237 113 303
rect 0 -17 3114 17
use sky130_sram_1kbyte_1rw1r_32x256_8_pdriver_3  sky130_sram_1kbyte_1rw1r_32x256_8_pdriver_3_0
timestamp 1676037725
transform 1 0 478 0 1 0
box -36 -17 2672 1471
use sky130_sram_1kbyte_1rw1r_32x256_8_pnand3  sky130_sram_1kbyte_1rw1r_32x256_8_pnand3_0
timestamp 1676037725
transform 1 0 0 0 1 0
box -36 -17 514 1471
<< labels >>
rlabel locali s 1758 707 1758 707 4 Z
rlabel locali s 96 270 96 270 4 A
rlabel locali s 229 394 229 394 4 B
rlabel locali s 362 518 362 518 4 C
rlabel locali s 1557 0 1557 0 4 gnd
rlabel locali s 1557 1414 1557 1414 4 vdd
<< properties >>
string FIXED_BBOX 0 0 3114 1414
string GDS_END 6270182
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_1kbyte_1rw1r_32x256_8.gds
string GDS_START 6268934
<< end >>
