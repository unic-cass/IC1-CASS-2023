magic
tech sky130B
magscale 1 2
timestamp 1676037725
<< dnwell >>
rect -40 86 86 3350
rect 4306 86 4432 3350
rect -40 -40 4432 86
<< nwell >>
rect -120 166 166 3350
rect 4226 166 4512 3350
rect -120 -120 4512 166
<< mvnsubdiff >>
rect 6 3316 40 3350
rect 6 3248 40 3282
rect 6 3180 40 3214
rect 6 3112 40 3146
rect 6 3044 40 3078
rect 6 2976 40 3010
rect 6 2908 40 2942
rect 6 2840 40 2874
rect 6 2772 40 2806
rect 6 2704 40 2738
rect 6 2636 40 2670
rect 6 2568 40 2602
rect 6 2500 40 2534
rect 6 2432 40 2466
rect 6 2364 40 2398
rect 6 2296 40 2330
rect 6 2228 40 2262
rect 6 2160 40 2194
rect 6 2092 40 2126
rect 6 2024 40 2058
rect 6 1956 40 1990
rect 6 1888 40 1922
rect 6 1820 40 1854
rect 6 1752 40 1786
rect 6 1684 40 1718
rect 6 1616 40 1650
rect 6 1548 40 1582
rect 6 1480 40 1514
rect 6 1412 40 1446
rect 6 1344 40 1378
rect 6 1276 40 1310
rect 6 1208 40 1242
rect 6 1140 40 1174
rect 6 1072 40 1106
rect 6 1004 40 1038
rect 6 936 40 970
rect 6 868 40 902
rect 6 800 40 834
rect 6 732 40 766
rect 6 664 40 698
rect 6 596 40 630
rect 6 528 40 562
rect 6 460 40 494
rect 6 392 40 426
rect 6 324 40 358
rect 6 256 40 290
rect 6 188 40 222
rect 6 120 40 154
rect 6 40 40 86
rect 4352 3304 4386 3350
rect 4352 3236 4386 3270
rect 4352 3168 4386 3202
rect 4352 3100 4386 3134
rect 4352 3032 4386 3066
rect 4352 2964 4386 2998
rect 4352 2896 4386 2930
rect 4352 2828 4386 2862
rect 4352 2760 4386 2794
rect 4352 2692 4386 2726
rect 4352 2624 4386 2658
rect 4352 2556 4386 2590
rect 4352 2488 4386 2522
rect 4352 2420 4386 2454
rect 4352 2352 4386 2386
rect 4352 2284 4386 2318
rect 4352 2216 4386 2250
rect 4352 2148 4386 2182
rect 4352 2080 4386 2114
rect 4352 2012 4386 2046
rect 4352 1944 4386 1978
rect 4352 1876 4386 1910
rect 4352 1808 4386 1842
rect 4352 1740 4386 1774
rect 4352 1672 4386 1706
rect 4352 1604 4386 1638
rect 4352 1536 4386 1570
rect 4352 1468 4386 1502
rect 4352 1400 4386 1434
rect 4352 1332 4386 1366
rect 4352 1264 4386 1298
rect 4352 1196 4386 1230
rect 4352 1128 4386 1162
rect 4352 1060 4386 1094
rect 4352 992 4386 1026
rect 4352 924 4386 958
rect 4352 856 4386 890
rect 4352 788 4386 822
rect 4352 720 4386 754
rect 4352 652 4386 686
rect 4352 584 4386 618
rect 4352 516 4386 550
rect 4352 448 4386 482
rect 4352 380 4386 414
rect 4352 312 4386 346
rect 4352 244 4386 278
rect 4352 176 4386 210
rect 4352 108 4386 142
rect 4352 40 4386 74
rect 6 6 74 40
rect 108 6 142 40
rect 176 6 210 40
rect 244 6 278 40
rect 312 6 346 40
rect 380 6 414 40
rect 448 6 482 40
rect 516 6 550 40
rect 584 6 618 40
rect 652 6 686 40
rect 720 6 754 40
rect 788 6 822 40
rect 856 6 890 40
rect 924 6 958 40
rect 992 6 1026 40
rect 1060 6 1094 40
rect 1128 6 1162 40
rect 1196 6 1230 40
rect 1264 6 1298 40
rect 1332 6 1366 40
rect 1400 6 1434 40
rect 1468 6 1502 40
rect 1536 6 1570 40
rect 1604 6 1638 40
rect 1672 6 1706 40
rect 1740 6 1774 40
rect 1808 6 1842 40
rect 1876 6 1910 40
rect 1944 6 1978 40
rect 2012 6 2046 40
rect 2080 6 2114 40
rect 2148 6 2182 40
rect 2216 6 2250 40
rect 2284 6 2318 40
rect 2352 6 2386 40
rect 2420 6 2454 40
rect 2488 6 2522 40
rect 2556 6 2590 40
rect 2624 6 2658 40
rect 2692 6 2726 40
rect 2760 6 2794 40
rect 2828 6 2862 40
rect 2896 6 2930 40
rect 2964 6 2998 40
rect 3032 6 3066 40
rect 3100 6 3134 40
rect 3168 6 3202 40
rect 3236 6 3270 40
rect 3304 6 3338 40
rect 3372 6 3406 40
rect 3440 6 3474 40
rect 3508 6 3542 40
rect 3576 6 3610 40
rect 3644 6 3678 40
rect 3712 6 3746 40
rect 3780 6 3814 40
rect 3848 6 3882 40
rect 3916 6 3950 40
rect 3984 6 4018 40
rect 4052 6 4086 40
rect 4120 6 4154 40
rect 4188 6 4222 40
rect 4256 6 4386 40
<< mvnsubdiffcont >>
rect 6 3282 40 3316
rect 6 3214 40 3248
rect 6 3146 40 3180
rect 6 3078 40 3112
rect 6 3010 40 3044
rect 6 2942 40 2976
rect 6 2874 40 2908
rect 6 2806 40 2840
rect 6 2738 40 2772
rect 6 2670 40 2704
rect 6 2602 40 2636
rect 6 2534 40 2568
rect 6 2466 40 2500
rect 6 2398 40 2432
rect 6 2330 40 2364
rect 6 2262 40 2296
rect 6 2194 40 2228
rect 6 2126 40 2160
rect 6 2058 40 2092
rect 6 1990 40 2024
rect 6 1922 40 1956
rect 6 1854 40 1888
rect 6 1786 40 1820
rect 6 1718 40 1752
rect 6 1650 40 1684
rect 6 1582 40 1616
rect 6 1514 40 1548
rect 6 1446 40 1480
rect 6 1378 40 1412
rect 6 1310 40 1344
rect 6 1242 40 1276
rect 6 1174 40 1208
rect 6 1106 40 1140
rect 6 1038 40 1072
rect 6 970 40 1004
rect 6 902 40 936
rect 6 834 40 868
rect 6 766 40 800
rect 6 698 40 732
rect 6 630 40 664
rect 6 562 40 596
rect 6 494 40 528
rect 6 426 40 460
rect 6 358 40 392
rect 6 290 40 324
rect 6 222 40 256
rect 6 154 40 188
rect 6 86 40 120
rect 4352 3270 4386 3304
rect 4352 3202 4386 3236
rect 4352 3134 4386 3168
rect 4352 3066 4386 3100
rect 4352 2998 4386 3032
rect 4352 2930 4386 2964
rect 4352 2862 4386 2896
rect 4352 2794 4386 2828
rect 4352 2726 4386 2760
rect 4352 2658 4386 2692
rect 4352 2590 4386 2624
rect 4352 2522 4386 2556
rect 4352 2454 4386 2488
rect 4352 2386 4386 2420
rect 4352 2318 4386 2352
rect 4352 2250 4386 2284
rect 4352 2182 4386 2216
rect 4352 2114 4386 2148
rect 4352 2046 4386 2080
rect 4352 1978 4386 2012
rect 4352 1910 4386 1944
rect 4352 1842 4386 1876
rect 4352 1774 4386 1808
rect 4352 1706 4386 1740
rect 4352 1638 4386 1672
rect 4352 1570 4386 1604
rect 4352 1502 4386 1536
rect 4352 1434 4386 1468
rect 4352 1366 4386 1400
rect 4352 1298 4386 1332
rect 4352 1230 4386 1264
rect 4352 1162 4386 1196
rect 4352 1094 4386 1128
rect 4352 1026 4386 1060
rect 4352 958 4386 992
rect 4352 890 4386 924
rect 4352 822 4386 856
rect 4352 754 4386 788
rect 4352 686 4386 720
rect 4352 618 4386 652
rect 4352 550 4386 584
rect 4352 482 4386 516
rect 4352 414 4386 448
rect 4352 346 4386 380
rect 4352 278 4386 312
rect 4352 210 4386 244
rect 4352 142 4386 176
rect 4352 74 4386 108
rect 74 6 108 40
rect 142 6 176 40
rect 210 6 244 40
rect 278 6 312 40
rect 346 6 380 40
rect 414 6 448 40
rect 482 6 516 40
rect 550 6 584 40
rect 618 6 652 40
rect 686 6 720 40
rect 754 6 788 40
rect 822 6 856 40
rect 890 6 924 40
rect 958 6 992 40
rect 1026 6 1060 40
rect 1094 6 1128 40
rect 1162 6 1196 40
rect 1230 6 1264 40
rect 1298 6 1332 40
rect 1366 6 1400 40
rect 1434 6 1468 40
rect 1502 6 1536 40
rect 1570 6 1604 40
rect 1638 6 1672 40
rect 1706 6 1740 40
rect 1774 6 1808 40
rect 1842 6 1876 40
rect 1910 6 1944 40
rect 1978 6 2012 40
rect 2046 6 2080 40
rect 2114 6 2148 40
rect 2182 6 2216 40
rect 2250 6 2284 40
rect 2318 6 2352 40
rect 2386 6 2420 40
rect 2454 6 2488 40
rect 2522 6 2556 40
rect 2590 6 2624 40
rect 2658 6 2692 40
rect 2726 6 2760 40
rect 2794 6 2828 40
rect 2862 6 2896 40
rect 2930 6 2964 40
rect 2998 6 3032 40
rect 3066 6 3100 40
rect 3134 6 3168 40
rect 3202 6 3236 40
rect 3270 6 3304 40
rect 3338 6 3372 40
rect 3406 6 3440 40
rect 3474 6 3508 40
rect 3542 6 3576 40
rect 3610 6 3644 40
rect 3678 6 3712 40
rect 3746 6 3780 40
rect 3814 6 3848 40
rect 3882 6 3916 40
rect 3950 6 3984 40
rect 4018 6 4052 40
rect 4086 6 4120 40
rect 4154 6 4188 40
rect 4222 6 4256 40
<< locali >>
rect 6 3342 40 3350
rect 4352 3342 4386 3350
rect 0 3316 46 3342
rect 0 3276 6 3316
rect 40 3276 46 3316
rect 0 3248 46 3276
rect 0 3203 6 3248
rect 40 3203 46 3248
rect 0 3180 46 3203
rect 0 3130 6 3180
rect 40 3130 46 3180
rect 0 3112 46 3130
rect 0 3057 6 3112
rect 40 3057 46 3112
rect 0 3044 46 3057
rect 0 2984 6 3044
rect 40 2984 46 3044
rect 0 2976 46 2984
rect 0 2911 6 2976
rect 40 2911 46 2976
rect 0 2908 46 2911
rect 0 2874 6 2908
rect 40 2874 46 2908
rect 0 2872 46 2874
rect 0 2806 6 2872
rect 40 2806 46 2872
rect 0 2799 46 2806
rect 0 2738 6 2799
rect 40 2738 46 2799
rect 0 2726 46 2738
rect 0 2670 6 2726
rect 40 2670 46 2726
rect 0 2653 46 2670
rect 0 2602 6 2653
rect 40 2602 46 2653
rect 0 2580 46 2602
rect 0 2534 6 2580
rect 40 2534 46 2580
rect 0 2507 46 2534
rect 0 2466 6 2507
rect 40 2466 46 2507
rect 0 2434 46 2466
rect 0 2398 6 2434
rect 40 2398 46 2434
rect 0 2364 46 2398
rect 0 2327 6 2364
rect 40 2327 46 2364
rect 0 2296 46 2327
rect 0 2254 6 2296
rect 40 2254 46 2296
rect 0 2228 46 2254
rect 0 2181 6 2228
rect 40 2181 46 2228
rect 0 2160 46 2181
rect 0 2108 6 2160
rect 40 2108 46 2160
rect 0 2092 46 2108
rect 0 2035 6 2092
rect 40 2035 46 2092
rect 0 2024 46 2035
rect 0 1962 6 2024
rect 40 1962 46 2024
rect 0 1956 46 1962
rect 0 1889 6 1956
rect 40 1889 46 1956
rect 0 1888 46 1889
rect 0 1854 6 1888
rect 40 1854 46 1888
rect 0 1850 46 1854
rect 0 1786 6 1850
rect 40 1786 46 1850
rect 0 1777 46 1786
rect 0 1718 6 1777
rect 40 1718 46 1777
rect 0 1704 46 1718
rect 0 1650 6 1704
rect 40 1650 46 1704
rect 0 1631 46 1650
rect 0 1582 6 1631
rect 40 1582 46 1631
rect 0 1558 46 1582
rect 0 1514 6 1558
rect 40 1514 46 1558
rect 0 1485 46 1514
rect 0 1446 6 1485
rect 40 1446 46 1485
rect 0 1412 46 1446
rect 0 1378 6 1412
rect 40 1378 46 1412
rect 0 1344 46 1378
rect 0 1305 6 1344
rect 40 1305 46 1344
rect 0 1276 46 1305
rect 0 1232 6 1276
rect 40 1232 46 1276
rect 0 1208 46 1232
rect 0 1159 6 1208
rect 40 1159 46 1208
rect 0 1140 46 1159
rect 0 1086 6 1140
rect 40 1086 46 1140
rect 0 1072 46 1086
rect 0 1014 6 1072
rect 40 1014 46 1072
rect 0 1004 46 1014
rect 0 942 6 1004
rect 40 942 46 1004
rect 0 936 46 942
rect 0 870 6 936
rect 40 870 46 936
rect 0 868 46 870
rect 0 834 6 868
rect 40 834 46 868
rect 0 832 46 834
rect 0 766 6 832
rect 40 766 46 832
rect 0 760 46 766
rect 0 698 6 760
rect 40 698 46 760
rect 0 688 46 698
rect 0 630 6 688
rect 40 630 46 688
rect 0 616 46 630
rect 0 562 6 616
rect 40 562 46 616
rect 0 544 46 562
rect 0 494 6 544
rect 40 494 46 544
rect 0 472 46 494
rect 0 426 6 472
rect 40 426 46 472
rect 0 400 46 426
rect 0 358 6 400
rect 40 358 46 400
rect 0 328 46 358
rect 0 290 6 328
rect 40 290 46 328
rect 0 256 46 290
rect 0 222 6 256
rect 40 222 46 256
rect 0 188 46 222
rect 0 150 6 188
rect 40 150 46 188
rect 0 120 46 150
rect 0 78 6 120
rect 40 78 46 120
rect 0 46 46 78
rect 4352 3310 4416 3342
rect 4352 3304 4376 3310
rect 4410 3276 4416 3310
rect 4386 3270 4416 3276
rect 4352 3238 4416 3270
rect 4352 3236 4376 3238
rect 4410 3204 4416 3238
rect 4386 3202 4416 3204
rect 4352 3168 4416 3202
rect 4386 3166 4416 3168
rect 4352 3132 4376 3134
rect 4410 3132 4416 3166
rect 4352 3100 4416 3132
rect 4386 3094 4416 3100
rect 4352 3060 4376 3066
rect 4410 3060 4416 3094
rect 4352 3032 4416 3060
rect 4386 3022 4416 3032
rect 4352 2988 4376 2998
rect 4410 2988 4416 3022
rect 4352 2964 4416 2988
rect 4386 2950 4416 2964
rect 4352 2916 4376 2930
rect 4410 2916 4416 2950
rect 4352 2896 4416 2916
rect 4386 2878 4416 2896
rect 4352 2844 4376 2862
rect 4410 2844 4416 2878
rect 4352 2828 4416 2844
rect 4386 2806 4416 2828
rect 4352 2772 4376 2794
rect 4410 2772 4416 2806
rect 4352 2760 4416 2772
rect 4386 2734 4416 2760
rect 4352 2700 4376 2726
rect 4410 2700 4416 2734
rect 4352 2692 4416 2700
rect 4386 2662 4416 2692
rect 4352 2628 4376 2658
rect 4410 2628 4416 2662
rect 4352 2624 4416 2628
rect 4386 2590 4416 2624
rect 4352 2556 4376 2590
rect 4410 2556 4416 2590
rect 4386 2522 4416 2556
rect 4352 2518 4416 2522
rect 4352 2488 4376 2518
rect 4410 2484 4416 2518
rect 4386 2454 4416 2484
rect 4352 2446 4416 2454
rect 4352 2420 4376 2446
rect 4410 2412 4416 2446
rect 4386 2386 4416 2412
rect 4352 2374 4416 2386
rect 4352 2352 4376 2374
rect 4410 2340 4416 2374
rect 4386 2318 4416 2340
rect 4352 2302 4416 2318
rect 4352 2284 4376 2302
rect 4410 2268 4416 2302
rect 4386 2250 4416 2268
rect 4352 2229 4416 2250
rect 4352 2216 4376 2229
rect 4410 2195 4416 2229
rect 4386 2182 4416 2195
rect 4352 2156 4416 2182
rect 4352 2148 4376 2156
rect 4410 2122 4416 2156
rect 4386 2114 4416 2122
rect 4352 2083 4416 2114
rect 4352 2080 4376 2083
rect 4410 2049 4416 2083
rect 4386 2046 4416 2049
rect 4352 2012 4416 2046
rect 4386 2010 4416 2012
rect 4352 1976 4376 1978
rect 4410 1976 4416 2010
rect 4352 1944 4416 1976
rect 4386 1937 4416 1944
rect 4352 1903 4376 1910
rect 4410 1903 4416 1937
rect 4352 1876 4416 1903
rect 4386 1864 4416 1876
rect 4352 1830 4376 1842
rect 4410 1830 4416 1864
rect 4352 1808 4416 1830
rect 4386 1791 4416 1808
rect 4352 1757 4376 1774
rect 4410 1757 4416 1791
rect 4352 1740 4416 1757
rect 4386 1718 4416 1740
rect 4352 1684 4376 1706
rect 4410 1684 4416 1718
rect 4352 1672 4416 1684
rect 4386 1645 4416 1672
rect 4352 1611 4376 1638
rect 4410 1611 4416 1645
rect 4352 1604 4416 1611
rect 4386 1572 4416 1604
rect 4352 1538 4376 1570
rect 4410 1538 4416 1572
rect 4352 1536 4416 1538
rect 4386 1502 4416 1536
rect 4352 1499 4416 1502
rect 4352 1468 4376 1499
rect 4410 1465 4416 1499
rect 4386 1434 4416 1465
rect 4352 1426 4416 1434
rect 4352 1400 4376 1426
rect 4410 1392 4416 1426
rect 4386 1366 4416 1392
rect 4352 1353 4416 1366
rect 4352 1332 4376 1353
rect 4410 1319 4416 1353
rect 4386 1298 4416 1319
rect 4352 1280 4416 1298
rect 4352 1264 4376 1280
rect 4410 1246 4416 1280
rect 4386 1230 4416 1246
rect 4352 1207 4416 1230
rect 4352 1196 4376 1207
rect 4410 1173 4416 1207
rect 4386 1162 4416 1173
rect 4352 1134 4416 1162
rect 4352 1128 4376 1134
rect 4410 1100 4416 1134
rect 4386 1094 4416 1100
rect 4352 1061 4416 1094
rect 4352 1060 4376 1061
rect 4410 1027 4416 1061
rect 4386 1026 4416 1027
rect 4352 992 4416 1026
rect 4386 988 4416 992
rect 4352 954 4376 958
rect 4410 954 4416 988
rect 4352 924 4416 954
rect 4386 915 4416 924
rect 4352 881 4376 890
rect 4410 881 4416 915
rect 4352 856 4416 881
rect 4386 842 4416 856
rect 4352 808 4376 822
rect 4410 808 4416 842
rect 4352 788 4416 808
rect 4386 769 4416 788
rect 4352 735 4376 754
rect 4410 735 4416 769
rect 4352 720 4416 735
rect 4386 696 4416 720
rect 4352 662 4376 686
rect 4410 662 4416 696
rect 4352 652 4416 662
rect 4386 623 4416 652
rect 4352 589 4376 618
rect 4410 589 4416 623
rect 4352 584 4416 589
rect 4386 550 4416 584
rect 4352 516 4376 550
rect 4410 516 4416 550
rect 4386 482 4416 516
rect 4352 477 4416 482
rect 4352 448 4376 477
rect 4410 443 4416 477
rect 4386 414 4416 443
rect 4352 404 4416 414
rect 4352 380 4376 404
rect 4410 370 4416 404
rect 4386 346 4416 370
rect 4352 331 4416 346
rect 4352 312 4376 331
rect 4410 297 4416 331
rect 4386 278 4416 297
rect 4352 258 4416 278
rect 4352 244 4376 258
rect 4410 224 4416 258
rect 4386 210 4416 224
rect 4352 185 4416 210
rect 4352 176 4376 185
rect 4410 151 4416 185
rect 4386 142 4416 151
rect 4352 112 4416 142
rect 4352 108 4376 112
rect 4410 78 4416 112
rect 4386 74 4416 78
rect 4352 46 4416 74
rect 0 40 4416 46
rect 0 6 74 40
rect 112 6 142 40
rect 185 6 210 40
rect 258 6 278 40
rect 331 6 346 40
rect 404 6 414 40
rect 477 6 482 40
rect 584 6 589 40
rect 652 6 662 40
rect 720 6 734 40
rect 788 6 806 40
rect 856 6 878 40
rect 924 6 950 40
rect 992 6 1022 40
rect 1060 6 1094 40
rect 1128 6 1162 40
rect 1200 6 1230 40
rect 1272 6 1298 40
rect 1344 6 1366 40
rect 1400 6 1408 40
rect 1468 6 1481 40
rect 1536 6 1554 40
rect 1604 6 1627 40
rect 1672 6 1700 40
rect 1740 6 1773 40
rect 1808 6 1842 40
rect 1880 6 1910 40
rect 1953 6 1978 40
rect 2026 6 2046 40
rect 2099 6 2114 40
rect 2172 6 2182 40
rect 2245 6 2250 40
rect 2352 6 2357 40
rect 2420 6 2430 40
rect 2488 6 2503 40
rect 2556 6 2576 40
rect 2624 6 2648 40
rect 2692 6 2720 40
rect 2760 6 2792 40
rect 2828 6 2862 40
rect 2898 6 2930 40
rect 2970 6 2998 40
rect 3042 6 3066 40
rect 3114 6 3134 40
rect 3186 6 3202 40
rect 3258 6 3270 40
rect 3330 6 3338 40
rect 3402 6 3406 40
rect 3508 6 3512 40
rect 3576 6 3584 40
rect 3644 6 3656 40
rect 3712 6 3728 40
rect 3780 6 3800 40
rect 3848 6 3872 40
rect 3916 6 3944 40
rect 3984 6 4016 40
rect 4052 6 4086 40
rect 4122 6 4154 40
rect 4194 6 4222 40
rect 4266 6 4304 40
rect 4338 6 4416 40
rect 0 0 4416 6
<< viali >>
rect 6 3282 40 3310
rect 6 3276 40 3282
rect 6 3214 40 3237
rect 6 3203 40 3214
rect 6 3146 40 3164
rect 6 3130 40 3146
rect 6 3078 40 3091
rect 6 3057 40 3078
rect 6 3010 40 3018
rect 6 2984 40 3010
rect 6 2942 40 2945
rect 6 2911 40 2942
rect 6 2840 40 2872
rect 6 2838 40 2840
rect 6 2772 40 2799
rect 6 2765 40 2772
rect 6 2704 40 2726
rect 6 2692 40 2704
rect 6 2636 40 2653
rect 6 2619 40 2636
rect 6 2568 40 2580
rect 6 2546 40 2568
rect 6 2500 40 2507
rect 6 2473 40 2500
rect 6 2432 40 2434
rect 6 2400 40 2432
rect 6 2330 40 2361
rect 6 2327 40 2330
rect 6 2262 40 2288
rect 6 2254 40 2262
rect 6 2194 40 2215
rect 6 2181 40 2194
rect 6 2126 40 2142
rect 6 2108 40 2126
rect 6 2058 40 2069
rect 6 2035 40 2058
rect 6 1990 40 1996
rect 6 1962 40 1990
rect 6 1922 40 1923
rect 6 1889 40 1922
rect 6 1820 40 1850
rect 6 1816 40 1820
rect 6 1752 40 1777
rect 6 1743 40 1752
rect 6 1684 40 1704
rect 6 1670 40 1684
rect 6 1616 40 1631
rect 6 1597 40 1616
rect 6 1548 40 1558
rect 6 1524 40 1548
rect 6 1480 40 1485
rect 6 1451 40 1480
rect 6 1378 40 1412
rect 6 1310 40 1339
rect 6 1305 40 1310
rect 6 1242 40 1266
rect 6 1232 40 1242
rect 6 1174 40 1193
rect 6 1159 40 1174
rect 6 1106 40 1120
rect 6 1086 40 1106
rect 6 1038 40 1048
rect 6 1014 40 1038
rect 6 970 40 976
rect 6 942 40 970
rect 6 902 40 904
rect 6 870 40 902
rect 6 800 40 832
rect 6 798 40 800
rect 6 732 40 760
rect 6 726 40 732
rect 6 664 40 688
rect 6 654 40 664
rect 6 596 40 616
rect 6 582 40 596
rect 6 528 40 544
rect 6 510 40 528
rect 6 460 40 472
rect 6 438 40 460
rect 6 392 40 400
rect 6 366 40 392
rect 6 324 40 328
rect 6 294 40 324
rect 6 222 40 256
rect 6 154 40 184
rect 6 150 40 154
rect 6 86 40 112
rect 6 78 40 86
rect 4376 3304 4410 3310
rect 4376 3276 4386 3304
rect 4386 3276 4410 3304
rect 4376 3236 4410 3238
rect 4376 3204 4386 3236
rect 4386 3204 4410 3236
rect 4376 3134 4386 3166
rect 4386 3134 4410 3166
rect 4376 3132 4410 3134
rect 4376 3066 4386 3094
rect 4386 3066 4410 3094
rect 4376 3060 4410 3066
rect 4376 2998 4386 3022
rect 4386 2998 4410 3022
rect 4376 2988 4410 2998
rect 4376 2930 4386 2950
rect 4386 2930 4410 2950
rect 4376 2916 4410 2930
rect 4376 2862 4386 2878
rect 4386 2862 4410 2878
rect 4376 2844 4410 2862
rect 4376 2794 4386 2806
rect 4386 2794 4410 2806
rect 4376 2772 4410 2794
rect 4376 2726 4386 2734
rect 4386 2726 4410 2734
rect 4376 2700 4410 2726
rect 4376 2658 4386 2662
rect 4386 2658 4410 2662
rect 4376 2628 4410 2658
rect 4376 2556 4410 2590
rect 4376 2488 4410 2518
rect 4376 2484 4386 2488
rect 4386 2484 4410 2488
rect 4376 2420 4410 2446
rect 4376 2412 4386 2420
rect 4386 2412 4410 2420
rect 4376 2352 4410 2374
rect 4376 2340 4386 2352
rect 4386 2340 4410 2352
rect 4376 2284 4410 2302
rect 4376 2268 4386 2284
rect 4386 2268 4410 2284
rect 4376 2216 4410 2229
rect 4376 2195 4386 2216
rect 4386 2195 4410 2216
rect 4376 2148 4410 2156
rect 4376 2122 4386 2148
rect 4386 2122 4410 2148
rect 4376 2080 4410 2083
rect 4376 2049 4386 2080
rect 4386 2049 4410 2080
rect 4376 1978 4386 2010
rect 4386 1978 4410 2010
rect 4376 1976 4410 1978
rect 4376 1910 4386 1937
rect 4386 1910 4410 1937
rect 4376 1903 4410 1910
rect 4376 1842 4386 1864
rect 4386 1842 4410 1864
rect 4376 1830 4410 1842
rect 4376 1774 4386 1791
rect 4386 1774 4410 1791
rect 4376 1757 4410 1774
rect 4376 1706 4386 1718
rect 4386 1706 4410 1718
rect 4376 1684 4410 1706
rect 4376 1638 4386 1645
rect 4386 1638 4410 1645
rect 4376 1611 4410 1638
rect 4376 1570 4386 1572
rect 4386 1570 4410 1572
rect 4376 1538 4410 1570
rect 4376 1468 4410 1499
rect 4376 1465 4386 1468
rect 4386 1465 4410 1468
rect 4376 1400 4410 1426
rect 4376 1392 4386 1400
rect 4386 1392 4410 1400
rect 4376 1332 4410 1353
rect 4376 1319 4386 1332
rect 4386 1319 4410 1332
rect 4376 1264 4410 1280
rect 4376 1246 4386 1264
rect 4386 1246 4410 1264
rect 4376 1196 4410 1207
rect 4376 1173 4386 1196
rect 4386 1173 4410 1196
rect 4376 1128 4410 1134
rect 4376 1100 4386 1128
rect 4386 1100 4410 1128
rect 4376 1060 4410 1061
rect 4376 1027 4386 1060
rect 4386 1027 4410 1060
rect 4376 958 4386 988
rect 4386 958 4410 988
rect 4376 954 4410 958
rect 4376 890 4386 915
rect 4386 890 4410 915
rect 4376 881 4410 890
rect 4376 822 4386 842
rect 4386 822 4410 842
rect 4376 808 4410 822
rect 4376 754 4386 769
rect 4386 754 4410 769
rect 4376 735 4410 754
rect 4376 686 4386 696
rect 4386 686 4410 696
rect 4376 662 4410 686
rect 4376 618 4386 623
rect 4386 618 4410 623
rect 4376 589 4410 618
rect 4376 516 4410 550
rect 4376 448 4410 477
rect 4376 443 4386 448
rect 4386 443 4410 448
rect 4376 380 4410 404
rect 4376 370 4386 380
rect 4386 370 4410 380
rect 4376 312 4410 331
rect 4376 297 4386 312
rect 4386 297 4410 312
rect 4376 244 4410 258
rect 4376 224 4386 244
rect 4386 224 4410 244
rect 4376 176 4410 185
rect 4376 151 4386 176
rect 4386 151 4410 176
rect 4376 108 4410 112
rect 4376 78 4386 108
rect 4386 78 4410 108
rect 78 6 108 40
rect 108 6 112 40
rect 151 6 176 40
rect 176 6 185 40
rect 224 6 244 40
rect 244 6 258 40
rect 297 6 312 40
rect 312 6 331 40
rect 370 6 380 40
rect 380 6 404 40
rect 443 6 448 40
rect 448 6 477 40
rect 516 6 550 40
rect 589 6 618 40
rect 618 6 623 40
rect 662 6 686 40
rect 686 6 696 40
rect 734 6 754 40
rect 754 6 768 40
rect 806 6 822 40
rect 822 6 840 40
rect 878 6 890 40
rect 890 6 912 40
rect 950 6 958 40
rect 958 6 984 40
rect 1022 6 1026 40
rect 1026 6 1056 40
rect 1094 6 1128 40
rect 1166 6 1196 40
rect 1196 6 1200 40
rect 1238 6 1264 40
rect 1264 6 1272 40
rect 1310 6 1332 40
rect 1332 6 1344 40
rect 1408 6 1434 40
rect 1434 6 1442 40
rect 1481 6 1502 40
rect 1502 6 1515 40
rect 1554 6 1570 40
rect 1570 6 1588 40
rect 1627 6 1638 40
rect 1638 6 1661 40
rect 1700 6 1706 40
rect 1706 6 1734 40
rect 1773 6 1774 40
rect 1774 6 1807 40
rect 1846 6 1876 40
rect 1876 6 1880 40
rect 1919 6 1944 40
rect 1944 6 1953 40
rect 1992 6 2012 40
rect 2012 6 2026 40
rect 2065 6 2080 40
rect 2080 6 2099 40
rect 2138 6 2148 40
rect 2148 6 2172 40
rect 2211 6 2216 40
rect 2216 6 2245 40
rect 2284 6 2318 40
rect 2357 6 2386 40
rect 2386 6 2391 40
rect 2430 6 2454 40
rect 2454 6 2464 40
rect 2503 6 2522 40
rect 2522 6 2537 40
rect 2576 6 2590 40
rect 2590 6 2610 40
rect 2648 6 2658 40
rect 2658 6 2682 40
rect 2720 6 2726 40
rect 2726 6 2754 40
rect 2792 6 2794 40
rect 2794 6 2826 40
rect 2864 6 2896 40
rect 2896 6 2898 40
rect 2936 6 2964 40
rect 2964 6 2970 40
rect 3008 6 3032 40
rect 3032 6 3042 40
rect 3080 6 3100 40
rect 3100 6 3114 40
rect 3152 6 3168 40
rect 3168 6 3186 40
rect 3224 6 3236 40
rect 3236 6 3258 40
rect 3296 6 3304 40
rect 3304 6 3330 40
rect 3368 6 3372 40
rect 3372 6 3402 40
rect 3440 6 3474 40
rect 3512 6 3542 40
rect 3542 6 3546 40
rect 3584 6 3610 40
rect 3610 6 3618 40
rect 3656 6 3678 40
rect 3678 6 3690 40
rect 3728 6 3746 40
rect 3746 6 3762 40
rect 3800 6 3814 40
rect 3814 6 3834 40
rect 3872 6 3882 40
rect 3882 6 3906 40
rect 3944 6 3950 40
rect 3950 6 3978 40
rect 4016 6 4018 40
rect 4018 6 4050 40
rect 4088 6 4120 40
rect 4120 6 4122 40
rect 4160 6 4188 40
rect 4188 6 4194 40
rect 4232 6 4256 40
rect 4256 6 4266 40
rect 4304 6 4338 40
<< metal1 >>
rect 0 3310 46 3342
rect 0 3276 6 3310
rect 40 3276 46 3310
rect 0 3237 46 3276
rect 0 3203 6 3237
rect 40 3203 46 3237
rect 0 3164 46 3203
rect 0 3130 6 3164
rect 40 3130 46 3164
rect 0 3091 46 3130
rect 0 3057 6 3091
rect 40 3057 46 3091
rect 0 3018 46 3057
rect 0 2984 6 3018
rect 40 2984 46 3018
rect 0 2945 46 2984
rect 0 2911 6 2945
rect 40 2911 46 2945
rect 0 2872 46 2911
rect 0 2838 6 2872
rect 40 2838 46 2872
rect 0 2799 46 2838
rect 0 2765 6 2799
rect 40 2765 46 2799
rect 0 2726 46 2765
rect 0 2692 6 2726
rect 40 2692 46 2726
rect 0 2653 46 2692
rect 0 2619 6 2653
rect 40 2619 46 2653
rect 0 2580 46 2619
rect 0 2546 6 2580
rect 40 2546 46 2580
rect 0 2507 46 2546
rect 0 2473 6 2507
rect 40 2473 46 2507
rect 0 2434 46 2473
rect 0 2400 6 2434
rect 40 2400 46 2434
rect 0 2361 46 2400
rect 0 2327 6 2361
rect 40 2327 46 2361
rect 0 2288 46 2327
rect 0 2254 6 2288
rect 40 2254 46 2288
rect 0 2215 46 2254
rect 0 2181 6 2215
rect 40 2181 46 2215
rect 0 2142 46 2181
rect 0 2108 6 2142
rect 40 2108 46 2142
rect 0 2069 46 2108
rect 0 2035 6 2069
rect 40 2035 46 2069
rect 0 1996 46 2035
rect 0 1962 6 1996
rect 40 1962 46 1996
rect 0 1923 46 1962
rect 0 1889 6 1923
rect 40 1889 46 1923
rect 0 1850 46 1889
rect 0 1816 6 1850
rect 40 1816 46 1850
rect 0 1777 46 1816
rect 0 1743 6 1777
rect 40 1743 46 1777
rect 0 1704 46 1743
rect 0 1670 6 1704
rect 40 1670 46 1704
rect 0 1631 46 1670
rect 0 1597 6 1631
rect 40 1597 46 1631
rect 0 1558 46 1597
rect 0 1524 6 1558
rect 40 1524 46 1558
rect 0 1485 46 1524
rect 0 1451 6 1485
rect 40 1451 46 1485
rect 0 1412 46 1451
rect 0 1378 6 1412
rect 40 1378 46 1412
rect 0 1339 46 1378
rect 0 1305 6 1339
rect 40 1305 46 1339
rect 0 1266 46 1305
rect 0 1232 6 1266
rect 40 1232 46 1266
rect 0 1193 46 1232
rect 0 1159 6 1193
rect 40 1159 46 1193
rect 0 1120 46 1159
rect 0 1086 6 1120
rect 40 1086 46 1120
rect 0 1048 46 1086
rect 0 1014 6 1048
rect 40 1014 46 1048
rect 0 976 46 1014
rect 0 942 6 976
rect 40 942 46 976
rect 0 904 46 942
rect 0 870 6 904
rect 40 870 46 904
rect 0 832 46 870
rect 0 798 6 832
rect 40 798 46 832
rect 0 760 46 798
rect 0 726 6 760
rect 40 726 46 760
rect 0 688 46 726
rect 0 654 6 688
rect 40 654 46 688
rect 0 616 46 654
rect 0 582 6 616
rect 40 582 46 616
rect 0 544 46 582
rect 0 510 6 544
rect 40 510 46 544
rect 0 472 46 510
rect 0 438 6 472
rect 40 438 46 472
rect 0 400 46 438
rect 0 366 6 400
rect 40 366 46 400
rect 0 328 46 366
rect 0 294 6 328
rect 40 294 46 328
rect 0 256 46 294
rect 0 222 6 256
rect 40 222 46 256
rect 0 184 46 222
rect 0 150 6 184
rect 40 150 46 184
rect 0 112 46 150
rect 0 78 6 112
rect 40 78 46 112
rect 0 46 46 78
rect 4370 3310 4416 3342
rect 4370 3276 4376 3310
rect 4410 3276 4416 3310
rect 4370 3238 4416 3276
rect 4370 3204 4376 3238
rect 4410 3204 4416 3238
rect 4370 3166 4416 3204
rect 4370 3132 4376 3166
rect 4410 3132 4416 3166
rect 4370 3094 4416 3132
rect 4370 3060 4376 3094
rect 4410 3060 4416 3094
rect 4370 3022 4416 3060
rect 4370 2988 4376 3022
rect 4410 2988 4416 3022
rect 4370 2950 4416 2988
rect 4370 2916 4376 2950
rect 4410 2916 4416 2950
rect 4370 2878 4416 2916
rect 4370 2844 4376 2878
rect 4410 2844 4416 2878
rect 4370 2806 4416 2844
rect 4370 2772 4376 2806
rect 4410 2772 4416 2806
rect 4370 2734 4416 2772
rect 4370 2700 4376 2734
rect 4410 2700 4416 2734
rect 4370 2662 4416 2700
rect 4370 2628 4376 2662
rect 4410 2628 4416 2662
rect 4370 2590 4416 2628
rect 4370 2556 4376 2590
rect 4410 2556 4416 2590
rect 4370 2518 4416 2556
rect 4370 2484 4376 2518
rect 4410 2484 4416 2518
rect 4370 2446 4416 2484
rect 4370 2412 4376 2446
rect 4410 2412 4416 2446
rect 4370 2374 4416 2412
rect 4370 2340 4376 2374
rect 4410 2340 4416 2374
rect 4370 2302 4416 2340
rect 4370 2268 4376 2302
rect 4410 2268 4416 2302
rect 4370 2229 4416 2268
rect 4370 2195 4376 2229
rect 4410 2195 4416 2229
rect 4370 2156 4416 2195
rect 4370 2122 4376 2156
rect 4410 2122 4416 2156
rect 4370 2083 4416 2122
rect 4370 2049 4376 2083
rect 4410 2049 4416 2083
rect 4370 2010 4416 2049
rect 4370 1976 4376 2010
rect 4410 1976 4416 2010
rect 4370 1937 4416 1976
rect 4370 1903 4376 1937
rect 4410 1903 4416 1937
rect 4370 1864 4416 1903
rect 4370 1830 4376 1864
rect 4410 1830 4416 1864
rect 4370 1791 4416 1830
rect 4370 1757 4376 1791
rect 4410 1757 4416 1791
rect 4370 1718 4416 1757
rect 4370 1684 4376 1718
rect 4410 1684 4416 1718
rect 4370 1645 4416 1684
rect 4370 1611 4376 1645
rect 4410 1611 4416 1645
rect 4370 1572 4416 1611
rect 4370 1538 4376 1572
rect 4410 1538 4416 1572
rect 4370 1499 4416 1538
rect 4370 1465 4376 1499
rect 4410 1465 4416 1499
rect 4370 1426 4416 1465
rect 4370 1392 4376 1426
rect 4410 1392 4416 1426
rect 4370 1353 4416 1392
rect 4370 1319 4376 1353
rect 4410 1319 4416 1353
rect 4370 1280 4416 1319
rect 4370 1246 4376 1280
rect 4410 1246 4416 1280
rect 4370 1207 4416 1246
rect 4370 1173 4376 1207
rect 4410 1173 4416 1207
rect 4370 1134 4416 1173
rect 4370 1100 4376 1134
rect 4410 1100 4416 1134
rect 4370 1061 4416 1100
rect 4370 1027 4376 1061
rect 4410 1027 4416 1061
rect 4370 988 4416 1027
rect 4370 954 4376 988
rect 4410 954 4416 988
rect 4370 915 4416 954
rect 4370 881 4376 915
rect 4410 881 4416 915
rect 4370 842 4416 881
rect 4370 808 4376 842
rect 4410 808 4416 842
rect 4370 769 4416 808
rect 4370 735 4376 769
rect 4410 735 4416 769
rect 4370 696 4416 735
rect 4370 662 4376 696
rect 4410 662 4416 696
rect 4370 623 4416 662
rect 4370 589 4376 623
rect 4410 589 4416 623
rect 4370 550 4416 589
rect 4370 516 4376 550
rect 4410 516 4416 550
rect 4370 477 4416 516
rect 4370 443 4376 477
rect 4410 443 4416 477
rect 4370 404 4416 443
rect 4370 370 4376 404
rect 4410 370 4416 404
rect 4370 331 4416 370
rect 4370 297 4376 331
rect 4410 297 4416 331
rect 4370 258 4416 297
rect 4370 224 4376 258
rect 4410 224 4416 258
rect 4370 185 4416 224
rect 4370 151 4376 185
rect 4410 151 4416 185
rect 4370 112 4416 151
rect 4370 78 4376 112
rect 4410 78 4416 112
rect 4370 46 4416 78
rect 0 40 4416 46
rect 0 6 78 40
rect 112 6 151 40
rect 185 6 224 40
rect 258 6 297 40
rect 331 6 370 40
rect 404 6 443 40
rect 477 6 516 40
rect 550 6 589 40
rect 623 6 662 40
rect 696 6 734 40
rect 768 6 806 40
rect 840 6 878 40
rect 912 6 950 40
rect 984 6 1022 40
rect 1056 6 1094 40
rect 1128 6 1166 40
rect 1200 6 1238 40
rect 1272 6 1310 40
rect 1344 6 1408 40
rect 1442 6 1481 40
rect 1515 6 1554 40
rect 1588 6 1627 40
rect 1661 6 1700 40
rect 1734 6 1773 40
rect 1807 6 1846 40
rect 1880 6 1919 40
rect 1953 6 1992 40
rect 2026 6 2065 40
rect 2099 6 2138 40
rect 2172 6 2211 40
rect 2245 6 2284 40
rect 2318 6 2357 40
rect 2391 6 2430 40
rect 2464 6 2503 40
rect 2537 6 2576 40
rect 2610 6 2648 40
rect 2682 6 2720 40
rect 2754 6 2792 40
rect 2826 6 2864 40
rect 2898 6 2936 40
rect 2970 6 3008 40
rect 3042 6 3080 40
rect 3114 6 3152 40
rect 3186 6 3224 40
rect 3258 6 3296 40
rect 3330 6 3368 40
rect 3402 6 3440 40
rect 3474 6 3512 40
rect 3546 6 3584 40
rect 3618 6 3656 40
rect 3690 6 3728 40
rect 3762 6 3800 40
rect 3834 6 3872 40
rect 3906 6 3944 40
rect 3978 6 4016 40
rect 4050 6 4088 40
rect 4122 6 4160 40
rect 4194 6 4232 40
rect 4266 6 4304 40
rect 4338 6 4416 40
rect 0 0 4416 6
<< properties >>
string GDS_END 29704758
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 29684210
<< end >>
