magic
tech sky130A
magscale 1 2
timestamp 1676037725
<< locali >>
rect 238 961 588 980
rect 116 823 182 889
rect 238 855 252 961
rect 574 855 588 961
rect 238 841 588 855
rect 644 823 710 889
rect 116 795 160 823
rect 666 795 710 823
rect 41 759 160 795
rect 41 725 60 759
rect 94 725 160 759
rect 41 687 160 725
rect 41 653 60 687
rect 94 653 160 687
rect 41 615 160 653
rect 41 581 60 615
rect 94 581 160 615
rect 41 543 160 581
rect 41 509 60 543
rect 94 509 160 543
rect 41 471 160 509
rect 41 437 60 471
rect 94 437 160 471
rect 41 399 160 437
rect 41 365 60 399
rect 94 365 160 399
rect 41 327 160 365
rect 41 293 60 327
rect 94 293 160 327
rect 41 255 160 293
rect 41 221 60 255
rect 94 221 160 255
rect 41 185 160 221
rect 666 759 785 795
rect 666 725 732 759
rect 766 725 785 759
rect 666 687 785 725
rect 666 653 732 687
rect 766 653 785 687
rect 666 615 785 653
rect 666 581 732 615
rect 766 581 785 615
rect 666 543 785 581
rect 666 509 732 543
rect 766 509 785 543
rect 666 471 785 509
rect 666 437 732 471
rect 766 437 785 471
rect 666 399 785 437
rect 666 365 732 399
rect 766 365 785 399
rect 666 327 785 365
rect 666 293 732 327
rect 766 293 785 327
rect 666 255 785 293
rect 666 221 732 255
rect 766 221 785 255
rect 666 185 785 221
rect 116 157 160 185
rect 666 157 710 185
rect 116 91 182 157
rect 238 125 588 139
rect 238 19 252 125
rect 574 19 588 125
rect 644 91 710 157
rect 238 0 588 19
<< viali >>
rect 252 855 574 961
rect 60 725 94 759
rect 60 653 94 687
rect 60 581 94 615
rect 60 509 94 543
rect 60 437 94 471
rect 60 365 94 399
rect 60 293 94 327
rect 60 221 94 255
rect 732 725 766 759
rect 732 653 766 687
rect 732 581 766 615
rect 732 509 766 543
rect 732 437 766 471
rect 732 365 766 399
rect 732 293 766 327
rect 732 221 766 255
rect 252 19 574 125
<< obsli1 >>
rect 212 185 246 795
rect 304 185 338 795
rect 396 185 430 795
rect 488 185 522 795
rect 580 185 614 795
<< metal1 >>
rect 236 961 590 980
rect 236 855 252 961
rect 574 855 590 961
rect 236 843 590 855
rect 41 759 100 771
rect 41 725 60 759
rect 94 725 100 759
rect 41 687 100 725
rect 41 653 60 687
rect 94 653 100 687
rect 41 615 100 653
rect 41 581 60 615
rect 94 581 100 615
rect 41 543 100 581
rect 41 509 60 543
rect 94 509 100 543
rect 41 471 100 509
rect 41 437 60 471
rect 94 437 100 471
rect 41 399 100 437
rect 41 365 60 399
rect 94 365 100 399
rect 41 327 100 365
rect 41 293 60 327
rect 94 293 100 327
rect 41 255 100 293
rect 41 221 60 255
rect 94 221 100 255
rect 41 209 100 221
rect 726 759 785 771
rect 726 725 732 759
rect 766 725 785 759
rect 726 687 785 725
rect 726 653 732 687
rect 766 653 785 687
rect 726 615 785 653
rect 726 581 732 615
rect 766 581 785 615
rect 726 543 785 581
rect 726 509 732 543
rect 766 509 785 543
rect 726 471 785 509
rect 726 437 732 471
rect 766 437 785 471
rect 726 399 785 437
rect 726 365 732 399
rect 766 365 785 399
rect 726 327 785 365
rect 726 293 732 327
rect 766 293 785 327
rect 726 255 785 293
rect 726 221 732 255
rect 766 221 785 255
rect 726 209 785 221
rect 236 125 590 137
rect 236 19 252 125
rect 574 19 590 125
rect 236 0 590 19
<< obsm1 >>
rect 203 209 255 771
rect 295 209 347 771
rect 387 209 439 771
rect 479 209 531 771
rect 571 209 623 771
<< metal2 >>
rect 14 515 812 771
rect 14 209 812 465
<< labels >>
rlabel viali s 732 725 766 759 6 BULK
port 4 nsew
rlabel viali s 732 653 766 687 6 BULK
port 4 nsew
rlabel viali s 732 581 766 615 6 BULK
port 4 nsew
rlabel viali s 732 509 766 543 6 BULK
port 4 nsew
rlabel viali s 732 437 766 471 6 BULK
port 4 nsew
rlabel viali s 732 365 766 399 6 BULK
port 4 nsew
rlabel viali s 732 293 766 327 6 BULK
port 4 nsew
rlabel viali s 732 221 766 255 6 BULK
port 4 nsew
rlabel viali s 60 725 94 759 6 BULK
port 4 nsew
rlabel viali s 60 653 94 687 6 BULK
port 4 nsew
rlabel viali s 60 581 94 615 6 BULK
port 4 nsew
rlabel viali s 60 509 94 543 6 BULK
port 4 nsew
rlabel viali s 60 437 94 471 6 BULK
port 4 nsew
rlabel viali s 60 365 94 399 6 BULK
port 4 nsew
rlabel viali s 60 293 94 327 6 BULK
port 4 nsew
rlabel viali s 60 221 94 255 6 BULK
port 4 nsew
rlabel locali s 666 795 710 823 6 BULK
port 4 nsew
rlabel locali s 666 185 785 795 6 BULK
port 4 nsew
rlabel locali s 666 157 710 185 6 BULK
port 4 nsew
rlabel locali s 644 823 710 889 6 BULK
port 4 nsew
rlabel locali s 644 91 710 157 6 BULK
port 4 nsew
rlabel locali s 116 823 182 889 6 BULK
port 4 nsew
rlabel locali s 116 795 160 823 6 BULK
port 4 nsew
rlabel locali s 116 157 160 185 6 BULK
port 4 nsew
rlabel locali s 116 91 182 157 6 BULK
port 4 nsew
rlabel locali s 41 185 160 795 6 BULK
port 4 nsew
rlabel metal1 s 726 209 785 771 6 BULK
port 4 nsew
rlabel metal1 s 41 209 100 771 6 BULK
port 4 nsew
rlabel metal2 s 14 515 812 771 6 DRAIN
port 1 nsew
rlabel viali s 252 855 574 961 6 GATE
port 2 nsew
rlabel viali s 252 19 574 125 6 GATE
port 2 nsew
rlabel locali s 238 841 588 980 6 GATE
port 2 nsew
rlabel locali s 238 0 588 139 6 GATE
port 2 nsew
rlabel metal1 s 236 843 590 980 6 GATE
port 2 nsew
rlabel metal1 s 236 0 590 137 6 GATE
port 2 nsew
rlabel metal2 s 14 209 812 465 6 SOURCE
port 3 nsew
<< properties >>
string FIXED_BBOX 0 0 826 980
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 9697378
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 9676500
string device primitive
<< end >>