VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO R4_butter
  CLASS BLOCK ;
  FOREIGN R4_butter ;
  ORIGIN 0.000 0.000 ;
  SIZE 182.000 BY 194.000 ;
  PIN Xio[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.000 49.000 182.000 49.600 ;
    END
  END Xio[0]
  PIN Xio[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.000 96.600 182.000 97.200 ;
    END
  END Xio[1]
  PIN Xio[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.000 144.200 182.000 144.800 ;
    END
  END Xio[2]
  PIN Xio[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.000 187.040 182.000 187.640 ;
    END
  END Xio[3]
  PIN Xro[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.000 44.240 182.000 44.840 ;
    END
  END Xro[0]
  PIN Xro[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.000 91.840 182.000 92.440 ;
    END
  END Xro[1]
  PIN Xro[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.000 139.440 182.000 140.040 ;
    END
  END Xro[2]
  PIN Xro[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.000 182.280 182.000 182.880 ;
    END
  END Xro[3]
  PIN c1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 190.000 22.910 194.000 ;
    END
  END c1
  PIN c2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.170 190.000 68.450 194.000 ;
    END
  END c2
  PIN c3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.710 190.000 113.990 194.000 ;
    END
  END c3
  PIN la_oenb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.050 0.000 12.330 4.000 ;
    END
  END la_oenb[0]
  PIN la_oenb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.590 0.000 34.870 4.000 ;
    END
  END la_oenb[1]
  PIN la_oenb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.130 0.000 57.410 4.000 ;
    END
  END la_oenb[2]
  PIN la_oenb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.670 0.000 79.950 4.000 ;
    END
  END la_oenb[3]
  PIN la_oenb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.210 0.000 102.490 4.000 ;
    END
  END la_oenb[4]
  PIN la_oenb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.750 0.000 125.030 4.000 ;
    END
  END la_oenb[5]
  PIN la_oenb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.290 0.000 147.570 4.000 ;
    END
  END la_oenb[6]
  PIN la_oenb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.830 0.000 170.110 4.000 ;
    END
  END la_oenb[7]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 182.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 182.480 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 182.480 ;
    END
  END vssd1
  PIN xi0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.000 10.920 182.000 11.520 ;
    END
  END xi0[0]
  PIN xi0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.000 58.520 182.000 59.120 ;
    END
  END xi0[1]
  PIN xi0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.000 106.120 182.000 106.720 ;
    END
  END xi0[2]
  PIN xi0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.000 153.720 182.000 154.320 ;
    END
  END xi0[3]
  PIN xi1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.000 20.440 182.000 21.040 ;
    END
  END xi1[0]
  PIN xi1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.000 68.040 182.000 68.640 ;
    END
  END xi1[1]
  PIN xi1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.000 115.640 182.000 116.240 ;
    END
  END xi1[2]
  PIN xi1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.000 163.240 182.000 163.840 ;
    END
  END xi1[3]
  PIN xi2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.000 29.960 182.000 30.560 ;
    END
  END xi2[0]
  PIN xi2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.000 77.560 182.000 78.160 ;
    END
  END xi2[1]
  PIN xi2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.000 125.160 182.000 125.760 ;
    END
  END xi2[2]
  PIN xi2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.000 172.760 182.000 173.360 ;
    END
  END xi2[3]
  PIN xi3[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.000 39.480 182.000 40.080 ;
    END
  END xi3[0]
  PIN xi3[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.000 87.080 182.000 87.680 ;
    END
  END xi3[1]
  PIN xi3[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.000 134.680 182.000 135.280 ;
    END
  END xi3[2]
  PIN xi3[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.250 190.000 159.530 194.000 ;
    END
  END xi3[3]
  PIN xr0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.000 6.160 182.000 6.760 ;
    END
  END xr0[0]
  PIN xr0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.000 53.760 182.000 54.360 ;
    END
  END xr0[1]
  PIN xr0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.000 101.360 182.000 101.960 ;
    END
  END xr0[2]
  PIN xr0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.000 148.960 182.000 149.560 ;
    END
  END xr0[3]
  PIN xr1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.000 15.680 182.000 16.280 ;
    END
  END xr1[0]
  PIN xr1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.000 63.280 182.000 63.880 ;
    END
  END xr1[1]
  PIN xr1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.000 110.880 182.000 111.480 ;
    END
  END xr1[2]
  PIN xr1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.000 158.480 182.000 159.080 ;
    END
  END xr1[3]
  PIN xr2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.000 25.200 182.000 25.800 ;
    END
  END xr2[0]
  PIN xr2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.000 72.800 182.000 73.400 ;
    END
  END xr2[1]
  PIN xr2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.000 120.400 182.000 121.000 ;
    END
  END xr2[2]
  PIN xr2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.000 168.000 182.000 168.600 ;
    END
  END xr2[3]
  PIN xr3[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.000 34.720 182.000 35.320 ;
    END
  END xr3[0]
  PIN xr3[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.000 82.320 182.000 82.920 ;
    END
  END xr3[1]
  PIN xr3[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.000 129.920 182.000 130.520 ;
    END
  END xr3[2]
  PIN xr3[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.000 177.520 182.000 178.120 ;
    END
  END xr3[3]
  OBS
      LAYER nwell ;
        RECT 5.330 180.825 176.370 182.430 ;
        RECT 5.330 175.385 176.370 178.215 ;
        RECT 5.330 169.945 176.370 172.775 ;
        RECT 5.330 164.505 176.370 167.335 ;
        RECT 5.330 159.065 176.370 161.895 ;
        RECT 5.330 153.625 176.370 156.455 ;
        RECT 5.330 148.185 176.370 151.015 ;
        RECT 5.330 142.745 176.370 145.575 ;
        RECT 5.330 137.305 176.370 140.135 ;
        RECT 5.330 131.865 176.370 134.695 ;
        RECT 5.330 126.425 176.370 129.255 ;
        RECT 5.330 120.985 176.370 123.815 ;
        RECT 5.330 115.545 176.370 118.375 ;
        RECT 5.330 110.105 176.370 112.935 ;
        RECT 5.330 104.665 176.370 107.495 ;
        RECT 5.330 99.225 176.370 102.055 ;
        RECT 5.330 93.785 176.370 96.615 ;
        RECT 5.330 88.345 176.370 91.175 ;
        RECT 5.330 82.905 176.370 85.735 ;
        RECT 5.330 77.465 176.370 80.295 ;
        RECT 5.330 72.025 176.370 74.855 ;
        RECT 5.330 66.585 176.370 69.415 ;
        RECT 5.330 61.145 176.370 63.975 ;
        RECT 5.330 55.705 176.370 58.535 ;
        RECT 5.330 50.265 176.370 53.095 ;
        RECT 5.330 44.825 176.370 47.655 ;
        RECT 5.330 39.385 176.370 42.215 ;
        RECT 5.330 33.945 176.370 36.775 ;
        RECT 5.330 28.505 176.370 31.335 ;
        RECT 5.330 23.065 176.370 25.895 ;
        RECT 5.330 17.625 176.370 20.455 ;
        RECT 5.330 12.185 176.370 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 176.180 182.325 ;
      LAYER met1 ;
        RECT 5.520 10.640 179.330 182.480 ;
      LAYER met2 ;
        RECT 12.060 189.720 22.350 190.810 ;
        RECT 23.190 189.720 67.890 190.810 ;
        RECT 68.730 189.720 113.430 190.810 ;
        RECT 114.270 189.720 158.970 190.810 ;
        RECT 159.810 189.720 179.300 190.810 ;
        RECT 12.060 4.280 179.300 189.720 ;
        RECT 12.610 4.000 34.310 4.280 ;
        RECT 35.150 4.000 56.850 4.280 ;
        RECT 57.690 4.000 79.390 4.280 ;
        RECT 80.230 4.000 101.930 4.280 ;
        RECT 102.770 4.000 124.470 4.280 ;
        RECT 125.310 4.000 147.010 4.280 ;
        RECT 147.850 4.000 169.550 4.280 ;
        RECT 170.390 4.000 179.300 4.280 ;
      LAYER met3 ;
        RECT 21.050 186.640 177.600 187.505 ;
        RECT 21.050 183.280 178.000 186.640 ;
        RECT 21.050 181.880 177.600 183.280 ;
        RECT 21.050 178.520 178.000 181.880 ;
        RECT 21.050 177.120 177.600 178.520 ;
        RECT 21.050 173.760 178.000 177.120 ;
        RECT 21.050 172.360 177.600 173.760 ;
        RECT 21.050 169.000 178.000 172.360 ;
        RECT 21.050 167.600 177.600 169.000 ;
        RECT 21.050 164.240 178.000 167.600 ;
        RECT 21.050 162.840 177.600 164.240 ;
        RECT 21.050 159.480 178.000 162.840 ;
        RECT 21.050 158.080 177.600 159.480 ;
        RECT 21.050 154.720 178.000 158.080 ;
        RECT 21.050 153.320 177.600 154.720 ;
        RECT 21.050 149.960 178.000 153.320 ;
        RECT 21.050 148.560 177.600 149.960 ;
        RECT 21.050 145.200 178.000 148.560 ;
        RECT 21.050 143.800 177.600 145.200 ;
        RECT 21.050 140.440 178.000 143.800 ;
        RECT 21.050 139.040 177.600 140.440 ;
        RECT 21.050 135.680 178.000 139.040 ;
        RECT 21.050 134.280 177.600 135.680 ;
        RECT 21.050 130.920 178.000 134.280 ;
        RECT 21.050 129.520 177.600 130.920 ;
        RECT 21.050 126.160 178.000 129.520 ;
        RECT 21.050 124.760 177.600 126.160 ;
        RECT 21.050 121.400 178.000 124.760 ;
        RECT 21.050 120.000 177.600 121.400 ;
        RECT 21.050 116.640 178.000 120.000 ;
        RECT 21.050 115.240 177.600 116.640 ;
        RECT 21.050 111.880 178.000 115.240 ;
        RECT 21.050 110.480 177.600 111.880 ;
        RECT 21.050 107.120 178.000 110.480 ;
        RECT 21.050 105.720 177.600 107.120 ;
        RECT 21.050 102.360 178.000 105.720 ;
        RECT 21.050 100.960 177.600 102.360 ;
        RECT 21.050 97.600 178.000 100.960 ;
        RECT 21.050 96.200 177.600 97.600 ;
        RECT 21.050 92.840 178.000 96.200 ;
        RECT 21.050 91.440 177.600 92.840 ;
        RECT 21.050 88.080 178.000 91.440 ;
        RECT 21.050 86.680 177.600 88.080 ;
        RECT 21.050 83.320 178.000 86.680 ;
        RECT 21.050 81.920 177.600 83.320 ;
        RECT 21.050 78.560 178.000 81.920 ;
        RECT 21.050 77.160 177.600 78.560 ;
        RECT 21.050 73.800 178.000 77.160 ;
        RECT 21.050 72.400 177.600 73.800 ;
        RECT 21.050 69.040 178.000 72.400 ;
        RECT 21.050 67.640 177.600 69.040 ;
        RECT 21.050 64.280 178.000 67.640 ;
        RECT 21.050 62.880 177.600 64.280 ;
        RECT 21.050 59.520 178.000 62.880 ;
        RECT 21.050 58.120 177.600 59.520 ;
        RECT 21.050 54.760 178.000 58.120 ;
        RECT 21.050 53.360 177.600 54.760 ;
        RECT 21.050 50.000 178.000 53.360 ;
        RECT 21.050 48.600 177.600 50.000 ;
        RECT 21.050 45.240 178.000 48.600 ;
        RECT 21.050 43.840 177.600 45.240 ;
        RECT 21.050 40.480 178.000 43.840 ;
        RECT 21.050 39.080 177.600 40.480 ;
        RECT 21.050 35.720 178.000 39.080 ;
        RECT 21.050 34.320 177.600 35.720 ;
        RECT 21.050 30.960 178.000 34.320 ;
        RECT 21.050 29.560 177.600 30.960 ;
        RECT 21.050 26.200 178.000 29.560 ;
        RECT 21.050 24.800 177.600 26.200 ;
        RECT 21.050 21.440 178.000 24.800 ;
        RECT 21.050 20.040 177.600 21.440 ;
        RECT 21.050 16.680 178.000 20.040 ;
        RECT 21.050 15.280 177.600 16.680 ;
        RECT 21.050 11.920 178.000 15.280 ;
        RECT 21.050 10.520 177.600 11.920 ;
        RECT 21.050 7.160 178.000 10.520 ;
        RECT 21.050 6.295 177.600 7.160 ;
  END
END R4_butter
END LIBRARY

