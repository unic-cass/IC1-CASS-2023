magic
tech sky130A
magscale 1 2
timestamp 1676037725
<< nwell >>
rect -66 377 2082 897
<< pwell >>
rect 1736 281 1994 283
rect 1412 269 1994 281
rect 4 242 418 269
rect 848 242 1994 269
rect 4 43 1994 242
rect -26 -43 2042 43
<< locali >>
rect 122 277 188 440
rect 672 293 738 395
rect 1647 625 1720 689
rect 1670 405 1720 625
rect 1670 345 1736 405
rect 1926 379 1999 747
rect 1945 243 1999 379
rect 1926 103 1999 243
<< obsli1 >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2016 831
rect 22 754 666 763
rect 22 729 172 754
rect 22 695 28 729
rect 62 695 100 729
rect 134 720 172 729
rect 206 720 244 754
rect 278 720 316 754
rect 350 720 399 754
rect 433 720 471 754
rect 505 729 666 754
rect 505 720 543 729
rect 134 711 543 720
rect 134 695 205 711
rect 22 689 205 695
rect 533 695 543 711
rect 577 695 615 729
rect 649 695 666 729
rect 1137 757 1892 763
rect 1137 743 1639 757
rect 1137 729 1287 743
rect 533 689 666 695
rect 22 440 88 689
rect 239 633 499 677
rect 334 377 400 599
rect 455 463 499 633
rect 600 497 666 689
rect 704 677 1103 711
rect 1137 695 1143 729
rect 1177 695 1215 729
rect 1249 709 1287 729
rect 1321 709 1359 743
rect 1393 729 1639 743
rect 1393 709 1431 729
rect 1249 695 1431 709
rect 1465 695 1503 729
rect 1537 723 1639 729
rect 1673 723 1711 757
rect 1745 729 1892 757
rect 1745 723 1783 729
rect 1537 695 1613 723
rect 1137 689 1613 695
rect 1754 695 1783 723
rect 1817 695 1855 729
rect 1889 695 1892 729
rect 1754 689 1892 695
rect 704 463 738 677
rect 455 429 738 463
rect 772 601 1035 643
rect 319 311 421 377
rect 28 125 94 234
rect 334 168 400 311
rect 455 216 494 429
rect 444 141 494 216
rect 528 259 594 393
rect 772 259 814 601
rect 528 225 814 259
rect 28 119 153 125
rect 28 85 35 119
rect 69 85 107 119
rect 141 85 153 119
rect 28 73 153 85
rect 231 107 373 134
rect 528 107 562 225
rect 231 73 562 107
rect 596 125 666 191
rect 764 141 814 225
rect 875 466 932 532
rect 1069 519 1103 677
rect 1027 485 1103 519
rect 875 273 909 466
rect 1027 389 1061 485
rect 1164 466 1230 689
rect 1332 417 1386 532
rect 1430 445 1496 689
rect 943 323 1061 389
rect 1103 375 1386 417
rect 1103 307 1169 375
rect 1332 365 1386 375
rect 1491 365 1557 411
rect 1225 273 1298 331
rect 875 239 1298 273
rect 596 119 730 125
rect 596 85 599 119
rect 633 85 671 119
rect 705 107 730 119
rect 875 107 932 239
rect 1164 125 1230 205
rect 705 105 785 107
rect 705 85 743 105
rect 596 71 743 85
rect 777 71 785 105
rect 596 51 785 71
rect 819 51 932 107
rect 966 119 1230 125
rect 966 105 1118 119
rect 966 71 974 105
rect 1008 71 1046 105
rect 1080 85 1118 105
rect 1152 85 1190 119
rect 1224 85 1230 119
rect 1080 71 1230 85
rect 1264 134 1298 239
rect 1332 323 1557 365
rect 1332 168 1386 323
rect 1491 277 1557 323
rect 1591 311 1636 591
rect 1754 439 1820 689
rect 1789 311 1911 345
rect 1591 277 1911 311
rect 1591 243 1636 277
rect 1430 177 1636 243
rect 1264 71 1382 134
rect 1754 125 1820 243
rect 1416 119 1892 125
rect 1416 105 1708 119
rect 1416 71 1420 105
rect 1454 71 1492 105
rect 1526 71 1564 105
rect 1598 71 1636 105
rect 1670 85 1708 105
rect 1742 85 1780 119
rect 1814 85 1852 119
rect 1886 85 1892 119
rect 1670 71 1892 85
rect 966 51 1230 71
rect 1416 51 1892 71
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
<< obsli1c >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 895 797 929 831
rect 991 797 1025 831
rect 1087 797 1121 831
rect 1183 797 1217 831
rect 1279 797 1313 831
rect 1375 797 1409 831
rect 1471 797 1505 831
rect 1567 797 1601 831
rect 1663 797 1697 831
rect 1759 797 1793 831
rect 1855 797 1889 831
rect 1951 797 1985 831
rect 28 695 62 729
rect 100 695 134 729
rect 172 720 206 754
rect 244 720 278 754
rect 316 720 350 754
rect 399 720 433 754
rect 471 720 505 754
rect 543 695 577 729
rect 615 695 649 729
rect 1143 695 1177 729
rect 1215 695 1249 729
rect 1287 709 1321 743
rect 1359 709 1393 743
rect 1431 695 1465 729
rect 1503 695 1537 729
rect 1639 723 1673 757
rect 1711 723 1745 757
rect 1783 695 1817 729
rect 1855 695 1889 729
rect 35 85 69 119
rect 107 85 141 119
rect 599 85 633 119
rect 671 85 705 119
rect 743 71 777 105
rect 974 71 1008 105
rect 1046 71 1080 105
rect 1118 85 1152 119
rect 1190 85 1224 119
rect 1420 71 1454 105
rect 1492 71 1526 105
rect 1564 71 1598 105
rect 1636 71 1670 105
rect 1708 85 1742 119
rect 1780 85 1814 119
rect 1852 85 1886 119
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
<< metal1 >>
rect 0 831 2016 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2016 831
rect 0 791 2016 797
rect 0 757 2016 763
rect 0 754 1639 757
rect 0 729 172 754
rect 0 695 28 729
rect 62 695 100 729
rect 134 720 172 729
rect 206 720 244 754
rect 278 720 316 754
rect 350 720 399 754
rect 433 720 471 754
rect 505 743 1639 754
rect 505 729 1287 743
rect 505 720 543 729
rect 134 695 543 720
rect 577 695 615 729
rect 649 695 1143 729
rect 1177 695 1215 729
rect 1249 709 1287 729
rect 1321 709 1359 743
rect 1393 729 1639 743
rect 1393 709 1431 729
rect 1249 695 1431 709
rect 1465 695 1503 729
rect 1537 723 1639 729
rect 1673 723 1711 757
rect 1745 729 2016 757
rect 1745 723 1783 729
rect 1537 695 1783 723
rect 1817 695 1855 729
rect 1889 695 2016 729
rect 0 689 2016 695
rect 0 119 2016 125
rect 0 85 35 119
rect 69 85 107 119
rect 141 85 599 119
rect 633 85 671 119
rect 705 105 1118 119
rect 705 85 743 105
rect 0 71 743 85
rect 777 71 974 105
rect 1008 71 1046 105
rect 1080 85 1118 105
rect 1152 85 1190 119
rect 1224 105 1708 119
rect 1224 85 1420 105
rect 1080 71 1420 85
rect 1454 71 1492 105
rect 1526 71 1564 105
rect 1598 71 1636 105
rect 1670 85 1708 105
rect 1742 85 1780 119
rect 1814 85 1852 119
rect 1886 85 2016 119
rect 1670 71 2016 85
rect 0 51 2016 71
rect 0 17 2016 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
rect 0 -23 2016 -17
<< labels >>
rlabel locali s 1670 345 1736 405 6 CLK
port 1 nsew clock input
rlabel locali s 672 293 738 395 6 CLK
port 1 nsew clock input
rlabel locali s 1670 405 1720 625 6 CLK
port 1 nsew clock input
rlabel locali s 1647 625 1720 689 6 CLK
port 1 nsew clock input
rlabel locali s 122 277 188 440 6 GATE
port 2 nsew signal input
rlabel metal1 s 0 51 2016 125 6 VGND
port 3 nsew ground bidirectional
rlabel metal1 s 0 -23 2016 23 8 VNB
port 4 nsew ground bidirectional
rlabel pwell s -26 -43 2042 43 8 VNB
port 4 nsew ground bidirectional
rlabel pwell s 4 43 1994 242 6 VNB
port 4 nsew ground bidirectional
rlabel pwell s 848 242 1994 269 6 VNB
port 4 nsew ground bidirectional
rlabel pwell s 4 242 418 269 6 VNB
port 4 nsew ground bidirectional
rlabel pwell s 1412 269 1994 281 6 VNB
port 4 nsew ground bidirectional
rlabel pwell s 1736 281 1994 283 6 VNB
port 4 nsew ground bidirectional
rlabel metal1 s 0 791 2016 837 6 VPB
port 5 nsew power bidirectional
rlabel nwell s -66 377 2082 897 6 VPB
port 5 nsew power bidirectional
rlabel metal1 s 0 689 2016 763 6 VPWR
port 6 nsew power bidirectional
rlabel locali s 1926 103 1999 243 6 GCLK
port 7 nsew signal output
rlabel locali s 1945 243 1999 379 6 GCLK
port 7 nsew signal output
rlabel locali s 1926 379 1999 747 6 GCLK
port 7 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 2016 814
string LEFclass CORE
string LEFsite unithv
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 1183864
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string GDS_START 1159928
<< end >>
