magic
tech sky130B
magscale 1 2
timestamp 1676037725
<< nwell >>
rect -38 261 774 582
<< pwell >>
rect 549 157 735 203
rect 1 21 735 157
rect 29 -17 63 21
<< scnmos >>
rect 79 47 109 131
rect 267 47 297 131
rect 339 47 369 131
rect 439 47 469 131
rect 527 47 557 131
rect 627 47 657 177
<< scpmoshvt >>
rect 79 413 109 497
rect 163 413 193 497
rect 287 413 317 497
rect 439 413 469 497
rect 532 413 562 497
rect 627 297 657 497
<< ndiff >>
rect 575 131 627 177
rect 27 101 79 131
rect 27 67 35 101
rect 69 67 79 101
rect 27 47 79 67
rect 109 93 161 131
rect 109 59 119 93
rect 153 59 161 93
rect 109 47 161 59
rect 215 101 267 131
rect 215 67 223 101
rect 257 67 267 101
rect 215 47 267 67
rect 297 47 339 131
rect 369 47 439 131
rect 469 47 527 131
rect 557 93 627 131
rect 557 59 567 93
rect 601 59 627 93
rect 557 47 627 59
rect 657 161 709 177
rect 657 127 667 161
rect 701 127 709 161
rect 657 93 709 127
rect 657 59 667 93
rect 701 59 709 93
rect 657 47 709 59
<< pdiff >>
rect 27 477 79 497
rect 27 443 35 477
rect 69 443 79 477
rect 27 413 79 443
rect 109 485 163 497
rect 109 451 119 485
rect 153 451 163 485
rect 109 413 163 451
rect 193 477 287 497
rect 193 443 230 477
rect 264 443 287 477
rect 193 413 287 443
rect 317 479 439 497
rect 317 445 327 479
rect 361 445 395 479
rect 429 445 439 479
rect 317 413 439 445
rect 469 477 532 497
rect 469 443 488 477
rect 522 443 532 477
rect 469 413 532 443
rect 562 479 627 497
rect 562 445 578 479
rect 612 445 627 479
rect 562 413 627 445
rect 577 297 627 413
rect 657 453 709 497
rect 657 419 667 453
rect 701 419 709 453
rect 657 349 709 419
rect 657 315 667 349
rect 701 315 709 349
rect 657 297 709 315
<< ndiffc >>
rect 35 67 69 101
rect 119 59 153 93
rect 223 67 257 101
rect 567 59 601 93
rect 667 127 701 161
rect 667 59 701 93
<< pdiffc >>
rect 35 443 69 477
rect 119 451 153 485
rect 230 443 264 477
rect 327 445 361 479
rect 395 445 429 479
rect 488 443 522 477
rect 578 445 612 479
rect 667 419 701 453
rect 667 315 701 349
<< poly >>
rect 79 497 109 523
rect 163 497 193 523
rect 287 497 317 523
rect 439 497 469 523
rect 532 497 562 523
rect 627 497 657 523
rect 79 265 109 413
rect 163 265 193 413
rect 287 281 317 413
rect 287 271 369 281
rect 21 249 109 265
rect 21 215 31 249
rect 65 215 109 249
rect 21 199 109 215
rect 152 249 206 265
rect 152 215 162 249
rect 196 215 206 249
rect 287 237 314 271
rect 348 237 369 271
rect 439 265 469 413
rect 532 265 562 413
rect 627 265 657 297
rect 287 227 369 237
rect 152 199 206 215
rect 79 131 109 199
rect 175 176 206 199
rect 175 146 297 176
rect 267 131 297 146
rect 339 131 369 227
rect 415 249 469 265
rect 415 215 425 249
rect 459 215 469 249
rect 415 199 469 215
rect 511 249 565 265
rect 511 215 521 249
rect 555 215 565 249
rect 511 199 565 215
rect 607 249 661 265
rect 607 215 617 249
rect 651 215 661 249
rect 607 199 661 215
rect 439 131 469 199
rect 527 131 557 199
rect 627 177 657 199
rect 79 21 109 47
rect 267 21 297 47
rect 339 21 369 47
rect 439 21 469 47
rect 527 21 557 47
rect 627 21 657 47
<< polycont >>
rect 31 215 65 249
rect 162 215 196 249
rect 314 237 348 271
rect 425 215 459 249
rect 521 215 555 249
rect 617 215 651 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 34 477 69 493
rect 34 443 35 477
rect 34 403 69 443
rect 103 485 169 527
rect 103 451 119 485
rect 153 451 169 485
rect 103 439 169 451
rect 230 477 264 493
rect 311 479 445 527
rect 311 445 327 479
rect 361 445 395 479
rect 429 445 445 479
rect 488 477 522 493
rect 230 409 264 443
rect 562 479 628 527
rect 562 445 578 479
rect 612 445 628 479
rect 667 453 719 493
rect 488 409 522 443
rect 701 419 719 453
rect 34 369 160 403
rect 17 249 90 335
rect 17 215 31 249
rect 65 215 90 249
rect 17 199 90 215
rect 126 265 160 369
rect 230 375 633 409
rect 126 249 196 265
rect 126 215 162 249
rect 126 199 196 215
rect 126 165 160 199
rect 34 131 160 165
rect 34 101 69 131
rect 230 117 264 375
rect 34 67 35 101
rect 218 101 264 117
rect 34 51 69 67
rect 103 59 119 93
rect 153 59 169 93
rect 103 17 169 59
rect 218 67 223 101
rect 257 67 264 101
rect 304 271 360 339
rect 304 237 314 271
rect 348 237 360 271
rect 304 84 360 237
rect 405 249 459 339
rect 405 215 425 249
rect 405 84 459 215
rect 497 249 565 339
rect 497 215 521 249
rect 555 215 565 249
rect 497 133 565 215
rect 599 265 633 375
rect 667 349 719 419
rect 701 315 719 349
rect 667 299 719 315
rect 599 249 651 265
rect 599 215 617 249
rect 599 199 651 215
rect 685 161 719 299
rect 651 127 667 161
rect 701 127 719 161
rect 651 93 719 127
rect 218 51 264 67
rect 551 59 567 93
rect 601 59 617 93
rect 651 59 667 93
rect 701 68 719 93
rect 701 59 718 68
rect 551 17 617 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional abutment
flabel locali s 406 289 440 323 0 FreeSans 200 0 0 0 C
port 3 nsew signal input
flabel locali s 29 289 63 323 0 FreeSans 200 0 0 0 A_N
port 1 nsew signal input
flabel locali s 673 85 707 119 0 FreeSans 200 0 0 0 X
port 9 nsew signal output
flabel locali s 673 357 707 391 0 FreeSans 200 0 0 0 X
port 9 nsew signal output
flabel locali s 673 425 707 459 0 FreeSans 200 0 0 0 X
port 9 nsew signal output
flabel locali s 29 221 63 255 0 FreeSans 200 0 0 0 A_N
port 1 nsew signal input
flabel locali s 500 221 534 255 0 FreeSans 200 0 0 0 D
port 4 nsew signal input
flabel locali s 500 289 534 323 0 FreeSans 200 0 0 0 D
port 4 nsew signal input
flabel locali s 406 85 440 119 0 FreeSans 200 0 0 0 C
port 3 nsew signal input
flabel locali s 406 153 440 187 0 FreeSans 200 0 0 0 C
port 3 nsew signal input
flabel locali s 305 85 339 119 0 FreeSans 200 0 0 0 B
port 2 nsew signal input
flabel locali s 305 153 339 187 0 FreeSans 200 0 0 0 B
port 2 nsew signal input
flabel locali s 305 221 339 255 0 FreeSans 200 0 0 0 B
port 2 nsew signal input
flabel locali s 305 289 339 323 0 FreeSans 200 0 0 0 B
port 2 nsew signal input
flabel locali s 500 153 534 187 0 FreeSans 200 0 0 0 D
port 4 nsew signal input
flabel locali s 406 221 440 255 0 FreeSans 200 0 0 0 C
port 3 nsew signal input
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
rlabel comment s 0 0 0 0 4 and4b_1
rlabel metal1 s 0 -48 736 48 1 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 496 736 592 1 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 736 544
string GDS_END 3065058
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3057504
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 18.400 0.000 
<< end >>
