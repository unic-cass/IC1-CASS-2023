magic
tech sky130B
magscale 1 2
timestamp 1676037725
<< metal1 >>
tri 7377 3657 7451 3731 se
rect 7451 3657 9696 3731
rect 0 3645 9696 3657
rect 0 3511 7361 3645
tri 7361 3511 7495 3645 nw
tri 8852 3611 8858 3617 se
tri 7593 3545 7659 3611 se
rect 7659 3565 8858 3611
tri 7659 3545 7679 3565 nw
tri 7527 3479 7593 3545 se
tri 7593 3479 7659 3545 nw
tri 7498 3450 7527 3479 se
rect 7527 3450 7564 3479
tri 7564 3450 7593 3479 nw
tri 6891 3427 6914 3450 se
rect 6914 3427 7518 3450
rect 4524 3402 5939 3427
tri 5939 3402 5964 3427 sw
tri 6866 3402 6891 3427 se
rect 6891 3404 7518 3427
tri 7518 3404 7564 3450 nw
rect 6891 3402 6911 3404
rect 4524 3381 6911 3402
tri 6911 3381 6934 3404 nw
tri 4652 3375 4658 3381 nw
tri 5919 3356 5944 3381 ne
rect 5944 3356 6886 3381
tri 6886 3356 6911 3381 nw
rect 9608 3199 9656 3237
tri 9622 3165 9656 3199 ne
tri 9656 3198 9695 3237 sw
rect 9656 3165 9709 3198
tri 7200 3093 7262 3155 se
rect 7262 3103 8720 3155
tri 9656 3112 9709 3165 ne
tri 9709 3152 9741 3184 sw
tri 10813 3152 10831 3170 se
rect 10831 3152 11287 3170
rect 9709 3112 11287 3152
tri 9709 3108 9713 3112 ne
rect 9713 3108 11287 3112
tri 7262 3093 7272 3103 nw
tri 7186 3079 7200 3093 se
rect 7200 3079 7211 3093
rect 6705 3042 7211 3079
tri 7211 3042 7262 3093 nw
tri 10765 3042 10831 3108 ne
rect 10831 3042 11287 3108
rect 6705 3027 7196 3042
tri 7196 3027 7211 3042 nw
rect 0 2833 11255 2999
rect 0 2797 851 2833
tri 851 2797 887 2833 nw
tri 1001 2797 1037 2833 ne
rect 1037 2797 11255 2833
tri 9550 2772 9575 2797 ne
tri 9627 2772 9652 2797 nw
tri 9627 2689 9652 2714 sw
tri 10118 2689 10155 2726 se
rect 9881 2637 10202 2689
rect 0 2428 9600 2473
tri 9600 2428 9645 2473 sw
tri 9811 2428 9856 2473 se
rect 9856 2428 11256 2473
rect 0 2271 11256 2428
rect -1317 1995 -1271 2136
rect -1137 2094 -1093 2136
tri -1093 2094 -1033 2154 sw
tri -918 2149 -824 2243 sw
rect 9642 2177 9770 2229
tri 9770 2177 9822 2229 sw
rect -918 2136 -824 2149
tri -891 2099 -854 2136 ne
rect -854 2135 -824 2136
tri -824 2135 -810 2149 sw
tri -1271 1995 -1206 2060 sw
rect -1137 2048 -893 2094
tri -993 2000 -945 2048 ne
rect -1317 1949 -1055 1995
rect -945 1965 -893 2048
tri -1080 1924 -1055 1949 ne
tri -1083 1810 -1053 1840 sw
tri -941 1810 -854 1897 se
rect -854 1849 -810 2135
rect 5927 2097 6439 2147
tri 6439 2097 6489 2147 sw
rect 7943 2146 8718 2149
tri 8718 2146 8721 2149 sw
tri 9449 2146 9452 2149 se
rect 9452 2146 9642 2149
rect 7943 2097 9642 2146
tri 9752 2107 9822 2177 ne
tri 9822 2150 9849 2177 sw
rect 9822 2107 9928 2150
tri 9822 2098 9831 2107 ne
rect 9831 2098 9928 2107
rect 5927 2095 6489 2097
tri 6417 2069 6443 2095 ne
rect 6443 2069 6489 2095
tri 6489 2069 6517 2097 sw
tri 10842 2069 10904 2131 se
tri 6443 2017 6495 2069 ne
rect 6495 2017 10904 2069
rect -854 1810 -849 1849
tri -849 1810 -810 1849 nw
tri -191 1810 -141 1860 se
tri -141 1810 -93 1858 nw
tri 8777 1834 8802 1859 ne
tri 9228 1834 9253 1859 nw
tri 11458 1831 11492 1865 se
rect -1083 1765 -894 1810
tri -894 1765 -849 1810 nw
tri -241 1760 -191 1810 se
tri -191 1760 -141 1810 nw
rect 9518 1779 9637 1831
tri 9637 1779 9689 1831 sw
rect 11223 1785 11492 1831
tri -291 1710 -241 1760 se
tri -241 1710 -191 1760 nw
tri -341 1660 -291 1710 se
tri -291 1660 -241 1710 nw
rect 1941 1672 3200 1724
tri -391 1610 -341 1660 se
tri -341 1610 -291 1660 nw
tri 3178 1650 3200 1672 ne
tri 3200 1657 3267 1724 sw
rect 7497 1704 7869 1756
tri 9337 1754 9362 1779 nw
tri 9615 1705 9689 1779 ne
tri 9689 1705 9763 1779 sw
tri 9804 1754 9829 1779 ne
rect 3200 1650 3267 1657
tri -441 1560 -391 1610 se
tri -391 1560 -341 1610 nw
tri -466 1535 -441 1560 se
rect -441 1535 -430 1560
tri -1456 1401 -1337 1520 ne
rect -1337 1169 -650 1520
tri -1378 1102 -1337 1143 sw
tri -516 1138 -466 1188 se
rect -466 1174 -430 1535
tri -430 1521 -391 1560 nw
rect 244 1539 290 1607
tri 3200 1583 3267 1650 ne
tri 3267 1583 3341 1657 sw
rect 6907 1607 7010 1628
tri 7010 1607 7031 1628 sw
rect 7497 1608 7552 1704
tri 7552 1653 7603 1704 nw
tri 9260 1675 9285 1700 se
tri 9337 1675 9362 1700 sw
tri 9689 1637 9757 1705 ne
rect 9757 1689 9763 1705
tri 9763 1689 9779 1705 sw
tri 9804 1689 9829 1714 se
rect 9757 1637 9881 1689
tri 244 1493 290 1539 ne
tri 290 1529 328 1567 sw
tri 3267 1531 3319 1583 ne
rect 3319 1531 3550 1583
rect 6907 1576 7031 1607
tri 6988 1533 7031 1576 ne
tri 7031 1533 7105 1607 sw
tri 9404 1598 9429 1623 ne
tri 9481 1598 9506 1623 nw
tri 9804 1612 9829 1637 ne
tri 9404 1533 9429 1558 se
tri 9481 1533 9506 1558 sw
tri 9804 1533 9829 1558 se
rect 290 1493 328 1529
tri 290 1455 328 1493 ne
tri 328 1455 402 1529 sw
tri 328 1403 380 1455 ne
rect 380 1403 1166 1455
tri 6775 1453 6810 1488 se
tri 6862 1453 6897 1488 sw
tri 7031 1481 7083 1533 ne
rect 7083 1481 9541 1533
rect 6159 1401 7277 1453
tri -466 1138 -430 1174 nw
tri 8502 1152 8565 1215 se
rect 8565 1169 8899 1215
tri 8565 1152 8582 1169 nw
tri 8491 1141 8502 1152 se
tri -552 1102 -516 1138 se
rect -516 1102 -502 1138
tri -502 1102 -466 1138 nw
rect -1378 1066 -538 1102
tri -538 1066 -502 1102 nw
rect 6256 1079 7255 1125
tri 7255 1079 7301 1125 sw
tri 7891 1096 7936 1141 se
rect 7936 1096 8502 1141
tri 7874 1079 7891 1096 se
rect 7891 1089 8502 1096
tri 8502 1089 8565 1152 nw
rect 10663 1150 11287 1196
tri 8904 1109 8942 1147 se
rect 7891 1079 7912 1089
rect 6256 1073 7301 1079
tri 7233 1009 7297 1073 ne
rect 7297 1022 7301 1073
tri 7301 1022 7358 1079 sw
tri 7817 1022 7874 1079 se
rect 7874 1055 7912 1079
tri 7912 1055 7946 1089 nw
tri 8638 1055 8692 1109 se
rect 8692 1071 8942 1109
tri 11225 1088 11287 1150 ne
tri 8692 1055 8708 1071 nw
rect 7874 1022 7879 1055
tri 7879 1022 7912 1055 nw
rect 7297 1009 7827 1022
rect -1395 885 -1361 942
tri -775 940 -718 997 sw
rect -775 910 -595 940
tri -595 910 -565 940 sw
tri -1395 851 -1361 885 ne
tri -1361 856 -1317 900 sw
rect -775 894 -565 910
tri -615 856 -577 894 ne
rect -577 856 -565 894
rect -1361 851 -1317 856
tri -1361 826 -1336 851 ne
rect -1336 826 -1317 851
tri -1317 826 -1287 856 sw
rect -1061 828 -624 856
tri -624 828 -596 856 sw
tri -577 844 -565 856 ne
tri -565 844 -499 910 sw
tri -1336 777 -1287 826 ne
tri -1287 777 -1238 826 sw
tri -1287 762 -1272 777 ne
rect -1272 669 -1238 777
rect -1061 810 -596 828
rect -1061 757 -1009 810
tri -1009 771 -970 810 nw
tri -757 718 -709 766 sw
tri -644 762 -596 810 ne
tri -596 809 -577 828 sw
tri -565 809 -530 844 ne
rect -530 809 -499 844
rect -596 762 -577 809
tri -577 762 -530 809 sw
tri -530 778 -499 809 ne
tri -499 778 -433 844 sw
tri -317 778 -290 805 se
rect -290 779 -244 991
rect -290 778 -245 779
tri -245 778 -244 779 nw
tri -596 718 -552 762 ne
rect -552 732 -530 762
tri -530 732 -500 762 sw
tri -499 732 -453 778 ne
rect -453 732 -291 778
tri -291 732 -245 778 nw
rect -552 718 -500 732
rect -757 688 -592 718
tri -592 688 -562 718 sw
tri -552 688 -522 718 ne
rect -522 696 -500 718
tri -500 696 -464 732 sw
tri -163 696 -131 728 se
rect -131 708 -85 991
tri 7297 970 7336 1009 ne
rect 7336 970 7827 1009
tri 7827 970 7879 1022 nw
tri 8592 1009 8638 1055 se
rect 8638 1009 8646 1055
tri 8646 1009 8692 1055 nw
tri 8920 1049 8942 1071 ne
rect 8163 957 8594 1009
tri 8594 957 8646 1009 nw
tri 8735 949 8801 1015 se
rect 8801 969 9720 1015
tri 8801 949 8821 969 nw
tri 8709 923 8735 949 se
rect 8735 923 8775 949
tri 8775 923 8801 949 nw
rect 8664 877 8729 923
tri 8729 877 8775 923 nw
rect -131 696 -97 708
tri -97 696 -85 708 nw
rect -522 688 -143 696
tri -1238 669 -1224 683 sw
rect -757 672 -562 688
tri -1272 621 -1224 669 ne
tri -1224 621 -1176 669 sw
tri -757 652 -737 672 nw
tri -612 622 -562 672 ne
tri -562 650 -524 688 sw
tri -522 650 -484 688 ne
rect -484 650 -143 688
tri -143 650 -97 696 nw
rect -562 622 -524 650
tri -524 622 -496 650 sw
tri -1224 587 -1190 621 ne
rect -1190 592 -609 621
tri -609 592 -580 621 sw
rect -1190 587 -580 592
tri -623 544 -580 587 ne
tri -580 576 -564 592 sw
tri -562 576 -516 622 ne
rect -516 576 -253 622
rect -580 544 -564 576
tri -564 544 -532 576 sw
tri 1899 544 1917 562 se
tri 4968 544 5011 587 se
rect 5011 544 5799 587
tri -580 510 -546 544 ne
rect -546 528 1035 544
tri 1035 528 1051 544 sw
tri 1281 528 1297 544 se
rect 1297 528 1917 544
rect -546 510 1917 528
rect 2892 535 5799 544
rect 2892 510 5008 535
tri 5008 510 5033 535 nw
tri 1021 494 1037 510 ne
rect 1037 494 1290 510
tri 1290 494 1306 510 nw
tri 3006 492 3024 510 nw
tri -1083 101 -1048 136 sw
rect -1083 55 -986 101
tri -1083 21 -1049 55 nw
rect -1321 -95 -1275 -28
tri -1275 -95 -1255 -75 sw
tri -1321 -161 -1255 -95 ne
tri -1255 -161 -1189 -95 sw
tri -1359 -253 -1308 -202 sw
tri -1255 -223 -1193 -161 ne
rect -1193 -177 -1189 -161
tri -1189 -177 -1173 -161 sw
rect -1193 -223 -1128 -177
tri -751 -253 -731 -233 se
rect -731 -253 2674 -233
rect -1359 -285 2674 -253
rect -1359 -305 -729 -285
tri -729 -305 -709 -285 nw
rect -1359 -311 -1354 -305
tri -1354 -311 -1348 -305 nw
tri -1300 -341 -1294 -335 se
rect -1294 -387 -1184 -335
<< metal2 >>
tri 8858 3534 8889 3565 ne
tri 4524 3328 4571 3375 ne
tri 4524 3189 4571 3236 se
rect 4571 3189 4627 3375
tri 4627 3350 4652 3375 nw
tri 8720 3286 8796 3362 ne
tri 4627 3189 4652 3214 sw
tri 8720 3155 8796 3231 se
rect 8796 3155 8848 3362
tri 3550 3089 3598 3137 ne
tri -1593 2447 -1511 2529 se
rect -1593 2343 -1511 2447
rect -1593 179 -1441 2343
tri -1441 2279 -1377 2343 nw
rect -945 1294 -893 1969
rect -141 1809 -89 1858
tri -89 1809 -67 1831 sw
tri -141 1735 -67 1809 ne
tri -67 1746 -4 1809 sw
rect -67 1735 -4 1746
tri -67 1724 -56 1735 ne
rect -56 1660 -4 1735
tri 1941 1643 1970 1672 ne
tri -945 1242 -893 1294 ne
tri -893 1272 -849 1316 sw
rect -893 1242 -849 1272
tri -893 1198 -849 1242 ne
tri -849 1198 -775 1272 sw
tri -849 1176 -827 1198 ne
rect -827 1022 -775 1198
tri 1917 562 1970 615 se
rect 1970 562 2033 1672
tri 2033 1643 2062 1672 nw
tri 3550 1583 3598 1631 se
rect 3598 1583 3646 3137
tri 3646 3105 3678 3137 nw
rect 8720 3103 8848 3155
tri 8720 3027 8796 3103 ne
tri 6680 3002 6705 3027 ne
tri 5799 2053 5841 2095 ne
tri 3646 1583 3678 1615 sw
tri 5799 587 5841 629 se
rect 5841 587 5894 2095
tri 5894 2062 5927 2095 nw
tri 7891 1756 7944 1809 se
rect 7944 1756 7991 2097
tri 7991 2044 8044 2097 nw
rect 8489 1954 8617 2017
tri 8395 1826 8489 1920 se
tri 8489 1826 8617 1954 nw
tri 7991 1756 7997 1762 sw
tri 6757 1708 6782 1733 sw
tri 8301 1732 8395 1826 se
tri 8395 1732 8489 1826 nw
tri 8233 1664 8301 1732 se
rect 8301 1664 8327 1732
tri 8327 1664 8395 1732 nw
tri 7437 1549 7497 1609 se
rect 7497 1587 7549 1608
rect 7497 1549 7511 1587
tri 7511 1549 7549 1587 nw
rect 6804 1214 6865 1529
tri 7363 1475 7437 1549 se
tri 7437 1475 7511 1549 nw
tri 7341 1453 7363 1475 se
rect 7277 1401 7363 1453
tri 7363 1401 7437 1475 nw
tri 6865 1215 6932 1282 sw
tri 8024 1205 8035 1216 ne
tri 6327 1048 6352 1073 nw
rect 8035 1009 8163 1216
tri 8163 1201 8178 1216 nw
tri 5894 587 5927 620 sw
tri 2033 562 2045 574 sw
tri 2879 449 2922 492 ne
tri 2852 -165 2922 -95 se
rect 2922 -112 2975 492
tri 2975 461 3006 492 nw
rect 7973 303 8131 848
tri 8208 458 8233 483 se
rect 8233 406 8300 1664
tri 8300 1637 8327 1664 nw
tri 8692 1598 8717 1623 nw
tri 8771 1453 8796 1478 se
rect 8796 1453 8848 3103
tri 8831 1335 8889 1393 se
rect 8889 1375 8929 3565
tri 8929 3533 8961 3565 nw
tri 9366 3519 9401 3554 se
rect 9401 3519 9754 3554
tri 9754 3519 9789 3554 sw
tri 9346 3499 9366 3519 se
rect 9366 3510 9789 3519
rect 9366 3499 9390 3510
rect 9346 3332 9390 3499
tri 9390 3481 9419 3510 nw
tri 9736 3457 9789 3510 ne
tri 9789 3413 9895 3519 sw
tri 9390 3332 9452 3394 sw
tri 9574 3332 9604 3362 ne
rect 9346 3319 9495 3332
tri 9346 3287 9378 3319 ne
rect 9378 3287 9495 3319
tri 9456 3248 9495 3287 ne
tri 9581 3248 9604 3271 se
rect 9604 3248 9670 3362
tri 9670 3248 9709 3287 sw
tri 9616 2703 9682 2769 se
rect 9682 2717 9755 2769
tri 9682 2703 9696 2717 nw
tri 9588 2675 9616 2703 se
rect 9616 2675 9634 2703
tri 9549 2504 9588 2543 se
rect 9588 2451 9634 2675
tri 9634 2655 9682 2703 nw
tri 9804 2612 9829 2637 ne
tri 9514 2169 9522 2177 ne
rect 9522 2007 9574 2177
tri 9574 2151 9600 2177 nw
tri 9642 2068 9671 2097 ne
rect 9671 2067 9740 2097
tri 9522 1955 9574 2007 ne
tri 9574 1967 9636 2029 sw
rect 9574 1955 9636 1967
tri 9574 1945 9584 1955 ne
tri 9559 1831 9584 1856 se
rect 9584 1779 9636 1955
tri 8988 1379 9062 1453 se
rect 9062 1401 9162 1453
tri 9062 1379 9084 1401 nw
tri 8889 1335 8929 1375 nw
tri 8790 1294 8831 1335 se
rect 8831 1294 8848 1335
tri 8848 1294 8889 1335 nw
tri 8942 1333 8988 1379 se
rect 8988 1333 8994 1379
rect 8790 1039 8830 1294
tri 8830 1276 8848 1294 nw
rect 8942 1177 8994 1333
tri 8994 1311 9062 1379 nw
rect 9671 1116 9723 2067
tri 9723 2050 9740 2067 nw
tri 9804 1831 9829 1856 se
rect 9829 1779 9881 2689
tri 9928 2150 10000 2222 se
rect 10000 2150 10052 2724
tri 10052 2150 10056 2154 sw
tri 10881 1831 10904 1854 se
rect 10904 1831 10956 2017
tri 10956 1831 11009 1884 sw
tri 9723 1116 9799 1192 sw
tri 8830 1039 8848 1057 sw
tri 8790 981 8848 1039 ne
tri 8848 981 8906 1039 sw
tri 8848 965 8864 981 ne
tri 8692 928 8717 953 sw
rect 8864 932 8906 981
tri 8906 932 8955 981 sw
tri 8131 303 8184 356 sw
rect 7973 244 8392 303
tri 7973 145 8072 244 ne
rect 8072 145 8392 244
tri 6327 92 6352 117 sw
tri 2922 -165 2975 -112 nw
tri 2784 -233 2852 -165 se
rect 2852 -233 2854 -165
tri 2854 -233 2922 -165 nw
rect 2674 -285 2802 -233
tri 2802 -285 2854 -233 nw
tri -1236 -335 -1206 -305 se
tri -1159 -335 -1129 -305 sw
tri -1236 -408 -1215 -387 ne
tri -1159 -417 -1129 -387 nw
<< metal3 >>
tri -907 2352 -817 2442 ne
tri -1258 1173 -1220 1211 ne
rect -1220 -267 -1154 1211
tri -1154 1159 -1102 1211 nw
rect -817 776 -751 2442
use sky130_fd_io__com_pdpredrvr_pbiasv2  sky130_fd_io__com_pdpredrvr_pbiasv2_0
timestamp 1676037725
transform -1 0 20068 0 1 -2980
box 11368 2942 20000 5606
use sky130_fd_io__gpiov2_octl_mux  sky130_fd_io__gpiov2_octl_mux_0
timestamp 1676037725
transform 1 0 -1627 0 -1 3513
box 1191 1040 1945 3147
use sky130_fd_io__gpiov2_pdpredrvr_strong_nr2  sky130_fd_io__gpiov2_pdpredrvr_strong_nr2_0
timestamp 1676037725
transform 1 0 3465 0 -1 -331
box 4776 -2127 7821 -314
use sky130_fd_io__gpiov2_pdpredrvr_strong_nr3  sky130_fd_io__gpiov2_pdpredrvr_strong_nr3_0
timestamp 1676037725
transform -1 0 12458 0 1 3202
box 1161 -1273 3472 675
use sky130_fd_io__hvsbt_inv_x1  sky130_fd_io__hvsbt_inv_x1_0
timestamp 1676037725
transform -1 0 -1117 0 -1 418
box 107 226 240 873
use sky130_fd_io__hvsbt_inv_x1  sky130_fd_io__hvsbt_inv_x1_1
timestamp 1676037725
transform -1 0 -1117 0 -1 2582
box 107 226 240 873
use sky130_fd_io__hvsbt_nand2  sky130_fd_io__hvsbt_nand2_0
timestamp 1676037725
transform 1 0 -1299 0 -1 418
box 107 226 460 873
use sky130_fd_io__hvsbt_nand2  sky130_fd_io__hvsbt_nand2_1
timestamp 1676037725
transform 1 0 -1299 0 -1 2582
box 107 226 460 873
use sky130_fd_io__tk_em1o_cdns_5595914180880  sky130_fd_io__tk_em1o_cdns_5595914180880_0
timestamp 1676037725
transform 0 1 9429 1 0 1506
box 0 0 1 1
use sky130_fd_io__tk_em1o_cdns_5595914180880  sky130_fd_io__tk_em1o_cdns_5595914180880_1
timestamp 1676037725
transform 0 1 9829 -1 0 1806
box 0 0 1 1
use sky130_fd_io__tk_em1o_cdns_5595914180880  sky130_fd_io__tk_em1o_cdns_5595914180880_2
timestamp 1676037725
transform 1 0 9509 0 1 1481
box 0 0 1 1
use sky130_fd_io__tk_em1s_cdns_5595914180882  sky130_fd_io__tk_em1s_cdns_5595914180882_0
timestamp 1676037725
transform -1 0 9455 0 -1 1675
box 0 0 1 1
use sky130_fd_io__tk_em1s_cdns_5595914180882  sky130_fd_io__tk_em1s_cdns_5595914180882_1
timestamp 1676037725
transform 0 -1 9627 1 0 2680
box 0 0 1 1
use sky130_fd_io__tk_em1s_cdns_5595914180882  sky130_fd_io__tk_em1s_cdns_5595914180882_2
timestamp 1676037725
transform -1 0 9518 0 1 1779
box 0 0 1 1
use sky130_fd_pr__model__nfet_highvoltage__example_55959141808139  sky130_fd_pr__model__nfet_highvoltage__example_55959141808139_0
timestamp 1676037725
transform 1 0 8867 0 1 1623
box -15 0 311 1
use sky130_fd_pr__model__nfet_highvoltage__example_55959141808183  sky130_fd_pr__model__nfet_highvoltage__example_55959141808183_0
timestamp 1676037725
transform 1 0 9247 0 1 1623
box -15 0 121 1
use sky130_fd_pr__model__nfet_highvoltage__example_55959141808369  sky130_fd_pr__model__nfet_highvoltage__example_55959141808369_0
timestamp 1676037725
transform 1 0 -1093 0 -1 596
box -1 0 121 1
use sky130_fd_pr__model__nfet_highvoltage__example_55959141808643  sky130_fd_pr__model__nfet_highvoltage__example_55959141808643_0
timestamp 1676037725
transform 1 0 -1373 0 -1 540
box -1 0 101 1
use sky130_fd_pr__model__pfet_highvoltage__example_55959141808141  sky130_fd_pr__model__pfet_highvoltage__example_55959141808141_0
timestamp 1676037725
transform 1 0 8867 0 -1 1363
box -15 0 -14 1
use sky130_fd_pr__model__pfet_highvoltage__example_55959141808141  sky130_fd_pr__model__pfet_highvoltage__example_55959141808141_1
timestamp 1676037725
transform -1 0 9163 0 -1 1363
box -15 0 -14 1
use sky130_fd_pr__model__pfet_highvoltage__example_55959141808184  sky130_fd_pr__model__pfet_highvoltage__example_55959141808184_0
timestamp 1676037725
transform 1 0 9247 0 -1 1363
box -15 0 121 1
use sky130_fd_pr__model__pfet_highvoltage__example_55959141808371  sky130_fd_pr__model__pfet_highvoltage__example_55959141808371_0
timestamp 1676037725
transform 1 0 -1093 0 -1 994
box -1 0 121 1
use sky130_fd_pr__model__pfet_highvoltage__example_55959141808371  sky130_fd_pr__model__pfet_highvoltage__example_55959141808371_1
timestamp 1676037725
transform 1 0 -1093 0 1 1062
box -1 0 121 1
use sky130_fd_pr__model__pfet_highvoltage__example_55959141808642  sky130_fd_pr__model__pfet_highvoltage__example_55959141808642_0
timestamp 1676037725
transform 1 0 -1373 0 -1 1394
box -1 0 101 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_0
timestamp 1676037725
transform 0 -1 -1228 -1 0 539
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_1
timestamp 1676037725
transform 0 -1 -1104 -1 0 539
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_2
timestamp 1676037725
transform 0 -1 -1104 1 0 1184
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_3
timestamp 1676037725
transform 0 -1 9222 -1 0 836
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_4
timestamp 1676037725
transform 1 0 9049 0 -1 1441
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_5
timestamp 1676037725
transform 1 0 8876 0 -1 1441
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_6
timestamp 1676037725
transform 0 1 9188 1 0 1741
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_7
timestamp 1676037725
transform 0 1 8808 1 0 1741
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_8
timestamp 1676037725
transform 1 0 8781 0 -1 1209
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_9
timestamp 1676037725
transform 1 0 6225 0 1 52
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_10
timestamp 1676037725
transform 1 0 9363 0 -1 1523
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_11
timestamp 1676037725
transform 0 -1 8726 -1 0 836
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_0
timestamp 1676037725
transform 1 0 9508 0 1 1779
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_1
timestamp 1676037725
transform -1 0 9881 0 1 2637
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_2
timestamp 1676037725
transform -1 0 9881 0 1 1779
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_3
timestamp 1676037725
transform -1 0 8848 0 1 1401
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_4
timestamp 1676037725
transform 1 0 6256 0 1 40
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_5
timestamp 1676037725
transform 1 0 6256 0 1 1073
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_6
timestamp 1676037725
transform 1 0 8172 0 1 406
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_7
timestamp 1676037725
transform 1 0 8628 0 1 876
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_8
timestamp 1676037725
transform 1 0 8628 0 1 1623
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_9
timestamp 1676037725
transform 1 0 6629 0 1 3027
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_10
timestamp 1676037725
transform 1 0 6705 0 1 1656
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_0
timestamp 1676037725
transform 0 -1 -999 -1 0 762
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_1
timestamp 1676037725
transform 0 1 8894 1 0 1395
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_2
timestamp 1676037725
transform 0 1 9070 1 0 1395
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_3
timestamp 1676037725
transform 0 1 9247 1 0 1395
box 0 0 1 1
<< properties >>
string GDS_END 49062696
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 49014006
<< end >>
