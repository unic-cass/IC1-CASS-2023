magic
tech sky130B
magscale 1 2
timestamp 1676037725
<< metal1 >>
rect 235 3186 2717 3214
tri 235 3162 259 3186 nw
tri 2693 3162 2717 3186 ne
tri 3235 3194 3241 3200 sw
rect 3235 3171 5474 3194
tri 5474 3171 5497 3194 sw
rect 3235 3160 5497 3171
tri 3235 3148 3247 3160 nw
rect 2605 3120 2607 3138
tri 2607 3120 2625 3138 sw
rect 2479 3099 5416 3120
tri 5416 3099 5437 3120 sw
tri 5454 3117 5497 3160 ne
tri 5497 3117 5551 3171 sw
rect 2479 3086 5437 3099
rect 5383 3052 5437 3086
tri 5497 3083 5531 3117 ne
rect 5531 3083 6021 3117
rect 5967 2987 6021 3083
tri 2179 2793 2203 2817 sw
rect 2179 2765 3322 2793
tri 2415 2532 2447 2564 ne
tri 2499 2532 2531 2564 nw
rect 2837 2563 4642 2607
tri 2883 2529 2917 2563 nw
tri 4634 2555 4642 2563 ne
rect 934 2487 2268 2515
tri 922 2416 962 2456 se
rect 962 2428 1214 2456
tri 962 2416 974 2428 nw
tri 921 2415 922 2416 se
rect 922 2415 944 2416
rect 785 2398 944 2415
tri 944 2398 962 2416 nw
rect 785 2369 915 2398
tri 915 2369 944 2398 nw
rect 1068 2394 1132 2400
tri 1132 2394 1138 2400 sw
tri 1148 2394 1182 2428 ne
rect 1182 2424 1214 2428
tri 1214 2424 1246 2456 sw
tri 2200 2439 2248 2487 ne
rect 2248 2472 2268 2487
tri 2268 2472 2311 2515 sw
rect 2248 2439 2311 2472
tri 3209 2495 3248 2534 se
rect 3248 2495 3594 2534
rect 3209 2492 3594 2495
rect 3209 2450 3255 2492
tri 3255 2461 3286 2492 nw
tri 3578 2476 3594 2492 ne
tri 3594 2480 3648 2534 sw
tri 4835 2489 4841 2495 se
rect 3594 2476 3648 2480
tri 3594 2464 3606 2476 ne
rect 1182 2406 1246 2424
tri 1356 2398 1390 2432 se
tri 2878 2405 2912 2439 se
rect 1068 2354 1138 2394
tri 1138 2354 1178 2394 sw
tri 2409 2359 2435 2385 se
rect 2435 2362 2502 2393
rect 2435 2359 2453 2362
tri 1123 2299 1178 2354 ne
tri 1178 2299 1233 2354 sw
tri 1365 2327 1390 2352 ne
tri 1840 2313 1886 2359 se
rect 1886 2313 2453 2359
tri 2453 2313 2502 2362 nw
tri 2911 2358 2912 2359 ne
tri 3175 2327 3209 2361 se
tri 1178 2269 1208 2299 ne
rect 1208 2297 1233 2299
tri 1233 2297 1235 2299 sw
tri 1824 2297 1840 2313 se
rect 1840 2297 1852 2313
rect 1208 2285 1852 2297
tri 1852 2285 1880 2313 nw
tri 3596 2297 3606 2307 se
rect 3606 2297 3648 2476
tri 4220 2451 4254 2485 ne
tri 4503 2475 4505 2477 se
rect 4505 2475 4711 2477
tri 4711 2475 4713 2477 sw
tri 4438 2410 4503 2475 se
rect 4503 2431 4713 2475
rect 4350 2409 4503 2410
tri 4503 2409 4525 2431 nw
tri 4691 2409 4713 2431 ne
tri 4713 2409 4779 2475 sw
rect 4350 2388 4482 2409
tri 4482 2388 4503 2409 nw
tri 4713 2389 4733 2409 ne
tri 4510 2335 4544 2369 se
rect 1208 2269 1836 2285
tri 1836 2269 1852 2285 nw
tri 1883 2269 1899 2285 se
rect 1899 2269 2969 2285
tri 1858 2244 1883 2269 se
rect 1883 2257 2969 2269
rect 1883 2244 1899 2257
tri 1899 2244 1912 2257 nw
tri 1855 2241 1858 2244 se
rect 1858 2241 1868 2244
rect 1143 2201 1224 2214
tri 1224 2201 1237 2214 sw
rect 1768 2213 1868 2241
tri 1868 2213 1899 2244 nw
tri 2949 2237 2969 2257 ne
tri 2969 2253 3001 2285 sw
tri 3268 2253 3302 2287 se
tri 3348 2253 3382 2287 sw
tri 3476 2253 3510 2287 se
tri 4132 2276 4169 2313 se
rect 4169 2276 4171 2313
rect 2969 2237 3207 2253
tri 2969 2225 2981 2237 ne
rect 2981 2225 3207 2237
rect 1143 2162 1237 2201
tri 1202 2127 1237 2162 ne
tri 1237 2127 1311 2201 sw
rect 3960 2183 4169 2276
tri 4510 2260 4544 2294 ne
tri 4667 2222 4733 2288 se
rect 4733 2268 4779 2409
tri 4835 2355 4841 2361 ne
tri 4733 2222 4779 2268 nw
tri 4654 2209 4667 2222 se
rect 4667 2209 4708 2222
tri 2779 2127 2803 2151 se
tri 3960 2146 3997 2183 nw
tri 1237 2099 1265 2127 ne
rect 1265 2099 2803 2127
tri 1150 1813 1200 1863 se
rect 1200 1835 2423 1863
tri 3088 1859 3122 1893 ne
tri 3174 1859 3208 1893 nw
tri 3469 1859 3503 1893 ne
tri 3832 1859 3866 1893 nw
tri 1200 1813 1222 1835 nw
tri 1100 1763 1150 1813 se
tri 1150 1763 1200 1813 nw
tri 2399 1811 2423 1835 ne
tri 1072 1735 1100 1763 se
rect 1100 1735 1122 1763
tri 1122 1735 1150 1763 nw
rect 1912 1761 2201 1807
tri 1165 1735 1167 1737 se
rect 1167 1735 1280 1737
tri 754 1590 780 1616 ne
tri 780 1594 842 1656 sw
rect 900 1628 946 1665
rect 780 1590 842 1594
tri 780 1532 838 1590 ne
rect 838 1543 842 1590
tri 842 1543 893 1594 sw
tri 900 1582 946 1628 ne
tri 946 1600 979 1633 sw
tri 1040 1600 1072 1632 se
rect 1072 1610 1100 1735
tri 1100 1713 1122 1735 nw
rect 946 1582 1072 1600
tri 1072 1582 1100 1610 nw
tri 1128 1698 1165 1735 se
rect 1165 1709 1280 1735
rect 1165 1698 1174 1709
tri 1174 1698 1185 1709 nw
tri 946 1572 956 1582 ne
rect 956 1572 1062 1582
tri 1062 1572 1072 1582 nw
tri 1091 1543 1128 1580 se
rect 1128 1564 1156 1698
tri 1156 1680 1174 1698 nw
tri 1242 1671 1280 1709 ne
tri 1280 1685 1332 1737 sw
tri 2175 1735 2201 1761 ne
rect 1280 1671 1381 1685
tri 1280 1603 1348 1671 ne
rect 1348 1616 1381 1671
tri 3168 1666 3202 1700 se
tri 1427 1616 1461 1650 sw
tri 2094 1616 2128 1650 se
tri 2173 1623 2200 1650 sw
rect 2173 1616 2460 1623
tri 2460 1616 2467 1623 sw
tri 2788 1616 2822 1650 se
rect 1128 1543 1135 1564
tri 1135 1543 1156 1564 nw
tri 1230 1560 1264 1594 sw
rect 1348 1591 2893 1616
rect 1348 1588 2140 1591
tri 2140 1588 2143 1591 nw
tri 2421 1588 2424 1591 ne
rect 2424 1588 2893 1591
tri 2152 1560 2153 1561 se
rect 838 1532 1107 1543
tri 838 1515 855 1532 ne
rect 855 1515 1107 1532
tri 1107 1515 1135 1543 nw
rect 1230 1532 2205 1560
tri 4578 1533 4654 1609 se
rect 4654 1587 4708 2209
tri 4708 2197 4733 2222 nw
tri 4654 1533 4708 1587 nw
tri 2119 1498 2153 1532 ne
tri 4530 1485 4578 1533 se
rect 4578 1485 4606 1533
tri 4606 1485 4654 1533 nw
rect 4517 1433 4554 1485
tri 4554 1433 4606 1485 nw
rect 7822 1313 8247 1347
tri 8247 1313 8281 1347 sw
rect 7822 1295 8281 1313
tri 6385 1238 6419 1272 ne
rect 6419 1154 6631 1272
tri 6631 1215 6688 1272 nw
tri 8183 1249 8229 1295 ne
tri 7181 1201 7187 1207 sw
tri 4725 1074 4774 1123 se
rect 4774 1074 4856 1123
tri 4687 1036 4725 1074 se
rect 4725 1036 4753 1074
tri 4753 1036 4791 1074 nw
tri 4621 970 4687 1036 se
tri 4687 970 4753 1036 nw
tri 4555 904 4621 970 se
rect 4621 968 4685 970
tri 4685 968 4687 970 nw
rect 4621 916 4633 968
tri 4633 916 4685 968 nw
tri 4686 916 4738 968 se
rect 4738 916 4806 968
tri 4621 904 4633 916 nw
tri 4535 884 4555 904 se
rect 4555 884 4600 904
rect 4447 883 4600 884
tri 4600 883 4621 904 nw
tri 4666 896 4686 916 se
rect 4686 896 4732 916
tri 4732 896 4752 916 nw
tri 4653 883 4666 896 se
rect 4447 838 4555 883
tri 4555 838 4600 883 nw
tri 4600 830 4653 883 se
rect 4653 830 4666 883
tri 4666 830 4732 896 nw
tri 4580 810 4600 830 se
rect 4447 764 4600 810
tri 4600 764 4666 830 nw
rect 8229 807 8281 1295
tri 2733 729 2747 743 se
rect 2747 729 3154 743
tri 3154 729 3168 743 sw
tri 3483 729 3490 736 se
rect 3490 729 3930 736
tri 2693 689 2733 729 se
rect 2733 715 3168 729
tri 2733 689 2759 715 nw
tri 3142 689 3168 715 ne
tri 3168 689 3208 729 sw
tri 3450 696 3483 729 se
rect 3483 708 3930 729
rect 3483 696 3490 708
tri 3490 696 3502 708 nw
tri 2654 650 2693 689 se
rect 2693 663 2707 689
tri 2707 663 2733 689 nw
tri 2757 673 2771 687 se
rect 2771 673 3130 687
tri 3130 673 3144 687 sw
tri 2747 663 2757 673 se
rect 2757 663 3144 673
tri 3144 663 3154 673 sw
tri 3168 663 3194 689 ne
rect 3194 663 3208 689
rect 2327 649 2693 650
tri 2693 649 2707 663 nw
rect 2327 622 2666 649
tri 2666 622 2693 649 nw
tri 2717 633 2747 663 se
rect 2747 659 3154 663
rect 2747 633 2757 659
tri 2757 633 2783 659 nw
tri 3118 633 3144 659 ne
rect 3144 633 3154 659
tri 3154 633 3184 663 sw
tri 3194 649 3208 663 ne
tri 3208 649 3248 689 sw
tri 3410 656 3450 696 se
tri 3450 656 3490 696 nw
tri 3507 673 3514 680 se
rect 3514 673 3832 680
tri 3490 656 3507 673 se
rect 3507 656 3832 673
tri 3403 649 3410 656 se
rect 3410 649 3415 656
tri 2706 622 2717 633 se
rect 2327 585 2373 622
tri 2677 593 2706 622 se
rect 2706 593 2717 622
tri 2717 593 2757 633 nw
tri 2651 567 2677 593 se
rect 2677 567 2691 593
tri 2691 567 2717 593 nw
tri 2611 527 2651 567 se
tri 2651 527 2691 567 nw
tri 2571 487 2611 527 se
tri 2611 487 2651 527 nw
tri 2531 447 2571 487 se
tri 2571 447 2611 487 nw
rect 3002 480 3111 610
tri 3144 593 3184 633 ne
tri 3184 622 3195 633 sw
tri 3208 622 3235 649 ne
rect 3235 622 3415 649
rect 3184 593 3195 622
tri 3195 593 3224 622 sw
tri 3235 621 3236 622 ne
rect 3236 621 3415 622
tri 3415 621 3450 656 nw
tri 3474 640 3490 656 se
rect 3490 652 3832 656
rect 3490 640 3514 652
tri 3514 640 3526 652 nw
tri 3455 621 3474 640 se
tri 3434 600 3455 621 se
rect 3455 600 3474 621
tri 3474 600 3514 640 nw
tri 3427 593 3434 600 se
rect 3434 593 3439 600
tri 3111 574 3130 593 sw
tri 3184 565 3212 593 ne
rect 3212 565 3439 593
tri 3439 565 3474 600 nw
tri 3111 503 3130 522 nw
tri 8152 503 8186 537 se
tri 8194 503 8229 538 se
tri 8238 503 8272 537 sw
tri 2518 434 2531 447 se
rect 2531 434 2558 447
tri 2558 434 2571 447 nw
rect 2319 406 2530 434
tri 2530 406 2558 434 nw
tri -317 135 -247 205 sw
rect 4331 163 5080 378
tri 5325 341 5359 375 nw
tri 5080 163 5081 164 nw
rect -317 83 872 135
tri 6461 22 6485 46 sw
tri 6461 -304 6485 -280 nw
<< metal2 >>
tri 1985 3324 2000 3339 se
rect 2000 3324 2442 3339
tri 1931 3270 1985 3324 se
rect 1985 3302 2442 3324
tri 2442 3302 2479 3339 sw
tri 1985 3270 2017 3302 nw
tri 1303 2881 1377 2955 se
rect 1377 2903 1555 2955
tri 1377 2881 1399 2903 nw
tri 1533 2881 1555 2903 ne
tri 1555 2882 1628 2955 sw
rect 1555 2881 1628 2882
tri 1239 2817 1303 2881 se
rect 1303 2817 1342 2881
tri 1342 2846 1377 2881 nw
tri 1555 2860 1576 2881 ne
tri 1345 2554 1419 2628 se
rect 1419 2606 1471 2765
tri 1471 2731 1505 2765 nw
tri 1566 2661 1576 2671 se
rect 1576 2661 1628 2881
tri 1897 2817 1931 2851 se
rect 1931 2817 1983 3270
tri 1983 3268 1985 3270 nw
tri 2405 3228 2479 3302 ne
tri 2479 3250 2531 3302 sw
tri 2684 3283 2703 3302 se
rect 2703 3283 3238 3302
tri 3238 3283 3257 3302 sw
rect 2479 3138 2531 3250
tri 2654 3253 2684 3283 se
rect 2684 3268 3257 3283
rect 2684 3253 2688 3268
tri 2531 3138 2565 3172 sw
tri 2619 2890 2654 2925 se
rect 2654 2890 2688 3253
tri 2688 3239 2717 3268 nw
tri 3224 3235 3257 3268 ne
tri 3257 3235 3305 3283 sw
tri 3257 3221 3271 3235 ne
tri 2579 2804 2613 2838 ne
rect 1419 2577 1442 2606
tri 1442 2577 1471 2606 nw
tri 1504 2599 1566 2661 se
tri 1566 2599 1628 2661 nw
tri 1977 2654 2051 2728 se
tri 2051 2654 2162 2765 nw
tri 1970 2647 1977 2654 se
rect 1977 2647 2022 2654
tri 1482 2577 1504 2599 se
tri 1419 2554 1442 2577 nw
tri 1271 2480 1345 2554 se
rect 1345 2525 1390 2554
tri 1390 2525 1419 2554 nw
tri 1442 2537 1482 2577 se
rect 1482 2537 1504 2577
tri 1504 2537 1566 2599 nw
tri 1430 2525 1442 2537 se
tri 1345 2480 1390 2525 nw
tri 1390 2485 1430 2525 se
rect 1430 2485 1442 2525
tri 1197 2406 1271 2480 se
tri 1271 2406 1345 2480 nw
rect 1390 2455 1442 2485
tri 1442 2475 1504 2537 nw
tri 1160 2369 1197 2406 se
rect 1197 2369 1212 2406
tri 1086 2075 1160 2149 se
rect 1160 2127 1212 2369
tri 1212 2347 1271 2406 nw
tri 1436 2141 1470 2175 se
rect 1470 2153 1522 2327
rect 1970 2176 2022 2647
tri 2022 2625 2051 2654 nw
rect 1470 2141 1510 2153
tri 1510 2141 1522 2153 nw
tri 1160 2075 1212 2127 nw
tri 1212 2075 1278 2141 se
rect 1278 2089 1458 2141
tri 1458 2089 1510 2141 nw
tri 1012 2001 1086 2075 se
rect 1086 2047 1132 2075
tri 1132 2047 1160 2075 nw
tri 1204 2067 1212 2075 se
rect 1212 2067 1278 2075
tri 1278 2067 1300 2089 nw
tri 1184 2047 1204 2067 se
rect 1204 2047 1206 2067
tri 1086 2001 1132 2047 nw
tri 982 1971 1012 2001 se
rect 1012 1971 1034 2001
rect 982 1765 1034 1971
tri 1034 1949 1086 2001 nw
tri 1132 1995 1184 2047 se
rect 1184 1995 1206 2047
tri 1206 1995 1278 2067 nw
tri 1058 1545 1132 1619 se
rect 1132 1597 1184 1995
tri 1184 1973 1206 1995 nw
tri 2423 1863 2447 1887 se
rect 2447 1863 2499 2482
tri 2499 1863 2533 1897 sw
rect 2613 1789 2665 2838
tri 2665 2815 2688 2838 nw
rect 2717 2584 2769 3162
tri 2769 3123 2808 3162 nw
tri 3107 3124 3131 3148 ne
rect 2974 2809 3068 2872
tri 3068 2838 3102 2872 nw
tri 2912 2727 2974 2789 se
rect 2974 2727 2986 2809
tri 2986 2727 3068 2809 nw
rect 2912 2486 2964 2727
tri 2964 2705 2986 2727 nw
rect 3131 2647 3183 3148
tri 3183 3096 3235 3148 nw
rect 3271 2968 3305 3235
tri 3305 2968 3309 2972 sw
rect 3271 2958 3309 2968
tri 3271 2920 3309 2958 ne
tri 3309 2920 3357 2968 sw
rect 3591 2920 3998 2924
tri 3998 2920 4002 2924 sw
tri 3309 2872 3357 2920 ne
tri 3357 2872 3405 2920 sw
rect 3591 2872 4002 2920
tri 3357 2824 3405 2872 ne
tri 3405 2824 3453 2872 sw
tri 3976 2846 4002 2872 ne
tri 4002 2846 4076 2920 sw
rect 4920 2882 4972 2974
rect 5026 2955 5156 2970
tri 4972 2882 4994 2904 sw
tri 3405 2790 3439 2824 ne
rect 3439 2790 3958 2824
tri 3131 2595 3183 2647 ne
tri 3183 2598 3254 2669 sw
rect 3183 2595 3254 2598
tri 3183 2576 3202 2595 ne
tri 2833 2058 2874 2099 ne
rect 2874 1967 2931 2099
tri 2874 1910 2931 1967 ne
tri 2931 1952 2963 1984 sw
rect 2931 1910 2963 1952
tri 2931 1878 2963 1910 ne
tri 2963 1878 3037 1952 sw
tri 2963 1856 2985 1878 ne
rect 2985 1744 3037 1878
rect 3202 1786 3254 2595
tri 3297 1861 3308 1872 se
rect 3308 1798 3336 2779
tri 3944 2776 3958 2790 ne
tri 3958 2780 4002 2824 sw
tri 4002 2780 4068 2846 ne
rect 4068 2780 4076 2846
rect 3958 2776 4002 2780
tri 3958 2772 3962 2776 ne
rect 3962 2772 4002 2776
tri 4002 2772 4010 2780 sw
tri 4068 2772 4076 2780 ne
tri 4076 2772 4150 2846 sw
tri 4920 2808 4994 2882 ne
tri 4994 2872 5004 2882 sw
tri 5026 2872 5109 2955 ne
rect 5109 2922 5156 2955
tri 5156 2922 5193 2959 sw
tri 6248 2922 6278 2952 se
rect 6278 2922 6330 2957
rect 5109 2908 6330 2922
rect 5109 2872 6294 2908
tri 6294 2872 6330 2908 nw
rect 4994 2844 5004 2872
tri 5004 2844 5032 2872 sw
tri 6392 2866 6432 2906 se
rect 6432 2884 6484 2957
rect 6432 2866 6466 2884
tri 6466 2866 6484 2884 nw
tri 6370 2844 6392 2866 se
rect 4994 2808 6392 2844
tri 4994 2792 5010 2808 ne
rect 5010 2792 6392 2808
tri 6392 2792 6466 2866 nw
tri 3962 2730 4004 2772 ne
rect 4004 2730 4010 2772
tri 4010 2730 4052 2772 sw
tri 4004 2682 4052 2730 ne
tri 4052 2706 4076 2730 sw
tri 4076 2706 4142 2772 ne
rect 4142 2706 4150 2772
rect 4052 2682 4076 2706
tri 4076 2682 4100 2706 sw
tri 4142 2698 4150 2706 ne
tri 4150 2698 4224 2772 sw
tri 4052 2634 4100 2682 ne
tri 4100 2634 4148 2682 sw
tri 4100 2586 4148 2634 ne
tri 4148 2632 4150 2634 sw
tri 4150 2632 4216 2698 ne
rect 4216 2632 4224 2698
rect 4148 2586 4150 2632
tri 4150 2586 4196 2632 sw
tri 4216 2624 4224 2632 ne
tri 4224 2624 4298 2698 sw
rect 3683 2560 4127 2563
tri 4127 2560 4130 2563 sw
tri 4148 2560 4174 2586 ne
rect 4174 2560 4196 2586
rect 3683 2538 4130 2560
tri 4130 2538 4152 2560 sw
tri 4174 2538 4196 2560 ne
tri 4196 2558 4224 2586 sw
tri 4224 2558 4290 2624 ne
rect 4290 2558 4298 2624
rect 4196 2538 4224 2558
tri 4224 2538 4244 2558 sw
tri 4290 2550 4298 2558 ne
tri 4298 2550 4372 2624 sw
rect 4770 2598 5978 2607
tri 5978 2598 5987 2607 sw
rect 4770 2555 5987 2598
rect 3683 2507 4152 2538
tri 4117 2490 4134 2507 ne
rect 4134 2494 4152 2507
tri 4152 2494 4196 2538 sw
tri 4196 2494 4240 2538 ne
rect 4240 2494 4244 2538
rect 4134 2490 4196 2494
tri 4196 2490 4200 2494 sw
tri 4240 2490 4244 2494 ne
tri 4244 2490 4292 2538 sw
tri 4134 2428 4196 2490 ne
rect 4196 2472 4200 2490
tri 4200 2472 4218 2490 sw
tri 4244 2472 4262 2490 ne
rect 4262 2484 4292 2490
tri 4292 2484 4298 2490 sw
tri 4298 2484 4364 2550 ne
rect 4364 2484 4372 2550
rect 4262 2472 4298 2484
rect 4196 2428 4218 2472
tri 4218 2428 4262 2472 sw
tri 4262 2442 4292 2472 ne
rect 4292 2442 4298 2472
tri 4298 2442 4340 2484 sw
tri 4364 2476 4372 2484 ne
tri 4372 2476 4446 2550 sw
tri 5956 2524 5987 2555 ne
tri 5987 2524 6061 2598 sw
tri 4822 2476 4835 2489 se
tri 4196 2362 4262 2428 ne
tri 4262 2406 4284 2428 sw
tri 4292 2406 4328 2442 ne
rect 4328 2424 4340 2442
tri 4340 2424 4358 2442 sw
tri 4372 2424 4424 2476 ne
rect 4424 2424 4835 2476
tri 5987 2450 6061 2524 ne
tri 6061 2450 6135 2524 sw
rect 4328 2406 4358 2424
rect 4262 2362 4284 2406
tri 4284 2362 4328 2406 sw
tri 4328 2394 4340 2406 ne
rect 4340 2394 4358 2406
tri 4358 2394 4388 2424 sw
tri 4340 2362 4372 2394 ne
rect 4372 2362 4388 2394
tri 3883 2276 3960 2353 sw
tri 4262 2296 4328 2362 ne
tri 4328 2346 4344 2362 sw
tri 4372 2346 4388 2362 ne
tri 4388 2346 4436 2394 sw
tri 4801 2390 4835 2424 ne
tri 6061 2376 6135 2450 ne
tri 6135 2376 6209 2450 sw
rect 4328 2312 4344 2346
tri 4344 2312 4378 2346 sw
tri 4388 2312 4422 2346 ne
rect 4422 2312 4462 2346
rect 4328 2296 4378 2312
tri 4378 2296 4394 2312 sw
tri 3546 2191 3596 2241 ne
rect 3827 2146 3908 2276
tri 4328 2230 4394 2296 ne
tri 4394 2294 4396 2296 sw
tri 4444 2294 4462 2312 ne
tri 6135 2302 6209 2376 ne
tri 6209 2302 6283 2376 sw
rect 4394 2230 4396 2294
tri 4396 2230 4460 2294 sw
tri 6209 2280 6231 2302 ne
tri 4394 2174 4450 2230 ne
rect 4450 2174 6097 2230
tri 6075 2152 6097 2174 ne
tri 6097 2153 6174 2230 sw
rect 6097 2152 6174 2153
tri 6097 2131 6118 2152 ne
tri 3408 2096 3425 2113 ne
tri 3336 1861 3349 1874 sw
rect 3425 1782 3477 2113
tri 3477 2028 3562 2113 nw
tri 3477 1706 3511 1740 sw
rect 3477 1654 5913 1706
tri 1132 1545 1184 1597 nw
tri 998 1485 1058 1545 se
rect 1058 1485 1113 1545
tri 1113 1526 1132 1545 nw
tri -341 211 -317 235 sw
rect 1580 213 1632 1644
tri 4525 1461 4549 1485 sw
rect 4525 1433 4948 1461
rect 2427 1199 2483 1240
tri 2427 1143 2483 1199 ne
tri 2483 1184 2520 1221 sw
rect 4920 1207 4948 1433
rect 6118 1363 6174 2152
rect 6231 1425 6283 2302
tri 6231 1373 6283 1425 ne
tri 6283 1421 6309 1447 sw
rect 6283 1373 6309 1421
tri 6174 1363 6179 1368 sw
rect 6118 1346 6179 1363
tri 6118 1285 6179 1346 ne
tri 6179 1285 6257 1363 sw
tri 6283 1347 6309 1373 ne
tri 6309 1347 6383 1421 sw
tri 6309 1295 6361 1347 ne
rect 6361 1295 7702 1347
tri 6179 1207 6257 1285 ne
tri 6257 1207 6335 1285 sw
rect 2483 1143 2520 1184
tri 2483 1106 2520 1143 ne
tri 2520 1106 2598 1184 sw
tri 6257 1155 6309 1207 ne
rect 6309 1155 7043 1207
tri 7609 1124 7610 1125 se
rect 7610 1124 7803 1125
tri 2520 1050 2576 1106 ne
rect 2576 1050 3157 1106
rect 4871 1073 7803 1124
rect 4871 1072 7631 1073
tri 7631 1072 7632 1073 nw
tri 3109 1002 3157 1050 ne
tri 7489 968 7490 969 se
rect 7490 968 7803 969
rect 4871 917 7803 968
rect 4871 916 7623 917
tri 7623 916 7624 917 nw
rect 4871 815 7615 818
tri 7615 815 7618 818 sw
rect 4871 766 7798 815
tri 7593 763 7596 766 ne
rect 7596 763 7798 766
rect 8229 696 8281 769
rect 4871 659 7687 663
tri 7687 659 7691 663 sw
rect 4871 611 7804 659
tri 8229 644 8281 696 ne
tri 8281 690 8309 718 sw
rect 8281 644 8309 690
tri 8281 616 8309 644 ne
tri 8309 616 8383 690 sw
tri 7665 607 7669 611 ne
rect 7669 607 7804 611
tri 8309 564 8361 616 ne
rect 8361 591 8578 616
tri 8578 591 8603 616 sw
rect 8361 564 8603 591
tri 8556 517 8603 564 ne
tri 8603 517 8677 591 sw
tri 8603 495 8625 517 ne
tri 8118 371 8186 439 se
rect 8186 417 8238 449
rect 8186 371 8192 417
tri 8192 371 8238 417 nw
tri 1632 213 1675 256 sw
tri 4094 213 4128 247 se
rect 1580 202 4184 213
tri 1580 161 1621 202 ne
rect 1621 161 4184 202
tri -341 59 -317 83 nw
tri 872 17 938 83 ne
rect 938 -80 970 83
tri 970 53 1000 83 nw
tri 3213 -34 3296 49 sw
tri 6485 -16 6519 18 sw
tri 8044 -11 8118 63 se
rect 8118 41 8170 371
tri 8170 349 8192 371 nw
tri 8118 -11 8170 41 nw
tri 8039 -16 8044 -11 se
rect 8044 -16 8061 -11
tri 938 -112 970 -80 ne
tri 970 -108 1012 -66 sw
rect 3213 -86 5865 -34
tri 3213 -105 3232 -86 nw
tri 5843 -108 5865 -86 ne
tri 5865 -105 5936 -34 sw
rect 6485 -68 8061 -16
tri 8061 -68 8118 -11 nw
tri 8551 -31 8625 43 se
rect 8625 21 8677 517
tri 8625 -31 8677 21 nw
tri 6485 -102 6519 -68 nw
tri 8477 -105 8551 -31 se
tri 8551 -105 8625 -31 nw
rect 5865 -108 5936 -105
rect 970 -112 1012 -108
tri 970 -148 1006 -112 ne
rect 1006 -148 1012 -112
tri 1012 -148 1052 -108 sw
tri 1006 -194 1052 -148 ne
tri 1052 -194 1098 -148 sw
tri 5865 -173 5930 -108 ne
rect 5930 -173 5936 -108
tri 5936 -173 6004 -105 sw
tri 8430 -152 8477 -105 se
rect 8477 -152 8504 -105
tri 8504 -152 8551 -105 nw
tri 1052 -240 1098 -194 ne
tri 1098 -240 1144 -194 sw
tri 1098 -286 1144 -240 ne
tri 1144 -286 1190 -240 sw
tri 5930 -247 6004 -173 ne
tri 6004 -247 6078 -173 sw
rect 6485 -204 8452 -152
tri 8452 -204 8504 -152 nw
tri 6485 -238 6519 -204 nw
tri 1144 -318 1176 -286 ne
rect 1176 -300 1324 -286
tri 1324 -300 1338 -286 sw
rect 1176 -318 1338 -300
tri 1310 -346 1338 -318 ne
tri 1338 -346 1384 -300 sw
tri 6004 -321 6078 -247 ne
tri 6078 -321 6152 -247 sw
tri 6400 -321 6433 -288 se
rect 6433 -310 6485 -280
rect 6433 -321 6474 -310
tri 6474 -321 6485 -310 nw
tri 1338 -392 1384 -346 ne
tri 1384 -392 1430 -346 sw
tri 6078 -373 6130 -321 ne
rect 6130 -373 6422 -321
tri 6422 -373 6474 -321 nw
tri 1384 -438 1430 -392 ne
tri 1430 -438 1476 -392 sw
tri 1430 -484 1476 -438 ne
tri 1476 -484 1522 -438 sw
tri 1476 -530 1522 -484 ne
tri 1522 -530 1568 -484 sw
tri 1522 -576 1568 -530 ne
tri 1568 -576 1614 -530 sw
tri 1568 -622 1614 -576 ne
tri 1614 -622 1660 -576 sw
tri 1614 -668 1660 -622 ne
tri 1660 -668 1706 -622 sw
tri 1660 -714 1706 -668 ne
tri 1706 -714 1752 -668 sw
tri 1706 -760 1752 -714 ne
tri 1752 -760 1798 -714 sw
tri 2186 -760 2250 -696 se
tri 1752 -792 1784 -760 ne
rect 1784 -792 2306 -760
<< metal3 >>
rect 3068 2502 3533 2568
tri 3068 2468 3102 2502 nw
tri 3180 2336 3274 2430 se
rect 3274 2364 3888 2430
tri 3274 2336 3302 2364 nw
tri 3161 2317 3180 2336 se
rect 3180 2317 3189 2336
tri 2609 2223 2703 2317 se
rect 2703 2251 3189 2317
tri 3189 2251 3274 2336 nw
tri 3778 2320 3822 2364 ne
rect 3822 2360 3888 2364
rect 3644 2252 3648 2302
tri 3648 2252 3698 2302 sw
tri 2703 2223 2731 2251 nw
rect 3644 2236 3698 2252
tri 2515 2129 2609 2223 se
tri 2609 2129 2703 2223 nw
tri 2421 2035 2515 2129 se
tri 2515 2035 2609 2129 nw
tri 2839 2080 2933 2174 se
rect 2933 2108 3412 2174
tri 3620 2158 3698 2236 ne
tri 3698 2158 3792 2252 sw
tri 2933 2080 2961 2108 nw
tri 2419 2033 2421 2035 se
rect 2421 2033 2485 2035
rect 2192 1622 2258 1668
rect 2419 1663 2485 2033
tri 2485 2005 2515 2035 nw
tri 2745 1986 2839 2080 se
tri 2839 1986 2933 2080 nw
tri 3698 2064 3792 2158 ne
tri 3792 2064 3886 2158 sw
tri 3792 2036 3820 2064 ne
tri 2651 1892 2745 1986 se
tri 2745 1892 2839 1986 nw
tri 2560 1801 2651 1892 se
rect 2651 1801 2654 1892
tri 2654 1801 2745 1892 nw
tri 2258 1622 2286 1650 sw
tri 2192 1528 2286 1622 ne
tri 2286 1528 2380 1622 sw
tri 2286 1434 2380 1528 ne
tri 2380 1434 2474 1528 sw
tri 2380 1392 2422 1434 ne
rect 2422 1420 2474 1434
tri 2474 1420 2488 1434 sw
rect 2422 1390 2488 1420
tri 2466 534 2560 628 se
rect 2560 600 2626 1801
tri 2626 1773 2654 1801 nw
tri 2560 534 2626 600 nw
rect 3820 660 3886 2064
tri 3886 660 3907 681 sw
rect 3820 653 3907 660
tri 3820 566 3907 653 ne
tri 3907 566 4001 660 sw
tri 2372 440 2466 534 se
tri 2466 440 2560 534 nw
tri 3907 472 4001 566 ne
tri 4001 472 4095 566 sw
tri 2278 346 2372 440 se
tri 2372 346 2466 440 nw
tri 4001 378 4095 472 ne
tri 4095 378 4189 472 sw
tri 4095 350 4123 378 ne
tri 2245 313 2278 346 se
rect 2278 313 2311 346
rect 2245 -760 2311 313
tri 2311 285 2372 346 nw
rect 4123 313 4189 378
use sky130_fd_io__gpiov2_amux_nand4  sky130_fd_io__gpiov2_amux_nand4_0
timestamp 1676037725
transform 1 0 5688 0 -1 3114
box 52 228 930 1718
use sky130_fd_io__gpiov2_amux_nand4  sky130_fd_io__gpiov2_amux_nand4_1
timestamp 1676037725
transform -1 0 5746 0 -1 3114
box 52 228 930 1718
use sky130_fd_io__gpiov2_amux_nand5  sky130_fd_io__gpiov2_amux_nand5_0
timestamp 1676037725
transform 0 1 4701 1 0 140
box 25 228 1061 1718
use sky130_fd_io__gpiov2_amux_nand5  sky130_fd_io__gpiov2_amux_nand5_1
timestamp 1676037725
transform 0 -1 8349 1 0 140
box 25 228 1061 1718
use sky130_fd_io__hvsbt_nand2  sky130_fd_io__hvsbt_nand2_0
timestamp 1676037725
transform -1 0 2178 0 1 139
box 107 226 460 873
use sky130_fd_io__hvsbt_nand2  sky130_fd_io__hvsbt_nand2_1
timestamp 1676037725
transform 1 0 1996 0 1 139
box 107 226 460 873
use sky130_fd_io__hvsbt_nand2  sky130_fd_io__hvsbt_nand2_2
timestamp 1676037725
transform -1 0 3457 0 1 139
box 107 226 460 873
use sky130_fd_io__hvsbt_nand2  sky130_fd_io__hvsbt_nand2_3
timestamp 1676037725
transform -1 0 2992 0 1 139
box 107 226 460 873
use sky130_fd_io__hvsbt_nor  sky130_fd_io__hvsbt_nor_0
timestamp 1676037725
transform 1 0 3391 0 1 139
box 107 226 460 873
use sky130_fd_io__hvsbt_nor  sky130_fd_io__hvsbt_nor_1
timestamp 1676037725
transform -1 0 4396 0 1 139
box 107 226 460 873
use sky130_fd_io__inv_1  sky130_fd_io__inv_1_0
timestamp 1676037725
transform 1 0 2512 0 1 1356
box -38 -49 326 715
use sky130_fd_io__inv_1  sky130_fd_io__inv_1_1
timestamp 1676037725
transform -1 0 1936 0 1 1356
box -38 -49 326 715
use sky130_fd_io__inv_1  sky130_fd_io__inv_1_2
timestamp 1676037725
transform 1 0 976 0 1 1356
box -38 -49 326 715
use sky130_fd_io__inv_1  sky130_fd_io__inv_1_3
timestamp 1676037725
transform -1 0 3760 0 1 1356
box -38 -49 326 715
use sky130_fd_io__inv_1  sky130_fd_io__inv_1_4
timestamp 1676037725
transform -1 0 4048 0 1 1356
box -38 -49 326 715
use sky130_fd_io__inv_1  sky130_fd_io__inv_1_5
timestamp 1676037725
transform -1 0 3088 0 -1 2688
box -38 -49 326 715
use sky130_fd_io__inv_1  sky130_fd_io__inv_1_6
timestamp 1676037725
transform 1 0 1936 0 1 1356
box -38 -49 326 715
use sky130_fd_io__inv_1  sky130_fd_io__inv_1_7
timestamp 1676037725
transform 1 0 4336 0 -1 2688
box -38 -49 326 715
use sky130_fd_io__inv_1  sky130_fd_io__inv_1_8
timestamp 1676037725
transform 1 0 1264 0 -1 2688
box -38 -49 326 715
use sky130_fd_io__inv_1  sky130_fd_io__inv_1_9
timestamp 1676037725
transform 1 0 2512 0 -1 2688
box -38 -49 326 715
use sky130_fd_io__inv_1  sky130_fd_io__inv_1_10
timestamp 1676037725
transform -1 0 4048 0 -1 2688
box -38 -49 326 715
use sky130_fd_io__inv_1  sky130_fd_io__inv_1_11
timestamp 1676037725
transform -1 0 3760 0 -1 2688
box -38 -49 326 715
use sky130_fd_io__inv_1  sky130_fd_io__inv_1_12
timestamp 1676037725
transform 1 0 688 0 -1 2688
box -38 -49 326 715
use sky130_fd_io__inv_1  sky130_fd_io__inv_1_13
timestamp 1676037725
transform 1 0 400 0 -1 2688
box -38 -49 326 715
use sky130_fd_io__inv_1  sky130_fd_io__inv_1_14
timestamp 1676037725
transform 1 0 3088 0 1 1356
box -38 -49 326 715
use sky130_fd_io__nand2_1  sky130_fd_io__nand2_1_0
timestamp 1676037725
transform 1 0 2224 0 -1 2688
box -38 -49 326 715
use sky130_fd_io__nand2_1  sky130_fd_io__nand2_1_1
timestamp 1676037725
transform 1 0 976 0 -1 2688
box -38 -49 326 715
use sky130_fd_io__nand2_1  sky130_fd_io__nand2_1_2
timestamp 1676037725
transform 1 0 4048 0 -1 2688
box -38 -49 326 715
use sky130_fd_io__nand2_1  sky130_fd_io__nand2_1_3
timestamp 1676037725
transform 1 0 3088 0 -1 2688
box -38 -49 326 715
use sky130_fd_io__nor2_1  sky130_fd_io__nor2_1_0
timestamp 1676037725
transform 1 0 688 0 1 1356
box -38 -49 326 715
use sky130_fd_io__nor2_1  sky130_fd_io__nor2_1_1
timestamp 1676037725
transform 1 0 1360 0 1 1356
box -38 -49 326 715
use sky130_fd_io__nor2_1  sky130_fd_io__nor2_1_2
timestamp 1676037725
transform 1 0 2800 0 1 1356
box -38 -49 326 715
use sky130_fd_io__nor2_1  sky130_fd_io__nor2_1_3
timestamp 1676037725
transform 1 0 2224 0 1 1356
box -38 -49 326 715
use sky130_fd_io__tap_1  sky130_fd_io__tap_1_0
timestamp 1676037725
transform 1 0 1264 0 1 1356
box -38 -49 134 715
use sky130_fd_io__tap_1  sky130_fd_io__tap_1_1
timestamp 1676037725
transform 1 0 3376 0 1 1356
box -38 -49 134 715
use sky130_fd_io__tap_1  sky130_fd_io__tap_1_2
timestamp 1676037725
transform 1 0 3376 0 -1 2688
box -38 -49 134 715
use sky130_fd_io__xor2_1  sky130_fd_io__xor2_1_0
timestamp 1676037725
transform 1 0 1552 0 -1 2688
box 0 0 1 1
<< properties >>
string GDS_END 43960948
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 43893108
<< end >>
