VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wb_buttons_leds
  CLASS BLOCK ;
  FOREIGN wb_buttons_leds ;
  ORIGIN 0.000 0.000 ;
  SIZE 2800.000 BY 1760.000 ;
  PIN buttons
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.510 0.000 58.790 4.000 ;
    END
  END buttons
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2099.530 1756.000 2099.810 1760.000 ;
    END
  END clk
  PIN i_wb_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 39.480 4.000 40.080 ;
    END
  END i_wb_addr[0]
  PIN i_wb_addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 216.280 4.000 216.880 ;
    END
  END i_wb_addr[10]
  PIN i_wb_addr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 233.960 4.000 234.560 ;
    END
  END i_wb_addr[11]
  PIN i_wb_addr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 251.640 4.000 252.240 ;
    END
  END i_wb_addr[12]
  PIN i_wb_addr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 269.320 4.000 269.920 ;
    END
  END i_wb_addr[13]
  PIN i_wb_addr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 287.000 4.000 287.600 ;
    END
  END i_wb_addr[14]
  PIN i_wb_addr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 304.680 4.000 305.280 ;
    END
  END i_wb_addr[15]
  PIN i_wb_addr[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 322.360 4.000 322.960 ;
    END
  END i_wb_addr[16]
  PIN i_wb_addr[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 340.040 4.000 340.640 ;
    END
  END i_wb_addr[17]
  PIN i_wb_addr[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 357.720 4.000 358.320 ;
    END
  END i_wb_addr[18]
  PIN i_wb_addr[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 375.400 4.000 376.000 ;
    END
  END i_wb_addr[19]
  PIN i_wb_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.160 4.000 57.760 ;
    END
  END i_wb_addr[1]
  PIN i_wb_addr[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 393.080 4.000 393.680 ;
    END
  END i_wb_addr[20]
  PIN i_wb_addr[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 410.760 4.000 411.360 ;
    END
  END i_wb_addr[21]
  PIN i_wb_addr[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 428.440 4.000 429.040 ;
    END
  END i_wb_addr[22]
  PIN i_wb_addr[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 446.120 4.000 446.720 ;
    END
  END i_wb_addr[23]
  PIN i_wb_addr[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 463.800 4.000 464.400 ;
    END
  END i_wb_addr[24]
  PIN i_wb_addr[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 481.480 4.000 482.080 ;
    END
  END i_wb_addr[25]
  PIN i_wb_addr[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 499.160 4.000 499.760 ;
    END
  END i_wb_addr[26]
  PIN i_wb_addr[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 516.840 4.000 517.440 ;
    END
  END i_wb_addr[27]
  PIN i_wb_addr[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 534.520 4.000 535.120 ;
    END
  END i_wb_addr[28]
  PIN i_wb_addr[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 552.200 4.000 552.800 ;
    END
  END i_wb_addr[29]
  PIN i_wb_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END i_wb_addr[2]
  PIN i_wb_addr[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 569.880 4.000 570.480 ;
    END
  END i_wb_addr[30]
  PIN i_wb_addr[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 587.560 4.000 588.160 ;
    END
  END i_wb_addr[31]
  PIN i_wb_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 92.520 4.000 93.120 ;
    END
  END i_wb_addr[3]
  PIN i_wb_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.200 4.000 110.800 ;
    END
  END i_wb_addr[4]
  PIN i_wb_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.880 4.000 128.480 ;
    END
  END i_wb_addr[5]
  PIN i_wb_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 145.560 4.000 146.160 ;
    END
  END i_wb_addr[6]
  PIN i_wb_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 4.000 163.840 ;
    END
  END i_wb_addr[7]
  PIN i_wb_addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.920 4.000 181.520 ;
    END
  END i_wb_addr[8]
  PIN i_wb_addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 198.600 4.000 199.200 ;
    END
  END i_wb_addr[9]
  PIN i_wb_cyc
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 176.160 2800.000 176.760 ;
    END
  END i_wb_cyc
  PIN i_wb_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 605.240 4.000 605.840 ;
    END
  END i_wb_data[0]
  PIN i_wb_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 782.040 4.000 782.640 ;
    END
  END i_wb_data[10]
  PIN i_wb_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 799.720 4.000 800.320 ;
    END
  END i_wb_data[11]
  PIN i_wb_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 817.400 4.000 818.000 ;
    END
  END i_wb_data[12]
  PIN i_wb_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 835.080 4.000 835.680 ;
    END
  END i_wb_data[13]
  PIN i_wb_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 852.760 4.000 853.360 ;
    END
  END i_wb_data[14]
  PIN i_wb_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 870.440 4.000 871.040 ;
    END
  END i_wb_data[15]
  PIN i_wb_data[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 888.120 4.000 888.720 ;
    END
  END i_wb_data[16]
  PIN i_wb_data[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 905.800 4.000 906.400 ;
    END
  END i_wb_data[17]
  PIN i_wb_data[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 923.480 4.000 924.080 ;
    END
  END i_wb_data[18]
  PIN i_wb_data[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 941.160 4.000 941.760 ;
    END
  END i_wb_data[19]
  PIN i_wb_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 622.920 4.000 623.520 ;
    END
  END i_wb_data[1]
  PIN i_wb_data[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 958.840 4.000 959.440 ;
    END
  END i_wb_data[20]
  PIN i_wb_data[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 976.520 4.000 977.120 ;
    END
  END i_wb_data[21]
  PIN i_wb_data[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 994.200 4.000 994.800 ;
    END
  END i_wb_data[22]
  PIN i_wb_data[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1011.880 4.000 1012.480 ;
    END
  END i_wb_data[23]
  PIN i_wb_data[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1029.560 4.000 1030.160 ;
    END
  END i_wb_data[24]
  PIN i_wb_data[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1047.240 4.000 1047.840 ;
    END
  END i_wb_data[25]
  PIN i_wb_data[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1064.920 4.000 1065.520 ;
    END
  END i_wb_data[26]
  PIN i_wb_data[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1082.600 4.000 1083.200 ;
    END
  END i_wb_data[27]
  PIN i_wb_data[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1100.280 4.000 1100.880 ;
    END
  END i_wb_data[28]
  PIN i_wb_data[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1117.960 4.000 1118.560 ;
    END
  END i_wb_data[29]
  PIN i_wb_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 640.600 4.000 641.200 ;
    END
  END i_wb_data[2]
  PIN i_wb_data[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1135.640 4.000 1136.240 ;
    END
  END i_wb_data[30]
  PIN i_wb_data[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1153.320 4.000 1153.920 ;
    END
  END i_wb_data[31]
  PIN i_wb_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 658.280 4.000 658.880 ;
    END
  END i_wb_data[3]
  PIN i_wb_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 675.960 4.000 676.560 ;
    END
  END i_wb_data[4]
  PIN i_wb_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 693.640 4.000 694.240 ;
    END
  END i_wb_data[5]
  PIN i_wb_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 711.320 4.000 711.920 ;
    END
  END i_wb_data[6]
  PIN i_wb_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 729.000 4.000 729.600 ;
    END
  END i_wb_data[7]
  PIN i_wb_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 746.680 4.000 747.280 ;
    END
  END i_wb_data[8]
  PIN i_wb_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 764.360 4.000 764.960 ;
    END
  END i_wb_data[9]
  PIN i_wb_stb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 527.720 2800.000 528.320 ;
    END
  END i_wb_stb
  PIN i_wb_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 879.280 2800.000 879.880 ;
    END
  END i_wb_we
  PIN led_enb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.290 0.000 170.570 4.000 ;
    END
  END led_enb[0]
  PIN led_enb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1288.090 0.000 1288.370 4.000 ;
    END
  END led_enb[10]
  PIN led_enb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1399.870 0.000 1400.150 4.000 ;
    END
  END led_enb[11]
  PIN led_enb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.070 0.000 282.350 4.000 ;
    END
  END led_enb[1]
  PIN led_enb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 393.850 0.000 394.130 4.000 ;
    END
  END led_enb[2]
  PIN led_enb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.630 0.000 505.910 4.000 ;
    END
  END led_enb[3]
  PIN led_enb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 617.410 0.000 617.690 4.000 ;
    END
  END led_enb[4]
  PIN led_enb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 729.190 0.000 729.470 4.000 ;
    END
  END led_enb[5]
  PIN led_enb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 840.970 0.000 841.250 4.000 ;
    END
  END led_enb[6]
  PIN led_enb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 952.750 0.000 953.030 4.000 ;
    END
  END led_enb[7]
  PIN led_enb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1064.530 0.000 1064.810 4.000 ;
    END
  END led_enb[8]
  PIN led_enb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1176.310 0.000 1176.590 4.000 ;
    END
  END led_enb[9]
  PIN leds[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1511.650 0.000 1511.930 4.000 ;
    END
  END leds[0]
  PIN leds[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2629.450 0.000 2629.730 4.000 ;
    END
  END leds[10]
  PIN leds[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2741.230 0.000 2741.510 4.000 ;
    END
  END leds[11]
  PIN leds[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1623.430 0.000 1623.710 4.000 ;
    END
  END leds[1]
  PIN leds[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1735.210 0.000 1735.490 4.000 ;
    END
  END leds[2]
  PIN leds[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1846.990 0.000 1847.270 4.000 ;
    END
  END leds[3]
  PIN leds[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1958.770 0.000 1959.050 4.000 ;
    END
  END leds[4]
  PIN leds[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2070.550 0.000 2070.830 4.000 ;
    END
  END leds[5]
  PIN leds[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2182.330 0.000 2182.610 4.000 ;
    END
  END leds[6]
  PIN leds[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2294.110 0.000 2294.390 4.000 ;
    END
  END leds[7]
  PIN leds[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2405.890 0.000 2406.170 4.000 ;
    END
  END leds[8]
  PIN leds[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2517.670 0.000 2517.950 4.000 ;
    END
  END leds[9]
  PIN o_wb_ack
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1230.840 2800.000 1231.440 ;
    END
  END o_wb_ack
  PIN o_wb_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1171.000 4.000 1171.600 ;
    END
  END o_wb_data[0]
  PIN o_wb_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1347.800 4.000 1348.400 ;
    END
  END o_wb_data[10]
  PIN o_wb_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1365.480 4.000 1366.080 ;
    END
  END o_wb_data[11]
  PIN o_wb_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1383.160 4.000 1383.760 ;
    END
  END o_wb_data[12]
  PIN o_wb_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1400.840 4.000 1401.440 ;
    END
  END o_wb_data[13]
  PIN o_wb_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1418.520 4.000 1419.120 ;
    END
  END o_wb_data[14]
  PIN o_wb_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1436.200 4.000 1436.800 ;
    END
  END o_wb_data[15]
  PIN o_wb_data[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1453.880 4.000 1454.480 ;
    END
  END o_wb_data[16]
  PIN o_wb_data[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1471.560 4.000 1472.160 ;
    END
  END o_wb_data[17]
  PIN o_wb_data[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1489.240 4.000 1489.840 ;
    END
  END o_wb_data[18]
  PIN o_wb_data[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1506.920 4.000 1507.520 ;
    END
  END o_wb_data[19]
  PIN o_wb_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1188.680 4.000 1189.280 ;
    END
  END o_wb_data[1]
  PIN o_wb_data[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1524.600 4.000 1525.200 ;
    END
  END o_wb_data[20]
  PIN o_wb_data[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1542.280 4.000 1542.880 ;
    END
  END o_wb_data[21]
  PIN o_wb_data[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1559.960 4.000 1560.560 ;
    END
  END o_wb_data[22]
  PIN o_wb_data[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1577.640 4.000 1578.240 ;
    END
  END o_wb_data[23]
  PIN o_wb_data[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1595.320 4.000 1595.920 ;
    END
  END o_wb_data[24]
  PIN o_wb_data[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1613.000 4.000 1613.600 ;
    END
  END o_wb_data[25]
  PIN o_wb_data[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1630.680 4.000 1631.280 ;
    END
  END o_wb_data[26]
  PIN o_wb_data[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1648.360 4.000 1648.960 ;
    END
  END o_wb_data[27]
  PIN o_wb_data[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1666.040 4.000 1666.640 ;
    END
  END o_wb_data[28]
  PIN o_wb_data[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1683.720 4.000 1684.320 ;
    END
  END o_wb_data[29]
  PIN o_wb_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1206.360 4.000 1206.960 ;
    END
  END o_wb_data[2]
  PIN o_wb_data[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1701.400 4.000 1702.000 ;
    END
  END o_wb_data[30]
  PIN o_wb_data[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1719.080 4.000 1719.680 ;
    END
  END o_wb_data[31]
  PIN o_wb_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1224.040 4.000 1224.640 ;
    END
  END o_wb_data[3]
  PIN o_wb_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1241.720 4.000 1242.320 ;
    END
  END o_wb_data[4]
  PIN o_wb_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1259.400 4.000 1260.000 ;
    END
  END o_wb_data[5]
  PIN o_wb_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1277.080 4.000 1277.680 ;
    END
  END o_wb_data[6]
  PIN o_wb_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1294.760 4.000 1295.360 ;
    END
  END o_wb_data[7]
  PIN o_wb_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1312.440 4.000 1313.040 ;
    END
  END o_wb_data[8]
  PIN o_wb_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1330.120 4.000 1330.720 ;
    END
  END o_wb_data[9]
  PIN o_wb_stall
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1582.400 2800.000 1583.000 ;
    END
  END o_wb_stall
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 699.750 1756.000 700.030 1760.000 ;
    END
  END reset
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.440 10.640 1405.040 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1557.040 10.640 1558.640 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1710.640 10.640 1712.240 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1864.240 10.640 1865.840 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2017.840 10.640 2019.440 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2171.440 10.640 2173.040 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2325.040 10.640 2326.640 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2478.640 10.640 2480.240 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2632.240 10.640 2633.840 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2785.840 10.640 2787.440 1749.200 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1326.640 10.640 1328.240 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1480.240 10.640 1481.840 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1633.840 10.640 1635.440 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1787.440 10.640 1789.040 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1941.040 10.640 1942.640 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2094.640 10.640 2096.240 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2248.240 10.640 2249.840 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2401.840 10.640 2403.440 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2555.440 10.640 2557.040 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2709.040 10.640 2710.640 1749.200 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 2794.040 1749.045 ;
      LAYER met1 ;
        RECT 4.670 4.460 2795.350 1749.200 ;
      LAYER met2 ;
        RECT 4.690 1755.720 699.470 1756.000 ;
        RECT 700.310 1755.720 2099.250 1756.000 ;
        RECT 2100.090 1755.720 2795.330 1756.000 ;
        RECT 4.690 4.280 2795.330 1755.720 ;
        RECT 4.690 4.000 58.230 4.280 ;
        RECT 59.070 4.000 170.010 4.280 ;
        RECT 170.850 4.000 281.790 4.280 ;
        RECT 282.630 4.000 393.570 4.280 ;
        RECT 394.410 4.000 505.350 4.280 ;
        RECT 506.190 4.000 617.130 4.280 ;
        RECT 617.970 4.000 728.910 4.280 ;
        RECT 729.750 4.000 840.690 4.280 ;
        RECT 841.530 4.000 952.470 4.280 ;
        RECT 953.310 4.000 1064.250 4.280 ;
        RECT 1065.090 4.000 1176.030 4.280 ;
        RECT 1176.870 4.000 1287.810 4.280 ;
        RECT 1288.650 4.000 1399.590 4.280 ;
        RECT 1400.430 4.000 1511.370 4.280 ;
        RECT 1512.210 4.000 1623.150 4.280 ;
        RECT 1623.990 4.000 1734.930 4.280 ;
        RECT 1735.770 4.000 1846.710 4.280 ;
        RECT 1847.550 4.000 1958.490 4.280 ;
        RECT 1959.330 4.000 2070.270 4.280 ;
        RECT 2071.110 4.000 2182.050 4.280 ;
        RECT 2182.890 4.000 2293.830 4.280 ;
        RECT 2294.670 4.000 2405.610 4.280 ;
        RECT 2406.450 4.000 2517.390 4.280 ;
        RECT 2518.230 4.000 2629.170 4.280 ;
        RECT 2630.010 4.000 2740.950 4.280 ;
        RECT 2741.790 4.000 2795.330 4.280 ;
      LAYER met3 ;
        RECT 4.000 1720.080 2796.000 1749.125 ;
        RECT 4.400 1718.680 2796.000 1720.080 ;
        RECT 4.000 1702.400 2796.000 1718.680 ;
        RECT 4.400 1701.000 2796.000 1702.400 ;
        RECT 4.000 1684.720 2796.000 1701.000 ;
        RECT 4.400 1683.320 2796.000 1684.720 ;
        RECT 4.000 1667.040 2796.000 1683.320 ;
        RECT 4.400 1665.640 2796.000 1667.040 ;
        RECT 4.000 1649.360 2796.000 1665.640 ;
        RECT 4.400 1647.960 2796.000 1649.360 ;
        RECT 4.000 1631.680 2796.000 1647.960 ;
        RECT 4.400 1630.280 2796.000 1631.680 ;
        RECT 4.000 1614.000 2796.000 1630.280 ;
        RECT 4.400 1612.600 2796.000 1614.000 ;
        RECT 4.000 1596.320 2796.000 1612.600 ;
        RECT 4.400 1594.920 2796.000 1596.320 ;
        RECT 4.000 1583.400 2796.000 1594.920 ;
        RECT 4.000 1582.000 2795.600 1583.400 ;
        RECT 4.000 1578.640 2796.000 1582.000 ;
        RECT 4.400 1577.240 2796.000 1578.640 ;
        RECT 4.000 1560.960 2796.000 1577.240 ;
        RECT 4.400 1559.560 2796.000 1560.960 ;
        RECT 4.000 1543.280 2796.000 1559.560 ;
        RECT 4.400 1541.880 2796.000 1543.280 ;
        RECT 4.000 1525.600 2796.000 1541.880 ;
        RECT 4.400 1524.200 2796.000 1525.600 ;
        RECT 4.000 1507.920 2796.000 1524.200 ;
        RECT 4.400 1506.520 2796.000 1507.920 ;
        RECT 4.000 1490.240 2796.000 1506.520 ;
        RECT 4.400 1488.840 2796.000 1490.240 ;
        RECT 4.000 1472.560 2796.000 1488.840 ;
        RECT 4.400 1471.160 2796.000 1472.560 ;
        RECT 4.000 1454.880 2796.000 1471.160 ;
        RECT 4.400 1453.480 2796.000 1454.880 ;
        RECT 4.000 1437.200 2796.000 1453.480 ;
        RECT 4.400 1435.800 2796.000 1437.200 ;
        RECT 4.000 1419.520 2796.000 1435.800 ;
        RECT 4.400 1418.120 2796.000 1419.520 ;
        RECT 4.000 1401.840 2796.000 1418.120 ;
        RECT 4.400 1400.440 2796.000 1401.840 ;
        RECT 4.000 1384.160 2796.000 1400.440 ;
        RECT 4.400 1382.760 2796.000 1384.160 ;
        RECT 4.000 1366.480 2796.000 1382.760 ;
        RECT 4.400 1365.080 2796.000 1366.480 ;
        RECT 4.000 1348.800 2796.000 1365.080 ;
        RECT 4.400 1347.400 2796.000 1348.800 ;
        RECT 4.000 1331.120 2796.000 1347.400 ;
        RECT 4.400 1329.720 2796.000 1331.120 ;
        RECT 4.000 1313.440 2796.000 1329.720 ;
        RECT 4.400 1312.040 2796.000 1313.440 ;
        RECT 4.000 1295.760 2796.000 1312.040 ;
        RECT 4.400 1294.360 2796.000 1295.760 ;
        RECT 4.000 1278.080 2796.000 1294.360 ;
        RECT 4.400 1276.680 2796.000 1278.080 ;
        RECT 4.000 1260.400 2796.000 1276.680 ;
        RECT 4.400 1259.000 2796.000 1260.400 ;
        RECT 4.000 1242.720 2796.000 1259.000 ;
        RECT 4.400 1241.320 2796.000 1242.720 ;
        RECT 4.000 1231.840 2796.000 1241.320 ;
        RECT 4.000 1230.440 2795.600 1231.840 ;
        RECT 4.000 1225.040 2796.000 1230.440 ;
        RECT 4.400 1223.640 2796.000 1225.040 ;
        RECT 4.000 1207.360 2796.000 1223.640 ;
        RECT 4.400 1205.960 2796.000 1207.360 ;
        RECT 4.000 1189.680 2796.000 1205.960 ;
        RECT 4.400 1188.280 2796.000 1189.680 ;
        RECT 4.000 1172.000 2796.000 1188.280 ;
        RECT 4.400 1170.600 2796.000 1172.000 ;
        RECT 4.000 1154.320 2796.000 1170.600 ;
        RECT 4.400 1152.920 2796.000 1154.320 ;
        RECT 4.000 1136.640 2796.000 1152.920 ;
        RECT 4.400 1135.240 2796.000 1136.640 ;
        RECT 4.000 1118.960 2796.000 1135.240 ;
        RECT 4.400 1117.560 2796.000 1118.960 ;
        RECT 4.000 1101.280 2796.000 1117.560 ;
        RECT 4.400 1099.880 2796.000 1101.280 ;
        RECT 4.000 1083.600 2796.000 1099.880 ;
        RECT 4.400 1082.200 2796.000 1083.600 ;
        RECT 4.000 1065.920 2796.000 1082.200 ;
        RECT 4.400 1064.520 2796.000 1065.920 ;
        RECT 4.000 1048.240 2796.000 1064.520 ;
        RECT 4.400 1046.840 2796.000 1048.240 ;
        RECT 4.000 1030.560 2796.000 1046.840 ;
        RECT 4.400 1029.160 2796.000 1030.560 ;
        RECT 4.000 1012.880 2796.000 1029.160 ;
        RECT 4.400 1011.480 2796.000 1012.880 ;
        RECT 4.000 995.200 2796.000 1011.480 ;
        RECT 4.400 993.800 2796.000 995.200 ;
        RECT 4.000 977.520 2796.000 993.800 ;
        RECT 4.400 976.120 2796.000 977.520 ;
        RECT 4.000 959.840 2796.000 976.120 ;
        RECT 4.400 958.440 2796.000 959.840 ;
        RECT 4.000 942.160 2796.000 958.440 ;
        RECT 4.400 940.760 2796.000 942.160 ;
        RECT 4.000 924.480 2796.000 940.760 ;
        RECT 4.400 923.080 2796.000 924.480 ;
        RECT 4.000 906.800 2796.000 923.080 ;
        RECT 4.400 905.400 2796.000 906.800 ;
        RECT 4.000 889.120 2796.000 905.400 ;
        RECT 4.400 887.720 2796.000 889.120 ;
        RECT 4.000 880.280 2796.000 887.720 ;
        RECT 4.000 878.880 2795.600 880.280 ;
        RECT 4.000 871.440 2796.000 878.880 ;
        RECT 4.400 870.040 2796.000 871.440 ;
        RECT 4.000 853.760 2796.000 870.040 ;
        RECT 4.400 852.360 2796.000 853.760 ;
        RECT 4.000 836.080 2796.000 852.360 ;
        RECT 4.400 834.680 2796.000 836.080 ;
        RECT 4.000 818.400 2796.000 834.680 ;
        RECT 4.400 817.000 2796.000 818.400 ;
        RECT 4.000 800.720 2796.000 817.000 ;
        RECT 4.400 799.320 2796.000 800.720 ;
        RECT 4.000 783.040 2796.000 799.320 ;
        RECT 4.400 781.640 2796.000 783.040 ;
        RECT 4.000 765.360 2796.000 781.640 ;
        RECT 4.400 763.960 2796.000 765.360 ;
        RECT 4.000 747.680 2796.000 763.960 ;
        RECT 4.400 746.280 2796.000 747.680 ;
        RECT 4.000 730.000 2796.000 746.280 ;
        RECT 4.400 728.600 2796.000 730.000 ;
        RECT 4.000 712.320 2796.000 728.600 ;
        RECT 4.400 710.920 2796.000 712.320 ;
        RECT 4.000 694.640 2796.000 710.920 ;
        RECT 4.400 693.240 2796.000 694.640 ;
        RECT 4.000 676.960 2796.000 693.240 ;
        RECT 4.400 675.560 2796.000 676.960 ;
        RECT 4.000 659.280 2796.000 675.560 ;
        RECT 4.400 657.880 2796.000 659.280 ;
        RECT 4.000 641.600 2796.000 657.880 ;
        RECT 4.400 640.200 2796.000 641.600 ;
        RECT 4.000 623.920 2796.000 640.200 ;
        RECT 4.400 622.520 2796.000 623.920 ;
        RECT 4.000 606.240 2796.000 622.520 ;
        RECT 4.400 604.840 2796.000 606.240 ;
        RECT 4.000 588.560 2796.000 604.840 ;
        RECT 4.400 587.160 2796.000 588.560 ;
        RECT 4.000 570.880 2796.000 587.160 ;
        RECT 4.400 569.480 2796.000 570.880 ;
        RECT 4.000 553.200 2796.000 569.480 ;
        RECT 4.400 551.800 2796.000 553.200 ;
        RECT 4.000 535.520 2796.000 551.800 ;
        RECT 4.400 534.120 2796.000 535.520 ;
        RECT 4.000 528.720 2796.000 534.120 ;
        RECT 4.000 527.320 2795.600 528.720 ;
        RECT 4.000 517.840 2796.000 527.320 ;
        RECT 4.400 516.440 2796.000 517.840 ;
        RECT 4.000 500.160 2796.000 516.440 ;
        RECT 4.400 498.760 2796.000 500.160 ;
        RECT 4.000 482.480 2796.000 498.760 ;
        RECT 4.400 481.080 2796.000 482.480 ;
        RECT 4.000 464.800 2796.000 481.080 ;
        RECT 4.400 463.400 2796.000 464.800 ;
        RECT 4.000 447.120 2796.000 463.400 ;
        RECT 4.400 445.720 2796.000 447.120 ;
        RECT 4.000 429.440 2796.000 445.720 ;
        RECT 4.400 428.040 2796.000 429.440 ;
        RECT 4.000 411.760 2796.000 428.040 ;
        RECT 4.400 410.360 2796.000 411.760 ;
        RECT 4.000 394.080 2796.000 410.360 ;
        RECT 4.400 392.680 2796.000 394.080 ;
        RECT 4.000 376.400 2796.000 392.680 ;
        RECT 4.400 375.000 2796.000 376.400 ;
        RECT 4.000 358.720 2796.000 375.000 ;
        RECT 4.400 357.320 2796.000 358.720 ;
        RECT 4.000 341.040 2796.000 357.320 ;
        RECT 4.400 339.640 2796.000 341.040 ;
        RECT 4.000 323.360 2796.000 339.640 ;
        RECT 4.400 321.960 2796.000 323.360 ;
        RECT 4.000 305.680 2796.000 321.960 ;
        RECT 4.400 304.280 2796.000 305.680 ;
        RECT 4.000 288.000 2796.000 304.280 ;
        RECT 4.400 286.600 2796.000 288.000 ;
        RECT 4.000 270.320 2796.000 286.600 ;
        RECT 4.400 268.920 2796.000 270.320 ;
        RECT 4.000 252.640 2796.000 268.920 ;
        RECT 4.400 251.240 2796.000 252.640 ;
        RECT 4.000 234.960 2796.000 251.240 ;
        RECT 4.400 233.560 2796.000 234.960 ;
        RECT 4.000 217.280 2796.000 233.560 ;
        RECT 4.400 215.880 2796.000 217.280 ;
        RECT 4.000 199.600 2796.000 215.880 ;
        RECT 4.400 198.200 2796.000 199.600 ;
        RECT 4.000 181.920 2796.000 198.200 ;
        RECT 4.400 180.520 2796.000 181.920 ;
        RECT 4.000 177.160 2796.000 180.520 ;
        RECT 4.000 175.760 2795.600 177.160 ;
        RECT 4.000 164.240 2796.000 175.760 ;
        RECT 4.400 162.840 2796.000 164.240 ;
        RECT 4.000 146.560 2796.000 162.840 ;
        RECT 4.400 145.160 2796.000 146.560 ;
        RECT 4.000 128.880 2796.000 145.160 ;
        RECT 4.400 127.480 2796.000 128.880 ;
        RECT 4.000 111.200 2796.000 127.480 ;
        RECT 4.400 109.800 2796.000 111.200 ;
        RECT 4.000 93.520 2796.000 109.800 ;
        RECT 4.400 92.120 2796.000 93.520 ;
        RECT 4.000 75.840 2796.000 92.120 ;
        RECT 4.400 74.440 2796.000 75.840 ;
        RECT 4.000 58.160 2796.000 74.440 ;
        RECT 4.400 56.760 2796.000 58.160 ;
        RECT 4.000 40.480 2796.000 56.760 ;
        RECT 4.400 39.080 2796.000 40.480 ;
        RECT 4.000 10.715 2796.000 39.080 ;
      LAYER met4 ;
        RECT 9.495 872.615 20.640 1314.945 ;
        RECT 23.040 872.615 97.440 1314.945 ;
        RECT 99.840 872.615 174.240 1314.945 ;
        RECT 176.640 872.615 251.040 1314.945 ;
        RECT 253.440 872.615 327.840 1314.945 ;
        RECT 330.240 872.615 404.640 1314.945 ;
        RECT 407.040 872.615 481.440 1314.945 ;
        RECT 483.840 872.615 558.240 1314.945 ;
        RECT 560.640 872.615 635.040 1314.945 ;
        RECT 637.440 872.615 711.840 1314.945 ;
        RECT 714.240 872.615 788.640 1314.945 ;
        RECT 791.040 872.615 842.425 1314.945 ;
  END
END wb_buttons_leds
END LIBRARY

