magic
tech sky130A
magscale 1 2
timestamp 1676037725
<< nwell >>
rect -38 261 1326 582
<< pwell >>
rect 1 21 1239 203
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 177
rect 163 47 193 177
rect 247 47 277 177
rect 331 47 361 177
rect 415 47 445 177
rect 511 47 541 177
rect 607 47 637 177
rect 691 47 721 177
rect 879 47 909 177
rect 963 47 993 177
rect 1047 47 1077 177
rect 1131 47 1161 177
<< scpmoshvt >>
rect 79 297 109 497
rect 163 297 193 497
rect 247 297 277 497
rect 331 297 361 497
rect 415 297 445 497
rect 511 297 541 497
rect 607 297 637 497
rect 691 297 721 497
rect 879 297 909 497
rect 963 297 993 497
rect 1047 297 1077 497
rect 1131 297 1161 497
<< ndiff >>
rect 27 165 79 177
rect 27 131 35 165
rect 69 131 79 165
rect 27 97 79 131
rect 27 63 35 97
rect 69 63 79 97
rect 27 47 79 63
rect 109 47 163 177
rect 193 47 247 177
rect 277 113 331 177
rect 277 79 287 113
rect 321 79 331 113
rect 277 47 331 79
rect 361 47 415 177
rect 445 47 511 177
rect 541 90 607 177
rect 541 56 559 90
rect 593 56 607 90
rect 541 47 607 56
rect 637 161 691 177
rect 637 127 647 161
rect 681 127 691 161
rect 637 93 691 127
rect 637 59 647 93
rect 681 59 691 93
rect 637 47 691 59
rect 721 97 879 177
rect 721 63 747 97
rect 781 63 819 97
rect 853 63 879 97
rect 721 47 879 63
rect 909 165 963 177
rect 909 131 919 165
rect 953 131 963 165
rect 909 47 963 131
rect 993 97 1047 177
rect 993 63 1003 97
rect 1037 63 1047 97
rect 993 47 1047 63
rect 1077 165 1131 177
rect 1077 131 1087 165
rect 1121 131 1131 165
rect 1077 47 1131 131
rect 1161 97 1213 177
rect 1161 63 1171 97
rect 1205 63 1213 97
rect 1161 47 1213 63
<< pdiff >>
rect 27 477 79 497
rect 27 443 35 477
rect 69 443 79 477
rect 27 407 79 443
rect 27 373 35 407
rect 69 373 79 407
rect 27 297 79 373
rect 109 459 163 497
rect 109 425 119 459
rect 153 425 163 459
rect 109 297 163 425
rect 193 477 247 497
rect 193 443 203 477
rect 237 443 247 477
rect 193 407 247 443
rect 193 373 203 407
rect 237 373 247 407
rect 193 297 247 373
rect 277 459 331 497
rect 277 425 287 459
rect 321 425 331 459
rect 277 297 331 425
rect 361 477 415 497
rect 361 443 371 477
rect 405 443 415 477
rect 361 407 415 443
rect 361 373 371 407
rect 405 373 415 407
rect 361 297 415 373
rect 445 459 511 497
rect 445 425 455 459
rect 489 425 511 459
rect 445 297 511 425
rect 541 477 607 497
rect 541 443 563 477
rect 597 443 607 477
rect 541 407 607 443
rect 541 373 563 407
rect 597 373 607 407
rect 541 297 607 373
rect 637 423 691 497
rect 637 389 647 423
rect 681 389 691 423
rect 637 343 691 389
rect 637 309 647 343
rect 681 309 691 343
rect 637 297 691 309
rect 721 477 773 497
rect 721 443 731 477
rect 765 443 773 477
rect 721 409 773 443
rect 721 375 731 409
rect 765 375 773 409
rect 721 297 773 375
rect 827 459 879 497
rect 827 425 835 459
rect 869 425 879 459
rect 827 297 879 425
rect 909 477 963 497
rect 909 443 919 477
rect 953 443 963 477
rect 909 407 963 443
rect 909 373 919 407
rect 953 373 963 407
rect 909 297 963 373
rect 993 459 1047 497
rect 993 425 1003 459
rect 1037 425 1047 459
rect 993 297 1047 425
rect 1077 477 1131 497
rect 1077 443 1087 477
rect 1121 443 1131 477
rect 1077 407 1131 443
rect 1077 373 1087 407
rect 1121 373 1131 407
rect 1077 297 1131 373
rect 1161 459 1261 497
rect 1161 425 1171 459
rect 1205 425 1261 459
rect 1161 297 1261 425
<< ndiffc >>
rect 35 131 69 165
rect 35 63 69 97
rect 287 79 321 113
rect 559 56 593 90
rect 647 127 681 161
rect 647 59 681 93
rect 747 63 781 97
rect 819 63 853 97
rect 919 131 953 165
rect 1003 63 1037 97
rect 1087 131 1121 165
rect 1171 63 1205 97
<< pdiffc >>
rect 35 443 69 477
rect 35 373 69 407
rect 119 425 153 459
rect 203 443 237 477
rect 203 373 237 407
rect 287 425 321 459
rect 371 443 405 477
rect 371 373 405 407
rect 455 425 489 459
rect 563 443 597 477
rect 563 373 597 407
rect 647 389 681 423
rect 647 309 681 343
rect 731 443 765 477
rect 731 375 765 409
rect 835 425 869 459
rect 919 443 953 477
rect 919 373 953 407
rect 1003 425 1037 459
rect 1087 443 1121 477
rect 1087 373 1121 407
rect 1171 425 1205 459
<< poly >>
rect 79 497 109 523
rect 163 497 193 523
rect 247 497 277 523
rect 331 497 361 523
rect 415 497 445 523
rect 511 497 541 523
rect 607 497 637 523
rect 691 497 721 523
rect 879 497 909 523
rect 963 497 993 523
rect 1047 497 1077 523
rect 1131 497 1161 523
rect 79 265 109 297
rect 163 265 193 297
rect 45 249 109 265
rect 45 215 55 249
rect 89 215 109 249
rect 45 199 109 215
rect 151 249 205 265
rect 151 215 161 249
rect 195 215 205 249
rect 151 199 205 215
rect 247 259 277 297
rect 331 259 361 297
rect 415 265 445 297
rect 511 265 541 297
rect 607 265 637 297
rect 691 265 721 297
rect 879 265 909 297
rect 963 265 993 297
rect 1047 265 1077 297
rect 1131 265 1161 297
rect 247 249 361 259
rect 247 215 287 249
rect 321 215 361 249
rect 247 205 361 215
rect 79 177 109 199
rect 163 177 193 199
rect 247 177 277 205
rect 331 177 361 205
rect 403 249 457 265
rect 403 215 413 249
rect 447 215 457 249
rect 403 199 457 215
rect 511 249 565 265
rect 511 215 521 249
rect 555 215 565 249
rect 511 199 565 215
rect 607 259 721 265
rect 607 249 781 259
rect 607 215 731 249
rect 765 215 781 249
rect 607 205 781 215
rect 871 249 1197 265
rect 871 215 881 249
rect 915 215 949 249
rect 983 215 1017 249
rect 1051 215 1085 249
rect 1119 215 1153 249
rect 1187 215 1197 249
rect 607 199 721 205
rect 871 199 1197 215
rect 415 177 445 199
rect 511 177 541 199
rect 607 177 637 199
rect 691 177 721 199
rect 879 177 909 199
rect 963 177 993 199
rect 1047 177 1077 199
rect 1131 177 1161 199
rect 79 21 109 47
rect 163 21 193 47
rect 247 21 277 47
rect 331 21 361 47
rect 415 21 445 47
rect 511 21 541 47
rect 607 21 637 47
rect 691 21 721 47
rect 879 21 909 47
rect 963 21 993 47
rect 1047 21 1077 47
rect 1131 21 1161 47
<< polycont >>
rect 55 215 89 249
rect 161 215 195 249
rect 287 215 321 249
rect 413 215 447 249
rect 521 215 555 249
rect 731 215 765 249
rect 881 215 915 249
rect 949 215 983 249
rect 1017 215 1051 249
rect 1085 215 1119 249
rect 1153 215 1187 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 35 477 69 493
rect 35 407 69 443
rect 103 459 169 527
rect 103 425 119 459
rect 153 425 169 459
rect 203 477 237 493
rect 203 407 237 443
rect 271 459 337 527
rect 271 425 287 459
rect 321 425 337 459
rect 371 477 405 493
rect 69 373 203 391
rect 371 407 405 443
rect 439 459 505 527
rect 439 425 455 459
rect 489 425 505 459
rect 563 477 765 493
rect 597 459 731 477
rect 237 373 371 391
rect 563 407 597 443
rect 405 373 563 391
rect 35 357 597 373
rect 631 389 647 423
rect 681 389 697 423
rect 631 343 697 389
rect 731 409 765 443
rect 819 459 885 527
rect 819 425 835 459
rect 869 425 885 459
rect 919 477 953 493
rect 919 407 953 443
rect 987 459 1053 527
rect 987 425 1003 459
rect 1037 425 1053 459
rect 1087 477 1121 493
rect 731 359 765 375
rect 907 373 919 391
rect 1087 407 1121 443
rect 1155 459 1221 527
rect 1155 425 1171 459
rect 1205 425 1221 459
rect 953 373 1087 391
rect 1121 373 1259 391
rect 907 357 1259 373
rect 30 289 571 323
rect 30 249 105 289
rect 271 249 341 255
rect 30 215 55 249
rect 89 215 105 249
rect 145 215 161 249
rect 195 215 211 249
rect 271 215 287 249
rect 321 215 341 249
rect 397 249 463 255
rect 397 215 413 249
rect 447 215 463 249
rect 505 249 571 289
rect 505 215 521 249
rect 555 215 571 249
rect 631 309 647 343
rect 681 325 697 343
rect 681 309 879 325
rect 631 291 879 309
rect 161 181 195 215
rect 397 181 434 215
rect 35 165 69 181
rect 161 147 434 181
rect 631 174 669 291
rect 845 265 879 291
rect 715 249 806 257
rect 715 215 731 249
rect 765 215 806 249
rect 470 161 669 174
rect 35 97 69 131
rect 470 140 647 161
rect 470 113 504 140
rect 271 79 287 113
rect 321 79 504 113
rect 631 127 647 140
rect 681 127 697 161
rect 763 149 806 215
rect 845 249 1187 265
rect 845 215 881 249
rect 915 215 949 249
rect 983 215 1017 249
rect 1051 215 1085 249
rect 1119 215 1153 249
rect 845 199 1187 215
rect 1225 165 1259 357
rect 901 131 919 165
rect 953 131 1087 165
rect 1121 131 1259 165
rect 540 90 597 106
rect 35 17 69 63
rect 540 56 559 90
rect 593 56 597 90
rect 631 93 697 127
rect 631 59 647 93
rect 681 59 697 93
rect 747 97 853 113
rect 781 63 819 97
rect 540 17 597 56
rect 747 17 853 63
rect 987 63 1003 97
rect 1037 63 1053 97
rect 987 17 1053 63
rect 1155 63 1171 97
rect 1205 63 1221 97
rect 1155 17 1221 63
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
<< metal1 >>
rect 0 561 1288 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 0 496 1288 527
rect 0 17 1288 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
rect 0 -48 1288 -17
<< labels >>
flabel locali s 766 153 800 187 0 FreeSans 200 0 0 0 B1
port 4 nsew signal input
flabel locali s 398 153 432 187 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 30 289 64 323 0 FreeSans 200 0 0 0 A3
port 3 nsew signal input
flabel locali s 306 221 340 255 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel locali s 30 221 64 255 0 FreeSans 200 0 0 0 A3
port 3 nsew signal input
flabel locali s 766 221 800 255 0 FreeSans 200 0 0 0 B1
port 4 nsew signal input
flabel locali s 1225 221 1259 255 0 FreeSans 200 0 0 0 X
port 9 nsew signal output
flabel locali s 1225 153 1259 187 0 FreeSans 200 0 0 0 X
port 9 nsew signal output
flabel locali s 1225 357 1259 391 0 FreeSans 200 0 0 0 X
port 9 nsew signal output
flabel locali s 398 221 432 255 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 1225 289 1259 323 0 FreeSans 200 0 0 0 X
port 9 nsew signal output
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 a31o_4
rlabel metal1 s 0 -48 1288 48 1 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1288 592 1 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1288 544
string GDS_END 4137538
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 4127676
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 32.200 0.000 
<< end >>
