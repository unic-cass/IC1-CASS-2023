// This is the unpowered netlist.
module egd_top_wrapper (la_data_in_65,
    wb_clk_i,
    la_data_in_58_43,
    la_data_in_60_59,
    la_data_out_23_16,
    la_data_out_26_24,
    la_data_out_30_27);
 input la_data_in_65;
 input wb_clk_i;
 input [15:0] la_data_in_58_43;
 input [1:0] la_data_in_60_59;
 output [7:0] la_data_out_23_16;
 output [2:0] la_data_out_26_24;
 output [3:0] la_data_out_30_27;

 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire clknet_0__2882_;
 wire clknet_0__2883_;
 wire clknet_0__2884_;
 wire clknet_0__2885_;
 wire clknet_0__2886_;
 wire clknet_0__2887_;
 wire clknet_0__2888_;
 wire clknet_0__2889_;
 wire clknet_0__2890_;
 wire clknet_0__2891_;
 wire clknet_0__2892_;
 wire clknet_0__2893_;
 wire clknet_0__2894_;
 wire clknet_0__2895_;
 wire clknet_0__2896_;
 wire clknet_0__2897_;
 wire clknet_0__2898_;
 wire clknet_0__2899_;
 wire clknet_1_0__leaf__2882_;
 wire clknet_1_0__leaf__2883_;
 wire clknet_1_0__leaf__2884_;
 wire clknet_1_0__leaf__2885_;
 wire clknet_1_0__leaf__2886_;
 wire clknet_1_0__leaf__2887_;
 wire clknet_1_0__leaf__2888_;
 wire clknet_1_0__leaf__2889_;
 wire clknet_1_0__leaf__2890_;
 wire clknet_1_0__leaf__2891_;
 wire clknet_1_0__leaf__2892_;
 wire clknet_1_0__leaf__2893_;
 wire clknet_1_0__leaf__2894_;
 wire clknet_1_0__leaf__2895_;
 wire clknet_1_0__leaf__2896_;
 wire clknet_1_0__leaf__2897_;
 wire clknet_1_0__leaf__2898_;
 wire clknet_1_0__leaf__2899_;
 wire clknet_1_1__leaf__2882_;
 wire clknet_1_1__leaf__2883_;
 wire clknet_1_1__leaf__2884_;
 wire clknet_1_1__leaf__2885_;
 wire clknet_1_1__leaf__2886_;
 wire clknet_1_1__leaf__2887_;
 wire clknet_1_1__leaf__2888_;
 wire clknet_1_1__leaf__2889_;
 wire clknet_1_1__leaf__2890_;
 wire clknet_1_1__leaf__2891_;
 wire clknet_1_1__leaf__2892_;
 wire clknet_1_1__leaf__2893_;
 wire clknet_1_1__leaf__2894_;
 wire clknet_1_1__leaf__2895_;
 wire clknet_1_1__leaf__2896_;
 wire clknet_1_1__leaf__2897_;
 wire clknet_1_1__leaf__2898_;
 wire clknet_1_1__leaf__2899_;
 wire \egd_top.BitStream_buffer.BS_buffer[0] ;
 wire \egd_top.BitStream_buffer.BS_buffer[100] ;
 wire \egd_top.BitStream_buffer.BS_buffer[101] ;
 wire \egd_top.BitStream_buffer.BS_buffer[102] ;
 wire \egd_top.BitStream_buffer.BS_buffer[103] ;
 wire \egd_top.BitStream_buffer.BS_buffer[104] ;
 wire \egd_top.BitStream_buffer.BS_buffer[105] ;
 wire \egd_top.BitStream_buffer.BS_buffer[106] ;
 wire \egd_top.BitStream_buffer.BS_buffer[107] ;
 wire \egd_top.BitStream_buffer.BS_buffer[108] ;
 wire \egd_top.BitStream_buffer.BS_buffer[109] ;
 wire \egd_top.BitStream_buffer.BS_buffer[10] ;
 wire \egd_top.BitStream_buffer.BS_buffer[110] ;
 wire \egd_top.BitStream_buffer.BS_buffer[111] ;
 wire \egd_top.BitStream_buffer.BS_buffer[112] ;
 wire \egd_top.BitStream_buffer.BS_buffer[113] ;
 wire \egd_top.BitStream_buffer.BS_buffer[114] ;
 wire \egd_top.BitStream_buffer.BS_buffer[115] ;
 wire \egd_top.BitStream_buffer.BS_buffer[116] ;
 wire \egd_top.BitStream_buffer.BS_buffer[117] ;
 wire \egd_top.BitStream_buffer.BS_buffer[118] ;
 wire \egd_top.BitStream_buffer.BS_buffer[119] ;
 wire \egd_top.BitStream_buffer.BS_buffer[11] ;
 wire \egd_top.BitStream_buffer.BS_buffer[120] ;
 wire \egd_top.BitStream_buffer.BS_buffer[121] ;
 wire \egd_top.BitStream_buffer.BS_buffer[122] ;
 wire \egd_top.BitStream_buffer.BS_buffer[123] ;
 wire \egd_top.BitStream_buffer.BS_buffer[124] ;
 wire \egd_top.BitStream_buffer.BS_buffer[125] ;
 wire \egd_top.BitStream_buffer.BS_buffer[126] ;
 wire \egd_top.BitStream_buffer.BS_buffer[127] ;
 wire \egd_top.BitStream_buffer.BS_buffer[12] ;
 wire \egd_top.BitStream_buffer.BS_buffer[13] ;
 wire \egd_top.BitStream_buffer.BS_buffer[14] ;
 wire \egd_top.BitStream_buffer.BS_buffer[15] ;
 wire \egd_top.BitStream_buffer.BS_buffer[16] ;
 wire \egd_top.BitStream_buffer.BS_buffer[17] ;
 wire \egd_top.BitStream_buffer.BS_buffer[18] ;
 wire \egd_top.BitStream_buffer.BS_buffer[19] ;
 wire \egd_top.BitStream_buffer.BS_buffer[1] ;
 wire \egd_top.BitStream_buffer.BS_buffer[20] ;
 wire \egd_top.BitStream_buffer.BS_buffer[21] ;
 wire \egd_top.BitStream_buffer.BS_buffer[22] ;
 wire \egd_top.BitStream_buffer.BS_buffer[23] ;
 wire \egd_top.BitStream_buffer.BS_buffer[24] ;
 wire \egd_top.BitStream_buffer.BS_buffer[25] ;
 wire \egd_top.BitStream_buffer.BS_buffer[26] ;
 wire \egd_top.BitStream_buffer.BS_buffer[27] ;
 wire \egd_top.BitStream_buffer.BS_buffer[28] ;
 wire \egd_top.BitStream_buffer.BS_buffer[29] ;
 wire \egd_top.BitStream_buffer.BS_buffer[2] ;
 wire \egd_top.BitStream_buffer.BS_buffer[30] ;
 wire \egd_top.BitStream_buffer.BS_buffer[31] ;
 wire \egd_top.BitStream_buffer.BS_buffer[32] ;
 wire \egd_top.BitStream_buffer.BS_buffer[33] ;
 wire \egd_top.BitStream_buffer.BS_buffer[34] ;
 wire \egd_top.BitStream_buffer.BS_buffer[35] ;
 wire \egd_top.BitStream_buffer.BS_buffer[36] ;
 wire \egd_top.BitStream_buffer.BS_buffer[37] ;
 wire \egd_top.BitStream_buffer.BS_buffer[38] ;
 wire \egd_top.BitStream_buffer.BS_buffer[39] ;
 wire \egd_top.BitStream_buffer.BS_buffer[3] ;
 wire \egd_top.BitStream_buffer.BS_buffer[40] ;
 wire \egd_top.BitStream_buffer.BS_buffer[41] ;
 wire \egd_top.BitStream_buffer.BS_buffer[42] ;
 wire \egd_top.BitStream_buffer.BS_buffer[43] ;
 wire \egd_top.BitStream_buffer.BS_buffer[44] ;
 wire \egd_top.BitStream_buffer.BS_buffer[45] ;
 wire \egd_top.BitStream_buffer.BS_buffer[46] ;
 wire \egd_top.BitStream_buffer.BS_buffer[47] ;
 wire \egd_top.BitStream_buffer.BS_buffer[48] ;
 wire \egd_top.BitStream_buffer.BS_buffer[49] ;
 wire \egd_top.BitStream_buffer.BS_buffer[4] ;
 wire \egd_top.BitStream_buffer.BS_buffer[50] ;
 wire \egd_top.BitStream_buffer.BS_buffer[51] ;
 wire \egd_top.BitStream_buffer.BS_buffer[52] ;
 wire \egd_top.BitStream_buffer.BS_buffer[53] ;
 wire \egd_top.BitStream_buffer.BS_buffer[54] ;
 wire \egd_top.BitStream_buffer.BS_buffer[55] ;
 wire \egd_top.BitStream_buffer.BS_buffer[56] ;
 wire \egd_top.BitStream_buffer.BS_buffer[57] ;
 wire \egd_top.BitStream_buffer.BS_buffer[58] ;
 wire \egd_top.BitStream_buffer.BS_buffer[59] ;
 wire \egd_top.BitStream_buffer.BS_buffer[5] ;
 wire \egd_top.BitStream_buffer.BS_buffer[60] ;
 wire \egd_top.BitStream_buffer.BS_buffer[61] ;
 wire \egd_top.BitStream_buffer.BS_buffer[62] ;
 wire \egd_top.BitStream_buffer.BS_buffer[63] ;
 wire \egd_top.BitStream_buffer.BS_buffer[64] ;
 wire \egd_top.BitStream_buffer.BS_buffer[65] ;
 wire \egd_top.BitStream_buffer.BS_buffer[66] ;
 wire \egd_top.BitStream_buffer.BS_buffer[67] ;
 wire \egd_top.BitStream_buffer.BS_buffer[68] ;
 wire \egd_top.BitStream_buffer.BS_buffer[69] ;
 wire \egd_top.BitStream_buffer.BS_buffer[6] ;
 wire \egd_top.BitStream_buffer.BS_buffer[70] ;
 wire \egd_top.BitStream_buffer.BS_buffer[71] ;
 wire \egd_top.BitStream_buffer.BS_buffer[72] ;
 wire \egd_top.BitStream_buffer.BS_buffer[73] ;
 wire \egd_top.BitStream_buffer.BS_buffer[74] ;
 wire \egd_top.BitStream_buffer.BS_buffer[75] ;
 wire \egd_top.BitStream_buffer.BS_buffer[76] ;
 wire \egd_top.BitStream_buffer.BS_buffer[77] ;
 wire \egd_top.BitStream_buffer.BS_buffer[78] ;
 wire \egd_top.BitStream_buffer.BS_buffer[79] ;
 wire \egd_top.BitStream_buffer.BS_buffer[7] ;
 wire \egd_top.BitStream_buffer.BS_buffer[80] ;
 wire \egd_top.BitStream_buffer.BS_buffer[81] ;
 wire \egd_top.BitStream_buffer.BS_buffer[82] ;
 wire \egd_top.BitStream_buffer.BS_buffer[83] ;
 wire \egd_top.BitStream_buffer.BS_buffer[84] ;
 wire \egd_top.BitStream_buffer.BS_buffer[85] ;
 wire \egd_top.BitStream_buffer.BS_buffer[86] ;
 wire \egd_top.BitStream_buffer.BS_buffer[87] ;
 wire \egd_top.BitStream_buffer.BS_buffer[88] ;
 wire \egd_top.BitStream_buffer.BS_buffer[89] ;
 wire \egd_top.BitStream_buffer.BS_buffer[8] ;
 wire \egd_top.BitStream_buffer.BS_buffer[90] ;
 wire \egd_top.BitStream_buffer.BS_buffer[91] ;
 wire \egd_top.BitStream_buffer.BS_buffer[92] ;
 wire \egd_top.BitStream_buffer.BS_buffer[93] ;
 wire \egd_top.BitStream_buffer.BS_buffer[94] ;
 wire \egd_top.BitStream_buffer.BS_buffer[95] ;
 wire \egd_top.BitStream_buffer.BS_buffer[96] ;
 wire \egd_top.BitStream_buffer.BS_buffer[97] ;
 wire \egd_top.BitStream_buffer.BS_buffer[98] ;
 wire \egd_top.BitStream_buffer.BS_buffer[99] ;
 wire \egd_top.BitStream_buffer.BS_buffer[9] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[10] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[11] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[12] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[13] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[14] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[15] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[1] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[2] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[3] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[4] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[5] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[6] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[7] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[8] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[9] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_valid_n ;
 wire \egd_top.BitStream_buffer.buffer_index[4] ;
 wire \egd_top.BitStream_buffer.buffer_index[5] ;
 wire \egd_top.BitStream_buffer.buffer_index[6] ;
 wire \egd_top.BitStream_buffer.exp_golomb_len[1] ;
 wire \egd_top.BitStream_buffer.exp_golomb_len[2] ;
 wire \egd_top.BitStream_buffer.exp_golomb_len[3] ;
 wire \egd_top.BitStream_buffer.pc[1] ;
 wire \egd_top.BitStream_buffer.pc[2] ;
 wire \egd_top.BitStream_buffer.pc[3] ;
 wire \egd_top.BitStream_buffer.pc[4] ;
 wire \egd_top.BitStream_buffer.pc[5] ;
 wire \egd_top.BitStream_buffer.pc[6] ;
 wire \egd_top.BitStream_buffer.pc_previous[0] ;
 wire \egd_top.BitStream_buffer.pc_previous[1] ;
 wire \egd_top.BitStream_buffer.pc_previous[2] ;
 wire \egd_top.BitStream_buffer.pc_previous[3] ;
 wire \egd_top.BitStream_buffer.pc_previous[4] ;
 wire \egd_top.BitStream_buffer.pc_previous[5] ;
 wire \egd_top.BitStream_buffer.pc_previous[6] ;
 wire \egd_top.exp_golomb_decoding.te_range[2] ;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_0760_));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(_1465_));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(_1494_));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(_1850_));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(_1853_));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(_1891_));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(_1993_));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(_2100_));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(_2130_));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(_2248_));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(_2322_));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_0790_));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(_2966_));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(_2966_));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(_2982_));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(_3001_));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(_3104_));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(_3104_));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(_3243_));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(_3282_));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(_3282_));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_0838_));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(_0669_));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(_1644_));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(_1780_));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(_1857_));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(_2170_));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(_2988_));
 sky130_fd_sc_hd__diode_2 ANTENNA_36 (.DIODE(_3114_));
 sky130_fd_sc_hd__diode_2 ANTENNA_37 (.DIODE(_3283_));
 sky130_fd_sc_hd__diode_2 ANTENNA_38 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_0859_));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(_1056_));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(_1174_));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(_1201_));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(_1302_));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(_1427_));
 sky130_fd_sc_hd__fill_2 FILLER_0_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_314 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_510 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_115 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_326 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_546 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_140 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_17 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_303 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_31 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_448 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_131 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_20 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_392 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_58 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_186 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_28 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_354 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_454 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_476 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_17 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_255 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_310 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_479 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_88 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_424 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_548 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_88 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_301 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_314 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_12 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_170 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_59 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_34 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_366 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_510 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_340 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_142 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_30 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_86 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_423 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_454 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_84 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_22 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_28 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_280 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_438 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_451 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_107 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_20 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_314 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_451 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_546 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_424 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_520 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_12 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_415 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_524 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_22 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_131 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_415 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_224 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_62 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_146 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_471 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_520 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_536 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_314 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_12 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_527 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_228 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_329 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_12 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_496 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_451 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_12 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_135 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_303 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_480 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_546 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_479 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_527 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_78 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_450 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_504 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_538 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_448 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_466 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_56 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_16 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_423 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_546 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_519 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_522 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_534 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_224 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_40 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_451 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_507 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_543 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_104 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_370 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_539 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_130 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_438 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_532 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_357 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_423 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_103 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_163 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_451 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_491 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_507 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_519 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_524 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_539 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_424 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_499 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_18 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_308 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_543 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_547 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_392 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_539 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_478 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_536 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_16 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_28 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_168 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_280 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_12 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_146 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_527 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_539 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_394 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_494 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_478 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_60 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_86 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_114 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_329 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_247 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_76 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_326 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_133 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_224 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_387 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_504 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_538 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_186 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_98 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__and3_1 _3342_ (.A(net33),
    .B(net32),
    .C(net31),
    .X(_2900_));
 sky130_fd_sc_hd__clkbuf_4 _3343_ (.A(net19),
    .X(_2901_));
 sky130_fd_sc_hd__clkbuf_4 _3344_ (.A(_2901_),
    .X(_2902_));
 sky130_fd_sc_hd__o21a_1 _3345_ (.A1(net34),
    .A2(_2900_),
    .B1(_2902_),
    .X(_0321_));
 sky130_fd_sc_hd__inv_2 _3346_ (.A(net34),
    .Y(_2903_));
 sky130_fd_sc_hd__buf_4 _3347_ (.A(net19),
    .X(_2904_));
 sky130_fd_sc_hd__clkinv_2 _3348_ (.A(_2904_),
    .Y(_2905_));
 sky130_fd_sc_hd__inv_2 _3349_ (.A(net31),
    .Y(_2906_));
 sky130_fd_sc_hd__or3b_1 _3350_ (.A(net34),
    .B(_2906_),
    .C_N(net32),
    .X(_2907_));
 sky130_fd_sc_hd__inv_2 _3351_ (.A(net33),
    .Y(_2908_));
 sky130_fd_sc_hd__and2_1 _3352_ (.A(_2907_),
    .B(_2908_),
    .X(_2909_));
 sky130_fd_sc_hd__a211oi_1 _3353_ (.A1(_2903_),
    .A2(_2900_),
    .B1(_2905_),
    .C1(_2909_),
    .Y(_0320_));
 sky130_fd_sc_hd__nor2_1 _3354_ (.A(net33),
    .B(net32),
    .Y(_2910_));
 sky130_fd_sc_hd__nor2_1 _3355_ (.A(_2903_),
    .B(_2910_),
    .Y(_2911_));
 sky130_fd_sc_hd__nor2_1 _3356_ (.A(_2906_),
    .B(_2911_),
    .Y(_2912_));
 sky130_fd_sc_hd__buf_2 _3357_ (.A(_2901_),
    .X(_2913_));
 sky130_fd_sc_hd__o211a_1 _3358_ (.A1(net32),
    .A2(_2912_),
    .B1(_2913_),
    .C1(_2907_),
    .X(_0319_));
 sky130_fd_sc_hd__a21o_1 _3359_ (.A1(_2911_),
    .A2(_2906_),
    .B1(_2905_),
    .X(_2914_));
 sky130_fd_sc_hd__nor2_1 _3360_ (.A(_2912_),
    .B(_2914_),
    .Y(_0318_));
 sky130_fd_sc_hd__nor2_1 _3361_ (.A(net29),
    .B(net28),
    .Y(_2915_));
 sky130_fd_sc_hd__inv_2 _3362_ (.A(net30),
    .Y(_2916_));
 sky130_fd_sc_hd__and2_1 _3363_ (.A(_2915_),
    .B(_2916_),
    .X(_2917_));
 sky130_fd_sc_hd__inv_2 _3364_ (.A(_2917_),
    .Y(_2918_));
 sky130_fd_sc_hd__nand2_1 _3365_ (.A(net30),
    .B(net29),
    .Y(_2919_));
 sky130_fd_sc_hd__nand2_4 _3366_ (.A(\egd_top.BitStream_buffer.pc[2] ),
    .B(\egd_top.BitStream_buffer.pc[3] ),
    .Y(_2920_));
 sky130_fd_sc_hd__inv_2 _3367_ (.A(\egd_top.BitStream_buffer.pc[1] ),
    .Y(_2921_));
 sky130_fd_sc_hd__inv_2 _3368_ (.A(net18),
    .Y(_2922_));
 sky130_fd_sc_hd__clkinv_4 _3369_ (.A(net17),
    .Y(_2923_));
 sky130_fd_sc_hd__nand2_1 _3370_ (.A(_2922_),
    .B(_2923_),
    .Y(_2924_));
 sky130_fd_sc_hd__nand2_4 _3371_ (.A(_2924_),
    .B(\egd_top.BitStream_buffer.pc_previous[0] ),
    .Y(_2925_));
 sky130_fd_sc_hd__nor2_4 _3372_ (.A(net18),
    .B(net17),
    .Y(_2926_));
 sky130_fd_sc_hd__inv_2 _3373_ (.A(\egd_top.BitStream_buffer.pc_previous[0] ),
    .Y(_2927_));
 sky130_fd_sc_hd__nand2_1 _3374_ (.A(_2926_),
    .B(_2927_),
    .Y(_2928_));
 sky130_fd_sc_hd__nand2_4 _3375_ (.A(_2925_),
    .B(_2928_),
    .Y(_2929_));
 sky130_fd_sc_hd__or2_1 _3376_ (.A(_2921_),
    .B(_2929_),
    .X(_2930_));
 sky130_fd_sc_hd__nor2_4 _3377_ (.A(_2920_),
    .B(_2930_),
    .Y(_2931_));
 sky130_fd_sc_hd__clkinv_2 _3378_ (.A(\egd_top.BitStream_buffer.pc[6] ),
    .Y(_2932_));
 sky130_fd_sc_hd__and3_2 _3379_ (.A(_2932_),
    .B(\egd_top.BitStream_buffer.pc[4] ),
    .C(\egd_top.BitStream_buffer.pc[5] ),
    .X(_2933_));
 sky130_fd_sc_hd__buf_4 _3380_ (.A(_2933_),
    .X(_2934_));
 sky130_fd_sc_hd__nand2_4 _3381_ (.A(_2931_),
    .B(_2934_),
    .Y(_2935_));
 sky130_fd_sc_hd__inv_2 _3382_ (.A(_2935_),
    .Y(_2936_));
 sky130_fd_sc_hd__nor2_1 _3383_ (.A(\egd_top.BitStream_buffer.pc[6] ),
    .B(_2936_),
    .Y(_2937_));
 sky130_fd_sc_hd__inv_2 _3384_ (.A(\egd_top.BitStream_buffer.buffer_index[5] ),
    .Y(_2938_));
 sky130_fd_sc_hd__inv_2 _3385_ (.A(\egd_top.BitStream_buffer.buffer_index[4] ),
    .Y(_2939_));
 sky130_fd_sc_hd__and3_1 _3386_ (.A(_2938_),
    .B(_2939_),
    .C(\egd_top.BitStream_buffer.buffer_index[6] ),
    .X(_2940_));
 sky130_fd_sc_hd__and4_1 _3387_ (.A(\egd_top.BitStream_buffer.pc_previous[0] ),
    .B(\egd_top.BitStream_buffer.pc_previous[1] ),
    .C(\egd_top.BitStream_buffer.pc_previous[2] ),
    .D(\egd_top.BitStream_buffer.pc_previous[3] ),
    .X(_2941_));
 sky130_fd_sc_hd__a31o_1 _3388_ (.A1(_2941_),
    .A2(\egd_top.BitStream_buffer.pc_previous[4] ),
    .A3(\egd_top.BitStream_buffer.pc_previous[5] ),
    .B1(\egd_top.BitStream_buffer.pc_previous[6] ),
    .X(_2942_));
 sky130_fd_sc_hd__or3b_1 _3389_ (.A(\egd_top.BitStream_buffer.pc[6] ),
    .B(_2936_),
    .C_N(_2942_),
    .X(_2943_));
 sky130_fd_sc_hd__or3_1 _3390_ (.A(\egd_top.BitStream_buffer.buffer_index[6] ),
    .B(\egd_top.BitStream_buffer.buffer_index[5] ),
    .C(\egd_top.BitStream_buffer.buffer_index[4] ),
    .X(_2944_));
 sky130_fd_sc_hd__a21o_1 _3391_ (.A1(_2944_),
    .A2(\egd_top.BitStream_buffer.pc_previous[6] ),
    .B1(_2932_),
    .X(_2945_));
 sky130_fd_sc_hd__a21oi_1 _3392_ (.A1(_2943_),
    .A2(_2945_),
    .B1(_2918_),
    .Y(_2946_));
 sky130_fd_sc_hd__a31o_1 _3393_ (.A1(_2917_),
    .A2(_2937_),
    .A3(_2940_),
    .B1(_2946_),
    .X(_2947_));
 sky130_fd_sc_hd__a21o_1 _3394_ (.A1(_2918_),
    .A2(_2919_),
    .B1(_2947_),
    .X(_2948_));
 sky130_fd_sc_hd__and4_1 _3395_ (.A(_2908_),
    .B(_2906_),
    .C(net34),
    .D(net32),
    .X(_2949_));
 sky130_fd_sc_hd__nand2_1 _3396_ (.A(_2948_),
    .B(_2949_),
    .Y(_2950_));
 sky130_fd_sc_hd__clkinv_2 _3397_ (.A(_2950_),
    .Y(_2951_));
 sky130_fd_sc_hd__nor2_1 _3398_ (.A(net30),
    .B(net28),
    .Y(_2952_));
 sky130_fd_sc_hd__nor2_1 _3399_ (.A(_2916_),
    .B(_2915_),
    .Y(_2953_));
 sky130_fd_sc_hd__nor2_1 _3400_ (.A(net30),
    .B(net29),
    .Y(_2954_));
 sky130_fd_sc_hd__o31ai_1 _3401_ (.A1(_2952_),
    .A2(_2953_),
    .A3(_2954_),
    .B1(_2951_),
    .Y(_2955_));
 sky130_fd_sc_hd__o211ai_2 _3402_ (.A1(net30),
    .A2(_2951_),
    .B1(_2902_),
    .C1(_2955_),
    .Y(_2956_));
 sky130_fd_sc_hd__inv_2 _3403_ (.A(_2956_),
    .Y(_0317_));
 sky130_fd_sc_hd__nand2_1 _3404_ (.A(net29),
    .B(net28),
    .Y(_2957_));
 sky130_fd_sc_hd__nand2_1 _3405_ (.A(_2957_),
    .B(_2916_),
    .Y(_2958_));
 sky130_fd_sc_hd__o21ai_1 _3406_ (.A1(_2915_),
    .A2(_2958_),
    .B1(_2951_),
    .Y(_2959_));
 sky130_fd_sc_hd__o211ai_2 _3407_ (.A1(net29),
    .A2(_2951_),
    .B1(_2902_),
    .C1(_2959_),
    .Y(_2960_));
 sky130_fd_sc_hd__inv_2 _3408_ (.A(_2960_),
    .Y(_0316_));
 sky130_fd_sc_hd__or2b_1 _3409_ (.A(_2954_),
    .B_N(_2919_),
    .X(_2961_));
 sky130_fd_sc_hd__o21ba_1 _3410_ (.A1(net28),
    .A2(_2961_),
    .B1_N(_2947_),
    .X(_2962_));
 sky130_fd_sc_hd__nand2_1 _3411_ (.A(_2951_),
    .B(_2962_),
    .Y(_2963_));
 sky130_fd_sc_hd__o211a_1 _3412_ (.A1(net28),
    .A2(_2951_),
    .B1(_2913_),
    .C1(_2963_),
    .X(_0315_));
 sky130_fd_sc_hd__inv_2 _3413_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_valid_n ),
    .Y(_2964_));
 sky130_fd_sc_hd__clkbuf_4 _3414_ (.A(_2964_),
    .X(_2965_));
 sky130_fd_sc_hd__o21ai_1 _3415_ (.A1(_2965_),
    .A2(_2949_),
    .B1(_2902_),
    .Y(_0314_));
 sky130_fd_sc_hd__buf_4 _3416_ (.A(net7),
    .X(_2966_));
 sky130_fd_sc_hd__inv_2 _3417_ (.A(\egd_top.BitStream_buffer.buffer_index[6] ),
    .Y(_2967_));
 sky130_fd_sc_hd__and2_1 _3418_ (.A(_2910_),
    .B(_2903_),
    .X(_2968_));
 sky130_fd_sc_hd__or2_1 _3419_ (.A(_2911_),
    .B(_2968_),
    .X(_2969_));
 sky130_fd_sc_hd__nand2_2 _3420_ (.A(_2969_),
    .B(_2961_),
    .Y(_2970_));
 sky130_fd_sc_hd__nand2_1 _3421_ (.A(_2970_),
    .B(\egd_top.BitStream_buffer.buffer_index[4] ),
    .Y(_2971_));
 sky130_fd_sc_hd__or2_1 _3422_ (.A(_2938_),
    .B(_2971_),
    .X(_2972_));
 sky130_fd_sc_hd__nor2_1 _3423_ (.A(_2967_),
    .B(_2972_),
    .Y(_2973_));
 sky130_fd_sc_hd__clkinv_2 _3424_ (.A(_2973_),
    .Y(_2974_));
 sky130_fd_sc_hd__buf_2 _3425_ (.A(_2974_),
    .X(_2975_));
 sky130_fd_sc_hd__clkbuf_4 _3426_ (.A(_2974_),
    .X(_2976_));
 sky130_fd_sc_hd__inv_2 _3427_ (.A(\egd_top.BitStream_buffer.BS_buffer[112] ),
    .Y(_2977_));
 sky130_fd_sc_hd__nand2_1 _3428_ (.A(_2976_),
    .B(_2977_),
    .Y(_2978_));
 sky130_fd_sc_hd__o211a_1 _3429_ (.A1(_2966_),
    .A2(_2975_),
    .B1(_2913_),
    .C1(_2978_),
    .X(_0313_));
 sky130_fd_sc_hd__buf_4 _3430_ (.A(net6),
    .X(_2979_));
 sky130_fd_sc_hd__clkinv_2 _3431_ (.A(\egd_top.BitStream_buffer.BS_buffer[113] ),
    .Y(_2980_));
 sky130_fd_sc_hd__nand2_1 _3432_ (.A(_2976_),
    .B(_2980_),
    .Y(_2981_));
 sky130_fd_sc_hd__o211a_1 _3433_ (.A1(_2979_),
    .A2(_2975_),
    .B1(_2913_),
    .C1(_2981_),
    .X(_0312_));
 sky130_fd_sc_hd__buf_4 _3434_ (.A(net5),
    .X(_2982_));
 sky130_fd_sc_hd__clkinv_2 _3435_ (.A(\egd_top.BitStream_buffer.BS_buffer[114] ),
    .Y(_2983_));
 sky130_fd_sc_hd__nand2_1 _3436_ (.A(_2976_),
    .B(_2983_),
    .Y(_2984_));
 sky130_fd_sc_hd__o211a_1 _3437_ (.A1(_2982_),
    .A2(_2975_),
    .B1(_2913_),
    .C1(_2984_),
    .X(_0311_));
 sky130_fd_sc_hd__buf_4 _3438_ (.A(net4),
    .X(_2985_));
 sky130_fd_sc_hd__inv_2 _3439_ (.A(\egd_top.BitStream_buffer.BS_buffer[115] ),
    .Y(_2986_));
 sky130_fd_sc_hd__nand2_1 _3440_ (.A(_2976_),
    .B(_2986_),
    .Y(_2987_));
 sky130_fd_sc_hd__o211a_1 _3441_ (.A1(_2985_),
    .A2(_2975_),
    .B1(_2913_),
    .C1(_2987_),
    .X(_0310_));
 sky130_fd_sc_hd__buf_4 _3442_ (.A(net3),
    .X(_2988_));
 sky130_fd_sc_hd__clkbuf_4 _3443_ (.A(_2974_),
    .X(_2989_));
 sky130_fd_sc_hd__inv_2 _3444_ (.A(\egd_top.BitStream_buffer.BS_buffer[116] ),
    .Y(_2990_));
 sky130_fd_sc_hd__nand2_1 _3445_ (.A(_2989_),
    .B(_2990_),
    .Y(_2991_));
 sky130_fd_sc_hd__o211a_1 _3446_ (.A1(_2988_),
    .A2(_2975_),
    .B1(_2913_),
    .C1(_2991_),
    .X(_0309_));
 sky130_fd_sc_hd__buf_4 _3447_ (.A(net2),
    .X(_2992_));
 sky130_fd_sc_hd__clkinv_2 _3448_ (.A(\egd_top.BitStream_buffer.BS_buffer[117] ),
    .Y(_2993_));
 sky130_fd_sc_hd__nand2_1 _3449_ (.A(_2989_),
    .B(_2993_),
    .Y(_2994_));
 sky130_fd_sc_hd__o211a_1 _3450_ (.A1(_2992_),
    .A2(_2975_),
    .B1(_2913_),
    .C1(_2994_),
    .X(_0308_));
 sky130_fd_sc_hd__buf_4 _3451_ (.A(net16),
    .X(_2995_));
 sky130_fd_sc_hd__inv_2 _3452_ (.A(\egd_top.BitStream_buffer.BS_buffer[118] ),
    .Y(_2996_));
 sky130_fd_sc_hd__nand2_1 _3453_ (.A(_2989_),
    .B(_2996_),
    .Y(_2997_));
 sky130_fd_sc_hd__o211a_1 _3454_ (.A1(_2995_),
    .A2(_2975_),
    .B1(_2913_),
    .C1(_2997_),
    .X(_0307_));
 sky130_fd_sc_hd__buf_4 _3455_ (.A(net15),
    .X(_2998_));
 sky130_fd_sc_hd__clkinv_2 _3456_ (.A(\egd_top.BitStream_buffer.BS_buffer[119] ),
    .Y(_2999_));
 sky130_fd_sc_hd__nand2_1 _3457_ (.A(_2989_),
    .B(_2999_),
    .Y(_3000_));
 sky130_fd_sc_hd__o211a_1 _3458_ (.A1(_2998_),
    .A2(_2975_),
    .B1(_2913_),
    .C1(_3000_),
    .X(_0306_));
 sky130_fd_sc_hd__buf_4 _3459_ (.A(net14),
    .X(_3001_));
 sky130_fd_sc_hd__clkbuf_4 _3460_ (.A(_2901_),
    .X(_3002_));
 sky130_fd_sc_hd__clkinv_2 _3461_ (.A(\egd_top.BitStream_buffer.BS_buffer[120] ),
    .Y(_3003_));
 sky130_fd_sc_hd__nand2_1 _3462_ (.A(_2989_),
    .B(_3003_),
    .Y(_3004_));
 sky130_fd_sc_hd__o211a_1 _3463_ (.A1(_3001_),
    .A2(_2975_),
    .B1(_3002_),
    .C1(_3004_),
    .X(_0305_));
 sky130_fd_sc_hd__buf_4 _3464_ (.A(net13),
    .X(_3005_));
 sky130_fd_sc_hd__clkinv_2 _3465_ (.A(\egd_top.BitStream_buffer.BS_buffer[121] ),
    .Y(_3006_));
 sky130_fd_sc_hd__nand2_1 _3466_ (.A(_2989_),
    .B(_3006_),
    .Y(_3007_));
 sky130_fd_sc_hd__o211a_1 _3467_ (.A1(_3005_),
    .A2(_2975_),
    .B1(_3002_),
    .C1(_3007_),
    .X(_0304_));
 sky130_fd_sc_hd__clkbuf_4 _3468_ (.A(net12),
    .X(_3008_));
 sky130_fd_sc_hd__clkinv_2 _3469_ (.A(\egd_top.BitStream_buffer.BS_buffer[122] ),
    .Y(_3009_));
 sky130_fd_sc_hd__nand2_1 _3470_ (.A(_2989_),
    .B(_3009_),
    .Y(_3010_));
 sky130_fd_sc_hd__o211a_1 _3471_ (.A1(_3008_),
    .A2(_2976_),
    .B1(_3002_),
    .C1(_3010_),
    .X(_0303_));
 sky130_fd_sc_hd__buf_4 _3472_ (.A(net11),
    .X(_3011_));
 sky130_fd_sc_hd__inv_2 _3473_ (.A(\egd_top.BitStream_buffer.BS_buffer[123] ),
    .Y(_3012_));
 sky130_fd_sc_hd__nand2_1 _3474_ (.A(_2989_),
    .B(_3012_),
    .Y(_3013_));
 sky130_fd_sc_hd__o211a_1 _3475_ (.A1(_3011_),
    .A2(_2976_),
    .B1(_3002_),
    .C1(_3013_),
    .X(_0302_));
 sky130_fd_sc_hd__buf_4 _3476_ (.A(net10),
    .X(_3014_));
 sky130_fd_sc_hd__inv_2 _3477_ (.A(\egd_top.BitStream_buffer.BS_buffer[124] ),
    .Y(_3015_));
 sky130_fd_sc_hd__nand2_1 _3478_ (.A(_2989_),
    .B(_3015_),
    .Y(_3016_));
 sky130_fd_sc_hd__o211a_1 _3479_ (.A1(_3014_),
    .A2(_2976_),
    .B1(_3002_),
    .C1(_3016_),
    .X(_0301_));
 sky130_fd_sc_hd__buf_4 _3480_ (.A(net9),
    .X(_3017_));
 sky130_fd_sc_hd__inv_2 _3481_ (.A(\egd_top.BitStream_buffer.BS_buffer[125] ),
    .Y(_3018_));
 sky130_fd_sc_hd__nand2_1 _3482_ (.A(_2989_),
    .B(_3018_),
    .Y(_3019_));
 sky130_fd_sc_hd__o211a_1 _3483_ (.A1(_3017_),
    .A2(_2976_),
    .B1(_3002_),
    .C1(_3019_),
    .X(_0300_));
 sky130_fd_sc_hd__buf_4 _3484_ (.A(net8),
    .X(_3020_));
 sky130_fd_sc_hd__inv_2 _3485_ (.A(\egd_top.BitStream_buffer.BS_buffer[126] ),
    .Y(_3021_));
 sky130_fd_sc_hd__nand2_1 _3486_ (.A(_2974_),
    .B(_3021_),
    .Y(_3022_));
 sky130_fd_sc_hd__o211a_1 _3487_ (.A1(_3020_),
    .A2(_2976_),
    .B1(_3002_),
    .C1(_3022_),
    .X(_0299_));
 sky130_fd_sc_hd__buf_4 _3488_ (.A(net1),
    .X(_3023_));
 sky130_fd_sc_hd__inv_2 _3489_ (.A(\egd_top.BitStream_buffer.BS_buffer[127] ),
    .Y(_3024_));
 sky130_fd_sc_hd__nand2_1 _3490_ (.A(_2974_),
    .B(_3024_),
    .Y(_3025_));
 sky130_fd_sc_hd__o211a_1 _3491_ (.A1(_3023_),
    .A2(_2976_),
    .B1(_3002_),
    .C1(_3025_),
    .X(_0298_));
 sky130_fd_sc_hd__clkbuf_4 _3492_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_valid_n ),
    .X(_3026_));
 sky130_fd_sc_hd__clkbuf_4 _3493_ (.A(_3026_),
    .X(_3027_));
 sky130_fd_sc_hd__buf_2 _3494_ (.A(\egd_top.BitStream_buffer.BS_buffer[96] ),
    .X(_3028_));
 sky130_fd_sc_hd__nand2_1 _3495_ (.A(_2929_),
    .B(_2921_),
    .Y(_3029_));
 sky130_fd_sc_hd__inv_2 _3496_ (.A(_3029_),
    .Y(_3030_));
 sky130_fd_sc_hd__clkinv_2 _3497_ (.A(\egd_top.BitStream_buffer.pc[2] ),
    .Y(_3031_));
 sky130_fd_sc_hd__clkinv_2 _3498_ (.A(\egd_top.BitStream_buffer.pc[3] ),
    .Y(_3032_));
 sky130_fd_sc_hd__and3_4 _3499_ (.A(_3030_),
    .B(_3031_),
    .C(_3032_),
    .X(_3033_));
 sky130_fd_sc_hd__inv_2 _3500_ (.A(\egd_top.BitStream_buffer.pc[5] ),
    .Y(_3034_));
 sky130_fd_sc_hd__or3_2 _3501_ (.A(\egd_top.BitStream_buffer.pc[4] ),
    .B(_2932_),
    .C(_3034_),
    .X(_3035_));
 sky130_fd_sc_hd__inv_2 _3502_ (.A(_3035_),
    .Y(_3036_));
 sky130_fd_sc_hd__and2_1 _3503_ (.A(_3033_),
    .B(_3036_),
    .X(_3037_));
 sky130_fd_sc_hd__clkbuf_2 _3504_ (.A(_3037_),
    .X(_3038_));
 sky130_fd_sc_hd__clkbuf_4 _3505_ (.A(_3038_),
    .X(_3039_));
 sky130_fd_sc_hd__buf_2 _3506_ (.A(\egd_top.BitStream_buffer.BS_buffer[97] ),
    .X(_3040_));
 sky130_fd_sc_hd__buf_4 _3507_ (.A(_3035_),
    .X(_3041_));
 sky130_fd_sc_hd__or2_1 _3508_ (.A(\egd_top.BitStream_buffer.pc[1] ),
    .B(_2929_),
    .X(_3042_));
 sky130_fd_sc_hd__inv_2 _3509_ (.A(_3042_),
    .Y(_3043_));
 sky130_fd_sc_hd__and3_1 _3510_ (.A(_3043_),
    .B(_3031_),
    .C(_3032_),
    .X(_3044_));
 sky130_fd_sc_hd__buf_6 _3511_ (.A(_3044_),
    .X(_3045_));
 sky130_fd_sc_hd__inv_2 _3512_ (.A(_3045_),
    .Y(_3046_));
 sky130_fd_sc_hd__nor2_2 _3513_ (.A(_3041_),
    .B(_3046_),
    .Y(_3047_));
 sky130_fd_sc_hd__buf_6 _3514_ (.A(_3047_),
    .X(_3048_));
 sky130_fd_sc_hd__clkinv_2 _3515_ (.A(\egd_top.BitStream_buffer.BS_buffer[98] ),
    .Y(_3049_));
 sky130_fd_sc_hd__nand2_1 _3516_ (.A(_2929_),
    .B(\egd_top.BitStream_buffer.pc[1] ),
    .Y(_3050_));
 sky130_fd_sc_hd__inv_2 _3517_ (.A(_3050_),
    .Y(_3051_));
 sky130_fd_sc_hd__and3_2 _3518_ (.A(_3051_),
    .B(_3031_),
    .C(_3032_),
    .X(_3052_));
 sky130_fd_sc_hd__clkinv_2 _3519_ (.A(_3052_),
    .Y(_3053_));
 sky130_fd_sc_hd__nor2_1 _3520_ (.A(_3035_),
    .B(_3053_),
    .Y(_3054_));
 sky130_fd_sc_hd__inv_2 _3521_ (.A(_3054_),
    .Y(_3055_));
 sky130_fd_sc_hd__clkbuf_4 _3522_ (.A(_3055_),
    .X(_3056_));
 sky130_fd_sc_hd__inv_2 _3523_ (.A(_2930_),
    .Y(_3057_));
 sky130_fd_sc_hd__and3_2 _3524_ (.A(_3057_),
    .B(_3031_),
    .C(_3032_),
    .X(_3058_));
 sky130_fd_sc_hd__clkinv_2 _3525_ (.A(_3058_),
    .Y(_3059_));
 sky130_fd_sc_hd__nor2_2 _3526_ (.A(_3041_),
    .B(_3059_),
    .Y(_3060_));
 sky130_fd_sc_hd__buf_6 _3527_ (.A(_3060_),
    .X(_3061_));
 sky130_fd_sc_hd__clkbuf_4 _3528_ (.A(\egd_top.BitStream_buffer.BS_buffer[99] ),
    .X(_3062_));
 sky130_fd_sc_hd__nand2_1 _3529_ (.A(_3061_),
    .B(_3062_),
    .Y(_3063_));
 sky130_fd_sc_hd__o21ai_1 _3530_ (.A1(_3049_),
    .A2(_3056_),
    .B1(_3063_),
    .Y(_3064_));
 sky130_fd_sc_hd__a221oi_1 _3531_ (.A1(_3028_),
    .A2(_3039_),
    .B1(_3040_),
    .B2(_3048_),
    .C1(_3064_),
    .Y(_3065_));
 sky130_fd_sc_hd__clkbuf_4 _3532_ (.A(\egd_top.BitStream_buffer.BS_buffer[108] ),
    .X(_3066_));
 sky130_fd_sc_hd__nor2_4 _3533_ (.A(_2920_),
    .B(_3029_),
    .Y(_3067_));
 sky130_fd_sc_hd__inv_2 _3534_ (.A(_3067_),
    .Y(_3068_));
 sky130_fd_sc_hd__nor2_2 _3535_ (.A(_3035_),
    .B(_3068_),
    .Y(_3069_));
 sky130_fd_sc_hd__clkbuf_4 _3536_ (.A(\egd_top.BitStream_buffer.BS_buffer[109] ),
    .X(_3070_));
 sky130_fd_sc_hd__nor2_4 _3537_ (.A(_2920_),
    .B(_3042_),
    .Y(_3071_));
 sky130_fd_sc_hd__clkinv_2 _3538_ (.A(_3071_),
    .Y(_3072_));
 sky130_fd_sc_hd__nor2_2 _3539_ (.A(_3041_),
    .B(_3072_),
    .Y(_3073_));
 sky130_fd_sc_hd__buf_4 _3540_ (.A(_3073_),
    .X(_3074_));
 sky130_fd_sc_hd__clkbuf_4 _3541_ (.A(\egd_top.BitStream_buffer.BS_buffer[110] ),
    .X(_3075_));
 sky130_fd_sc_hd__nor2_2 _3542_ (.A(_2920_),
    .B(_3050_),
    .Y(_3076_));
 sky130_fd_sc_hd__inv_2 _3543_ (.A(_3076_),
    .Y(_3077_));
 sky130_fd_sc_hd__nor2_2 _3544_ (.A(_3041_),
    .B(_3077_),
    .Y(_3078_));
 sky130_fd_sc_hd__clkinv_2 _3545_ (.A(_2931_),
    .Y(_3079_));
 sky130_fd_sc_hd__nor2_2 _3546_ (.A(_3041_),
    .B(_3079_),
    .Y(_3080_));
 sky130_fd_sc_hd__buf_4 _3547_ (.A(_3080_),
    .X(_3081_));
 sky130_fd_sc_hd__clkbuf_4 _3548_ (.A(\egd_top.BitStream_buffer.BS_buffer[111] ),
    .X(_3082_));
 sky130_fd_sc_hd__a22o_1 _3549_ (.A1(_3075_),
    .A2(_3078_),
    .B1(_3081_),
    .B2(_3082_),
    .X(_3083_));
 sky130_fd_sc_hd__a221oi_1 _3550_ (.A1(_3066_),
    .A2(_3069_),
    .B1(_3070_),
    .B2(_3074_),
    .C1(_3083_),
    .Y(_3084_));
 sky130_fd_sc_hd__clkinv_2 _3551_ (.A(\egd_top.BitStream_buffer.BS_buffer[103] ),
    .Y(_3085_));
 sky130_fd_sc_hd__and3_1 _3552_ (.A(_3057_),
    .B(\egd_top.BitStream_buffer.pc[2] ),
    .C(_3032_),
    .X(_3086_));
 sky130_fd_sc_hd__buf_6 _3553_ (.A(_3086_),
    .X(_3087_));
 sky130_fd_sc_hd__nand2_2 _3554_ (.A(_3087_),
    .B(_3036_),
    .Y(_3088_));
 sky130_fd_sc_hd__clkbuf_4 _3555_ (.A(_3088_),
    .X(_3089_));
 sky130_fd_sc_hd__and3_2 _3556_ (.A(_3030_),
    .B(\egd_top.BitStream_buffer.pc[2] ),
    .C(_3032_),
    .X(_3090_));
 sky130_fd_sc_hd__inv_2 _3557_ (.A(_3090_),
    .Y(_3091_));
 sky130_fd_sc_hd__nor2_2 _3558_ (.A(_3041_),
    .B(_3091_),
    .Y(_3092_));
 sky130_fd_sc_hd__buf_4 _3559_ (.A(_3092_),
    .X(_3093_));
 sky130_fd_sc_hd__clkbuf_4 _3560_ (.A(\egd_top.BitStream_buffer.BS_buffer[100] ),
    .X(_3094_));
 sky130_fd_sc_hd__nand2_1 _3561_ (.A(_3093_),
    .B(_3094_),
    .Y(_3095_));
 sky130_fd_sc_hd__and3_2 _3562_ (.A(_3051_),
    .B(\egd_top.BitStream_buffer.pc[2] ),
    .C(_3032_),
    .X(_3096_));
 sky130_fd_sc_hd__inv_2 _3563_ (.A(_3096_),
    .Y(_3097_));
 sky130_fd_sc_hd__nor2_2 _3564_ (.A(_3041_),
    .B(_3097_),
    .Y(_3098_));
 sky130_fd_sc_hd__buf_4 _3565_ (.A(_3098_),
    .X(_3099_));
 sky130_fd_sc_hd__buf_2 _3566_ (.A(\egd_top.BitStream_buffer.BS_buffer[102] ),
    .X(_3100_));
 sky130_fd_sc_hd__nand2_1 _3567_ (.A(_3099_),
    .B(_3100_),
    .Y(_3101_));
 sky130_fd_sc_hd__inv_2 _3568_ (.A(\egd_top.BitStream_buffer.BS_buffer[101] ),
    .Y(_3102_));
 sky130_fd_sc_hd__and3_1 _3569_ (.A(_3043_),
    .B(\egd_top.BitStream_buffer.pc[2] ),
    .C(_3032_),
    .X(_3103_));
 sky130_fd_sc_hd__buf_6 _3570_ (.A(_3103_),
    .X(_3104_));
 sky130_fd_sc_hd__nand2_1 _3571_ (.A(_3104_),
    .B(_3036_),
    .Y(_3105_));
 sky130_fd_sc_hd__buf_2 _3572_ (.A(_3105_),
    .X(_3106_));
 sky130_fd_sc_hd__or2_1 _3573_ (.A(_3102_),
    .B(_3106_),
    .X(_3107_));
 sky130_fd_sc_hd__o2111a_1 _3574_ (.A1(_3085_),
    .A2(_3089_),
    .B1(_3095_),
    .C1(_3101_),
    .D1(_3107_),
    .X(_3108_));
 sky130_fd_sc_hd__clkbuf_4 _3575_ (.A(\egd_top.BitStream_buffer.BS_buffer[106] ),
    .X(_3109_));
 sky130_fd_sc_hd__and3_2 _3576_ (.A(_3051_),
    .B(_3031_),
    .C(\egd_top.BitStream_buffer.pc[3] ),
    .X(_3110_));
 sky130_fd_sc_hd__clkinv_2 _3577_ (.A(_3110_),
    .Y(_3111_));
 sky130_fd_sc_hd__nor2_2 _3578_ (.A(_3041_),
    .B(_3111_),
    .Y(_3112_));
 sky130_fd_sc_hd__buf_2 _3579_ (.A(_3112_),
    .X(_3113_));
 sky130_fd_sc_hd__and3_4 _3580_ (.A(_3057_),
    .B(_3031_),
    .C(\egd_top.BitStream_buffer.pc[3] ),
    .X(_3114_));
 sky130_fd_sc_hd__inv_2 _3581_ (.A(_3114_),
    .Y(_3115_));
 sky130_fd_sc_hd__nor2_2 _3582_ (.A(_3041_),
    .B(_3115_),
    .Y(_3116_));
 sky130_fd_sc_hd__buf_2 _3583_ (.A(_3116_),
    .X(_3117_));
 sky130_fd_sc_hd__clkbuf_4 _3584_ (.A(\egd_top.BitStream_buffer.BS_buffer[107] ),
    .X(_3118_));
 sky130_fd_sc_hd__clkinv_2 _3585_ (.A(\egd_top.BitStream_buffer.BS_buffer[105] ),
    .Y(_3119_));
 sky130_fd_sc_hd__and3_1 _3586_ (.A(_3043_),
    .B(_3031_),
    .C(\egd_top.BitStream_buffer.pc[3] ),
    .X(_3120_));
 sky130_fd_sc_hd__buf_6 _3587_ (.A(_3120_),
    .X(_3121_));
 sky130_fd_sc_hd__nand2_2 _3588_ (.A(_3121_),
    .B(_3036_),
    .Y(_3122_));
 sky130_fd_sc_hd__buf_2 _3589_ (.A(_3122_),
    .X(_3123_));
 sky130_fd_sc_hd__and3_2 _3590_ (.A(_3030_),
    .B(_3031_),
    .C(\egd_top.BitStream_buffer.pc[3] ),
    .X(_3124_));
 sky130_fd_sc_hd__inv_2 _3591_ (.A(_3124_),
    .Y(_3125_));
 sky130_fd_sc_hd__nor2_2 _3592_ (.A(_3041_),
    .B(_3125_),
    .Y(_3126_));
 sky130_fd_sc_hd__buf_2 _3593_ (.A(_3126_),
    .X(_3127_));
 sky130_fd_sc_hd__clkbuf_4 _3594_ (.A(\egd_top.BitStream_buffer.BS_buffer[104] ),
    .X(_3128_));
 sky130_fd_sc_hd__nand2_1 _3595_ (.A(_3127_),
    .B(_3128_),
    .Y(_3129_));
 sky130_fd_sc_hd__o21ai_1 _3596_ (.A1(_3119_),
    .A2(_3123_),
    .B1(_3129_),
    .Y(_3130_));
 sky130_fd_sc_hd__a221oi_1 _3597_ (.A1(_3109_),
    .A2(_3113_),
    .B1(_3117_),
    .B2(_3118_),
    .C1(_3130_),
    .Y(_3131_));
 sky130_fd_sc_hd__and4_1 _3598_ (.A(_3065_),
    .B(_3084_),
    .C(_3108_),
    .D(_3131_),
    .X(_3132_));
 sky130_fd_sc_hd__clkbuf_4 _3599_ (.A(\egd_top.BitStream_buffer.BS_buffer[122] ),
    .X(_3133_));
 sky130_fd_sc_hd__and3_2 _3600_ (.A(\egd_top.BitStream_buffer.pc[6] ),
    .B(\egd_top.BitStream_buffer.pc[4] ),
    .C(\egd_top.BitStream_buffer.pc[5] ),
    .X(_3134_));
 sky130_fd_sc_hd__and2_1 _3601_ (.A(_3110_),
    .B(_3134_),
    .X(_3135_));
 sky130_fd_sc_hd__clkbuf_2 _3602_ (.A(_3135_),
    .X(_3136_));
 sky130_fd_sc_hd__buf_4 _3603_ (.A(_3136_),
    .X(_3137_));
 sky130_fd_sc_hd__clkbuf_4 _3604_ (.A(\egd_top.BitStream_buffer.BS_buffer[123] ),
    .X(_3138_));
 sky130_fd_sc_hd__and2_1 _3605_ (.A(_3114_),
    .B(_3134_),
    .X(_3139_));
 sky130_fd_sc_hd__buf_2 _3606_ (.A(_3139_),
    .X(_3140_));
 sky130_fd_sc_hd__buf_6 _3607_ (.A(_3140_),
    .X(_3141_));
 sky130_fd_sc_hd__buf_2 _3608_ (.A(_3134_),
    .X(_3142_));
 sky130_fd_sc_hd__and2_1 _3609_ (.A(_3124_),
    .B(_3142_),
    .X(_3143_));
 sky130_fd_sc_hd__buf_2 _3610_ (.A(_3143_),
    .X(_3144_));
 sky130_fd_sc_hd__inv_2 _3611_ (.A(_3144_),
    .Y(_3145_));
 sky130_fd_sc_hd__and2_1 _3612_ (.A(_3121_),
    .B(_3134_),
    .X(_3146_));
 sky130_fd_sc_hd__buf_6 _3613_ (.A(_3146_),
    .X(_3147_));
 sky130_fd_sc_hd__buf_6 _3614_ (.A(_3147_),
    .X(_3148_));
 sky130_fd_sc_hd__clkbuf_4 _3615_ (.A(\egd_top.BitStream_buffer.BS_buffer[121] ),
    .X(_3149_));
 sky130_fd_sc_hd__nand2_1 _3616_ (.A(_3148_),
    .B(_3149_),
    .Y(_3150_));
 sky130_fd_sc_hd__o21ai_1 _3617_ (.A1(_3003_),
    .A2(_3145_),
    .B1(_3150_),
    .Y(_3151_));
 sky130_fd_sc_hd__a221oi_1 _3618_ (.A1(_3133_),
    .A2(_3137_),
    .B1(_3138_),
    .B2(_3141_),
    .C1(_3151_),
    .Y(_3152_));
 sky130_fd_sc_hd__clkbuf_4 _3619_ (.A(\egd_top.BitStream_buffer.BS_buffer[114] ),
    .X(_3153_));
 sky130_fd_sc_hd__and2_1 _3620_ (.A(_3052_),
    .B(_3142_),
    .X(_3154_));
 sky130_fd_sc_hd__buf_2 _3621_ (.A(_3154_),
    .X(_3155_));
 sky130_fd_sc_hd__buf_4 _3622_ (.A(_3155_),
    .X(_3156_));
 sky130_fd_sc_hd__clkbuf_4 _3623_ (.A(\egd_top.BitStream_buffer.BS_buffer[115] ),
    .X(_3157_));
 sky130_fd_sc_hd__and2_1 _3624_ (.A(_3058_),
    .B(_3142_),
    .X(_3158_));
 sky130_fd_sc_hd__buf_2 _3625_ (.A(_3158_),
    .X(_3159_));
 sky130_fd_sc_hd__buf_4 _3626_ (.A(_3159_),
    .X(_3160_));
 sky130_fd_sc_hd__and2_1 _3627_ (.A(_3045_),
    .B(_3142_),
    .X(_3161_));
 sky130_fd_sc_hd__buf_4 _3628_ (.A(_3161_),
    .X(_3162_));
 sky130_fd_sc_hd__buf_6 _3629_ (.A(_3162_),
    .X(_3163_));
 sky130_fd_sc_hd__clkbuf_4 _3630_ (.A(\egd_top.BitStream_buffer.BS_buffer[113] ),
    .X(_3164_));
 sky130_fd_sc_hd__nand2_1 _3631_ (.A(_3163_),
    .B(_3164_),
    .Y(_3165_));
 sky130_fd_sc_hd__and2_1 _3632_ (.A(_3033_),
    .B(_3134_),
    .X(_3166_));
 sky130_fd_sc_hd__buf_2 _3633_ (.A(_3166_),
    .X(_3167_));
 sky130_fd_sc_hd__clkbuf_4 _3634_ (.A(_3167_),
    .X(_3168_));
 sky130_fd_sc_hd__clkbuf_4 _3635_ (.A(\egd_top.BitStream_buffer.BS_buffer[112] ),
    .X(_3169_));
 sky130_fd_sc_hd__nand2_1 _3636_ (.A(_3168_),
    .B(_3169_),
    .Y(_3170_));
 sky130_fd_sc_hd__nand2_1 _3637_ (.A(_3165_),
    .B(_3170_),
    .Y(_3171_));
 sky130_fd_sc_hd__a221oi_2 _3638_ (.A1(_3153_),
    .A2(_3156_),
    .B1(_3157_),
    .B2(_3160_),
    .C1(_3171_),
    .Y(_3172_));
 sky130_fd_sc_hd__clkbuf_4 _3639_ (.A(\egd_top.BitStream_buffer.BS_buffer[124] ),
    .X(_3173_));
 sky130_fd_sc_hd__and2_1 _3640_ (.A(_3067_),
    .B(_3134_),
    .X(_3174_));
 sky130_fd_sc_hd__clkbuf_2 _3641_ (.A(_3174_),
    .X(_3175_));
 sky130_fd_sc_hd__buf_2 _3642_ (.A(_3175_),
    .X(_3176_));
 sky130_fd_sc_hd__clkbuf_4 _3643_ (.A(\egd_top.BitStream_buffer.BS_buffer[125] ),
    .X(_3177_));
 sky130_fd_sc_hd__and2_1 _3644_ (.A(_3071_),
    .B(_3142_),
    .X(_3178_));
 sky130_fd_sc_hd__clkbuf_2 _3645_ (.A(_3178_),
    .X(_3179_));
 sky130_fd_sc_hd__buf_4 _3646_ (.A(_3179_),
    .X(_3180_));
 sky130_fd_sc_hd__and2_2 _3647_ (.A(_3076_),
    .B(_3134_),
    .X(_3181_));
 sky130_fd_sc_hd__inv_2 _3648_ (.A(_3181_),
    .Y(_3182_));
 sky130_fd_sc_hd__clkbuf_4 _3649_ (.A(_3182_),
    .X(_3183_));
 sky130_fd_sc_hd__and2_1 _3650_ (.A(_2931_),
    .B(_3134_),
    .X(_3184_));
 sky130_fd_sc_hd__clkbuf_2 _3651_ (.A(_3184_),
    .X(_3185_));
 sky130_fd_sc_hd__clkbuf_4 _3652_ (.A(_3185_),
    .X(_3186_));
 sky130_fd_sc_hd__clkbuf_4 _3653_ (.A(\egd_top.BitStream_buffer.BS_buffer[127] ),
    .X(_3187_));
 sky130_fd_sc_hd__nand2_1 _3654_ (.A(_3186_),
    .B(_3187_),
    .Y(_3188_));
 sky130_fd_sc_hd__o21ai_1 _3655_ (.A1(_3021_),
    .A2(_3183_),
    .B1(_3188_),
    .Y(_3189_));
 sky130_fd_sc_hd__a221oi_1 _3656_ (.A1(_3173_),
    .A2(_3176_),
    .B1(_3177_),
    .B2(_3180_),
    .C1(_3189_),
    .Y(_3190_));
 sky130_fd_sc_hd__clkbuf_4 _3657_ (.A(\egd_top.BitStream_buffer.BS_buffer[118] ),
    .X(_3191_));
 sky130_fd_sc_hd__and2_1 _3658_ (.A(_3096_),
    .B(_3142_),
    .X(_3192_));
 sky130_fd_sc_hd__buf_2 _3659_ (.A(_3192_),
    .X(_3193_));
 sky130_fd_sc_hd__clkbuf_4 _3660_ (.A(_3193_),
    .X(_3194_));
 sky130_fd_sc_hd__and2_1 _3661_ (.A(_3087_),
    .B(_3142_),
    .X(_3195_));
 sky130_fd_sc_hd__buf_2 _3662_ (.A(_3195_),
    .X(_3196_));
 sky130_fd_sc_hd__buf_6 _3663_ (.A(_3196_),
    .X(_3197_));
 sky130_fd_sc_hd__clkbuf_4 _3664_ (.A(\egd_top.BitStream_buffer.BS_buffer[119] ),
    .X(_3198_));
 sky130_fd_sc_hd__nand2_2 _3665_ (.A(_3104_),
    .B(_3142_),
    .Y(_3199_));
 sky130_fd_sc_hd__clkbuf_4 _3666_ (.A(_3199_),
    .X(_3200_));
 sky130_fd_sc_hd__and2_1 _3667_ (.A(_3090_),
    .B(_3134_),
    .X(_3201_));
 sky130_fd_sc_hd__clkbuf_2 _3668_ (.A(_3201_),
    .X(_3202_));
 sky130_fd_sc_hd__clkbuf_4 _3669_ (.A(_3202_),
    .X(_3203_));
 sky130_fd_sc_hd__clkbuf_4 _3670_ (.A(\egd_top.BitStream_buffer.BS_buffer[116] ),
    .X(_3204_));
 sky130_fd_sc_hd__nand2_1 _3671_ (.A(_3203_),
    .B(_3204_),
    .Y(_3205_));
 sky130_fd_sc_hd__o21ai_1 _3672_ (.A1(_2993_),
    .A2(_3200_),
    .B1(_3205_),
    .Y(_3206_));
 sky130_fd_sc_hd__a221oi_1 _3673_ (.A1(_3191_),
    .A2(_3194_),
    .B1(_3197_),
    .B2(_3198_),
    .C1(_3206_),
    .Y(_3207_));
 sky130_fd_sc_hd__and4_1 _3674_ (.A(_3152_),
    .B(_3172_),
    .C(_3190_),
    .D(_3207_),
    .X(_3208_));
 sky130_fd_sc_hd__nand2_1 _3675_ (.A(_3132_),
    .B(_3208_),
    .Y(_3209_));
 sky130_fd_sc_hd__buf_2 _3676_ (.A(\egd_top.BitStream_buffer.BS_buffer[68] ),
    .X(_3210_));
 sky130_fd_sc_hd__inv_2 _3677_ (.A(\egd_top.BitStream_buffer.pc[4] ),
    .Y(_3211_));
 sky130_fd_sc_hd__and3_2 _3678_ (.A(_3211_),
    .B(_3034_),
    .C(\egd_top.BitStream_buffer.pc[6] ),
    .X(_3212_));
 sky130_fd_sc_hd__buf_2 _3679_ (.A(_3212_),
    .X(_3213_));
 sky130_fd_sc_hd__and2_1 _3680_ (.A(_3090_),
    .B(_3213_),
    .X(_3214_));
 sky130_fd_sc_hd__clkbuf_2 _3681_ (.A(_3214_),
    .X(_3215_));
 sky130_fd_sc_hd__buf_2 _3682_ (.A(_3215_),
    .X(_3216_));
 sky130_fd_sc_hd__buf_2 _3683_ (.A(\egd_top.BitStream_buffer.BS_buffer[69] ),
    .X(_3217_));
 sky130_fd_sc_hd__nand2_1 _3684_ (.A(_3104_),
    .B(_3213_),
    .Y(_3218_));
 sky130_fd_sc_hd__inv_2 _3685_ (.A(_3218_),
    .Y(_3219_));
 sky130_fd_sc_hd__buf_2 _3686_ (.A(_3219_),
    .X(_3220_));
 sky130_fd_sc_hd__buf_2 _3687_ (.A(\egd_top.BitStream_buffer.BS_buffer[70] ),
    .X(_3221_));
 sky130_fd_sc_hd__and2_1 _3688_ (.A(_3096_),
    .B(_3213_),
    .X(_3222_));
 sky130_fd_sc_hd__clkbuf_2 _3689_ (.A(_3222_),
    .X(_3223_));
 sky130_fd_sc_hd__buf_6 _3690_ (.A(_3223_),
    .X(_3224_));
 sky130_fd_sc_hd__nand2_1 _3691_ (.A(_3087_),
    .B(_3213_),
    .Y(_3225_));
 sky130_fd_sc_hd__inv_2 _3692_ (.A(_3225_),
    .Y(_3226_));
 sky130_fd_sc_hd__buf_2 _3693_ (.A(\egd_top.BitStream_buffer.BS_buffer[71] ),
    .X(_3227_));
 sky130_fd_sc_hd__a22o_1 _3694_ (.A1(_3221_),
    .A2(_3224_),
    .B1(_3226_),
    .B2(_3227_),
    .X(_3228_));
 sky130_fd_sc_hd__a221oi_1 _3695_ (.A1(_3210_),
    .A2(_3216_),
    .B1(_3217_),
    .B2(_3220_),
    .C1(_3228_),
    .Y(_3229_));
 sky130_fd_sc_hd__buf_2 _3696_ (.A(\egd_top.BitStream_buffer.BS_buffer[66] ),
    .X(_3230_));
 sky130_fd_sc_hd__and2_1 _3697_ (.A(_3052_),
    .B(_3213_),
    .X(_3231_));
 sky130_fd_sc_hd__clkbuf_2 _3698_ (.A(_3231_),
    .X(_3232_));
 sky130_fd_sc_hd__buf_2 _3699_ (.A(_3232_),
    .X(_3233_));
 sky130_fd_sc_hd__and2_1 _3700_ (.A(_3058_),
    .B(_3213_),
    .X(_3234_));
 sky130_fd_sc_hd__clkbuf_2 _3701_ (.A(_3234_),
    .X(_3235_));
 sky130_fd_sc_hd__buf_2 _3702_ (.A(_3235_),
    .X(_3236_));
 sky130_fd_sc_hd__buf_2 _3703_ (.A(\egd_top.BitStream_buffer.BS_buffer[67] ),
    .X(_3237_));
 sky130_fd_sc_hd__clkinv_2 _3704_ (.A(\egd_top.BitStream_buffer.BS_buffer[65] ),
    .Y(_3238_));
 sky130_fd_sc_hd__nand2_2 _3705_ (.A(_3045_),
    .B(_3213_),
    .Y(_3239_));
 sky130_fd_sc_hd__buf_2 _3706_ (.A(_3239_),
    .X(_3240_));
 sky130_fd_sc_hd__and2_1 _3707_ (.A(_3033_),
    .B(_3212_),
    .X(_3241_));
 sky130_fd_sc_hd__clkbuf_2 _3708_ (.A(_3241_),
    .X(_3242_));
 sky130_fd_sc_hd__buf_6 _3709_ (.A(_3242_),
    .X(_3243_));
 sky130_fd_sc_hd__buf_2 _3710_ (.A(\egd_top.BitStream_buffer.BS_buffer[64] ),
    .X(_3244_));
 sky130_fd_sc_hd__nand2_1 _3711_ (.A(_3243_),
    .B(_3244_),
    .Y(_3245_));
 sky130_fd_sc_hd__o21ai_1 _3712_ (.A1(_3238_),
    .A2(_3240_),
    .B1(_3245_),
    .Y(_3246_));
 sky130_fd_sc_hd__a221oi_1 _3713_ (.A1(_3230_),
    .A2(_3233_),
    .B1(_3236_),
    .B2(_3237_),
    .C1(_3246_),
    .Y(_3247_));
 sky130_fd_sc_hd__clkbuf_4 _3714_ (.A(\egd_top.BitStream_buffer.BS_buffer[74] ),
    .X(_3248_));
 sky130_fd_sc_hd__and2_1 _3715_ (.A(_3110_),
    .B(_3212_),
    .X(_3249_));
 sky130_fd_sc_hd__clkbuf_2 _3716_ (.A(_3249_),
    .X(_3250_));
 sky130_fd_sc_hd__buf_6 _3717_ (.A(_3250_),
    .X(_3251_));
 sky130_fd_sc_hd__buf_2 _3718_ (.A(\egd_top.BitStream_buffer.BS_buffer[75] ),
    .X(_3252_));
 sky130_fd_sc_hd__and2_1 _3719_ (.A(_3114_),
    .B(_3212_),
    .X(_3253_));
 sky130_fd_sc_hd__buf_2 _3720_ (.A(_3253_),
    .X(_3254_));
 sky130_fd_sc_hd__buf_4 _3721_ (.A(_3254_),
    .X(_3255_));
 sky130_fd_sc_hd__clkbuf_4 _3722_ (.A(\egd_top.BitStream_buffer.BS_buffer[72] ),
    .X(_3256_));
 sky130_fd_sc_hd__clkinv_2 _3723_ (.A(_3256_),
    .Y(_3257_));
 sky130_fd_sc_hd__and2_1 _3724_ (.A(_3124_),
    .B(_3212_),
    .X(_3258_));
 sky130_fd_sc_hd__buf_2 _3725_ (.A(_3258_),
    .X(_3259_));
 sky130_fd_sc_hd__inv_2 _3726_ (.A(_3259_),
    .Y(_3260_));
 sky130_fd_sc_hd__and2_1 _3727_ (.A(_3121_),
    .B(_3212_),
    .X(_3261_));
 sky130_fd_sc_hd__clkbuf_2 _3728_ (.A(_3261_),
    .X(_3262_));
 sky130_fd_sc_hd__buf_6 _3729_ (.A(_3262_),
    .X(_3263_));
 sky130_fd_sc_hd__clkbuf_4 _3730_ (.A(\egd_top.BitStream_buffer.BS_buffer[73] ),
    .X(_3264_));
 sky130_fd_sc_hd__nand2_1 _3731_ (.A(_3263_),
    .B(_3264_),
    .Y(_3265_));
 sky130_fd_sc_hd__o21ai_1 _3732_ (.A1(_3257_),
    .A2(_3260_),
    .B1(_3265_),
    .Y(_3266_));
 sky130_fd_sc_hd__a221oi_1 _3733_ (.A1(_3248_),
    .A2(_3251_),
    .B1(_3252_),
    .B2(_3255_),
    .C1(_3266_),
    .Y(_3267_));
 sky130_fd_sc_hd__clkbuf_4 _3734_ (.A(\egd_top.BitStream_buffer.BS_buffer[76] ),
    .X(_3268_));
 sky130_fd_sc_hd__nand2_1 _3735_ (.A(_3067_),
    .B(_3213_),
    .Y(_3269_));
 sky130_fd_sc_hd__inv_2 _3736_ (.A(_3269_),
    .Y(_3270_));
 sky130_fd_sc_hd__buf_2 _3737_ (.A(_3270_),
    .X(_3271_));
 sky130_fd_sc_hd__buf_2 _3738_ (.A(\egd_top.BitStream_buffer.BS_buffer[77] ),
    .X(_3272_));
 sky130_fd_sc_hd__nand2_1 _3739_ (.A(_3071_),
    .B(_3213_),
    .Y(_3273_));
 sky130_fd_sc_hd__inv_2 _3740_ (.A(_3273_),
    .Y(_3274_));
 sky130_fd_sc_hd__buf_2 _3741_ (.A(_3274_),
    .X(_3275_));
 sky130_fd_sc_hd__clkbuf_4 _3742_ (.A(\egd_top.BitStream_buffer.BS_buffer[79] ),
    .X(_3276_));
 sky130_fd_sc_hd__clkinv_2 _3743_ (.A(_3276_),
    .Y(_3277_));
 sky130_fd_sc_hd__nand2_1 _3744_ (.A(_2931_),
    .B(_3213_),
    .Y(_3278_));
 sky130_fd_sc_hd__clkbuf_4 _3745_ (.A(_3278_),
    .X(_3279_));
 sky130_fd_sc_hd__and2_1 _3746_ (.A(_3076_),
    .B(_3212_),
    .X(_3280_));
 sky130_fd_sc_hd__clkbuf_2 _3747_ (.A(_3280_),
    .X(_3281_));
 sky130_fd_sc_hd__buf_2 _3748_ (.A(_3281_),
    .X(_3282_));
 sky130_fd_sc_hd__buf_2 _3749_ (.A(\egd_top.BitStream_buffer.BS_buffer[78] ),
    .X(_3283_));
 sky130_fd_sc_hd__nand2_1 _3750_ (.A(_3282_),
    .B(_3283_),
    .Y(_3284_));
 sky130_fd_sc_hd__o21ai_1 _3751_ (.A1(_3277_),
    .A2(_3279_),
    .B1(_3284_),
    .Y(_3285_));
 sky130_fd_sc_hd__a221oi_1 _3752_ (.A1(_3268_),
    .A2(_3271_),
    .B1(_3272_),
    .B2(_3275_),
    .C1(_3285_),
    .Y(_3286_));
 sky130_fd_sc_hd__and4_1 _3753_ (.A(_3229_),
    .B(_3247_),
    .C(_3267_),
    .D(_3286_),
    .X(_3287_));
 sky130_fd_sc_hd__buf_2 _3754_ (.A(\egd_top.BitStream_buffer.BS_buffer[82] ),
    .X(_3288_));
 sky130_fd_sc_hd__or3_2 _3755_ (.A(\egd_top.BitStream_buffer.pc[5] ),
    .B(_2932_),
    .C(_3211_),
    .X(_3289_));
 sky130_fd_sc_hd__buf_4 _3756_ (.A(_3289_),
    .X(_3290_));
 sky130_fd_sc_hd__nor2_2 _3757_ (.A(_3290_),
    .B(_3053_),
    .Y(_3291_));
 sky130_fd_sc_hd__buf_4 _3758_ (.A(_3291_),
    .X(_3292_));
 sky130_fd_sc_hd__buf_2 _3759_ (.A(\egd_top.BitStream_buffer.BS_buffer[83] ),
    .X(_3293_));
 sky130_fd_sc_hd__nor2_2 _3760_ (.A(_3290_),
    .B(_3059_),
    .Y(_3294_));
 sky130_fd_sc_hd__buf_6 _3761_ (.A(_3294_),
    .X(_3295_));
 sky130_fd_sc_hd__inv_2 _3762_ (.A(\egd_top.BitStream_buffer.BS_buffer[80] ),
    .Y(_3296_));
 sky130_fd_sc_hd__clkinv_2 _3763_ (.A(_3289_),
    .Y(_3297_));
 sky130_fd_sc_hd__nand2_2 _3764_ (.A(_3033_),
    .B(_3297_),
    .Y(_3298_));
 sky130_fd_sc_hd__buf_2 _3765_ (.A(_3298_),
    .X(_3299_));
 sky130_fd_sc_hd__nor2_2 _3766_ (.A(_3290_),
    .B(_3046_),
    .Y(_3300_));
 sky130_fd_sc_hd__buf_6 _3767_ (.A(_3300_),
    .X(_3301_));
 sky130_fd_sc_hd__clkbuf_4 _3768_ (.A(\egd_top.BitStream_buffer.BS_buffer[81] ),
    .X(_3302_));
 sky130_fd_sc_hd__nand2_1 _3769_ (.A(_3301_),
    .B(_3302_),
    .Y(_3303_));
 sky130_fd_sc_hd__o21ai_1 _3770_ (.A1(_3296_),
    .A2(_3299_),
    .B1(_3303_),
    .Y(_3304_));
 sky130_fd_sc_hd__a221oi_1 _3771_ (.A1(_3288_),
    .A2(_3292_),
    .B1(_3293_),
    .B2(_3295_),
    .C1(_3304_),
    .Y(_3305_));
 sky130_fd_sc_hd__clkinv_2 _3772_ (.A(\egd_top.BitStream_buffer.BS_buffer[87] ),
    .Y(_3306_));
 sky130_fd_sc_hd__nand2_2 _3773_ (.A(_3087_),
    .B(_3297_),
    .Y(_3307_));
 sky130_fd_sc_hd__clkbuf_4 _3774_ (.A(_3307_),
    .X(_3308_));
 sky130_fd_sc_hd__nor2_2 _3775_ (.A(_3290_),
    .B(_3097_),
    .Y(_3309_));
 sky130_fd_sc_hd__buf_4 _3776_ (.A(_3309_),
    .X(_3310_));
 sky130_fd_sc_hd__buf_2 _3777_ (.A(\egd_top.BitStream_buffer.BS_buffer[86] ),
    .X(_3311_));
 sky130_fd_sc_hd__nand2_1 _3778_ (.A(_3310_),
    .B(_3311_),
    .Y(_3312_));
 sky130_fd_sc_hd__nor2_2 _3779_ (.A(_3289_),
    .B(_3091_),
    .Y(_3313_));
 sky130_fd_sc_hd__clkbuf_4 _3780_ (.A(_3313_),
    .X(_3314_));
 sky130_fd_sc_hd__clkbuf_4 _3781_ (.A(\egd_top.BitStream_buffer.BS_buffer[84] ),
    .X(_3315_));
 sky130_fd_sc_hd__nand2_1 _3782_ (.A(_3314_),
    .B(_3315_),
    .Y(_3316_));
 sky130_fd_sc_hd__clkinv_2 _3783_ (.A(\egd_top.BitStream_buffer.BS_buffer[85] ),
    .Y(_3317_));
 sky130_fd_sc_hd__nand2_2 _3784_ (.A(_3104_),
    .B(_3297_),
    .Y(_3318_));
 sky130_fd_sc_hd__buf_2 _3785_ (.A(_3318_),
    .X(_3319_));
 sky130_fd_sc_hd__or2_1 _3786_ (.A(_3317_),
    .B(_3319_),
    .X(_3320_));
 sky130_fd_sc_hd__o2111a_1 _3787_ (.A1(_3306_),
    .A2(_3308_),
    .B1(_3312_),
    .C1(_3316_),
    .D1(_3320_),
    .X(_3321_));
 sky130_fd_sc_hd__clkbuf_4 _3788_ (.A(\egd_top.BitStream_buffer.BS_buffer[90] ),
    .X(_3322_));
 sky130_fd_sc_hd__nor2_2 _3789_ (.A(_3290_),
    .B(_3111_),
    .Y(_3323_));
 sky130_fd_sc_hd__buf_2 _3790_ (.A(_3323_),
    .X(_3324_));
 sky130_fd_sc_hd__nor2_2 _3791_ (.A(_3290_),
    .B(_3115_),
    .Y(_3325_));
 sky130_fd_sc_hd__buf_2 _3792_ (.A(_3325_),
    .X(_3326_));
 sky130_fd_sc_hd__buf_2 _3793_ (.A(\egd_top.BitStream_buffer.BS_buffer[91] ),
    .X(_3327_));
 sky130_fd_sc_hd__clkinv_2 _3794_ (.A(\egd_top.BitStream_buffer.BS_buffer[89] ),
    .Y(_3328_));
 sky130_fd_sc_hd__nand2_2 _3795_ (.A(_3121_),
    .B(_3297_),
    .Y(_3329_));
 sky130_fd_sc_hd__clkbuf_4 _3796_ (.A(_3329_),
    .X(_3330_));
 sky130_fd_sc_hd__nand2_1 _3797_ (.A(_3124_),
    .B(_3297_),
    .Y(_3331_));
 sky130_fd_sc_hd__clkinv_2 _3798_ (.A(_3331_),
    .Y(_3332_));
 sky130_fd_sc_hd__buf_2 _3799_ (.A(_3332_),
    .X(_3333_));
 sky130_fd_sc_hd__buf_2 _3800_ (.A(\egd_top.BitStream_buffer.BS_buffer[88] ),
    .X(_3334_));
 sky130_fd_sc_hd__nand2_1 _3801_ (.A(_3333_),
    .B(_3334_),
    .Y(_3335_));
 sky130_fd_sc_hd__o21ai_1 _3802_ (.A1(_3328_),
    .A2(_3330_),
    .B1(_3335_),
    .Y(_3336_));
 sky130_fd_sc_hd__a221oi_1 _3803_ (.A1(_3322_),
    .A2(_3324_),
    .B1(_3326_),
    .B2(_3327_),
    .C1(_3336_),
    .Y(_3337_));
 sky130_fd_sc_hd__buf_2 _3804_ (.A(\egd_top.BitStream_buffer.BS_buffer[94] ),
    .X(_3338_));
 sky130_fd_sc_hd__nor2_2 _3805_ (.A(_3290_),
    .B(_3077_),
    .Y(_3339_));
 sky130_fd_sc_hd__buf_2 _3806_ (.A(_3339_),
    .X(_3340_));
 sky130_fd_sc_hd__buf_2 _3807_ (.A(\egd_top.BitStream_buffer.BS_buffer[95] ),
    .X(_3341_));
 sky130_fd_sc_hd__nor2_2 _3808_ (.A(_3290_),
    .B(_3079_),
    .Y(_0322_));
 sky130_fd_sc_hd__clkbuf_4 _3809_ (.A(_0322_),
    .X(_0323_));
 sky130_fd_sc_hd__inv_2 _3810_ (.A(\egd_top.BitStream_buffer.BS_buffer[93] ),
    .Y(_0324_));
 sky130_fd_sc_hd__nor2_1 _3811_ (.A(_3290_),
    .B(_3072_),
    .Y(_0325_));
 sky130_fd_sc_hd__inv_2 _3812_ (.A(_0325_),
    .Y(_0326_));
 sky130_fd_sc_hd__clkbuf_4 _3813_ (.A(_0326_),
    .X(_0327_));
 sky130_fd_sc_hd__nor2_2 _3814_ (.A(_3290_),
    .B(_3068_),
    .Y(_0328_));
 sky130_fd_sc_hd__buf_4 _3815_ (.A(_0328_),
    .X(_0329_));
 sky130_fd_sc_hd__clkbuf_4 _3816_ (.A(\egd_top.BitStream_buffer.BS_buffer[92] ),
    .X(_0330_));
 sky130_fd_sc_hd__nand2_1 _3817_ (.A(_0329_),
    .B(_0330_),
    .Y(_0331_));
 sky130_fd_sc_hd__o21ai_1 _3818_ (.A1(_0324_),
    .A2(_0327_),
    .B1(_0331_),
    .Y(_0332_));
 sky130_fd_sc_hd__a221oi_1 _3819_ (.A1(_3338_),
    .A2(_3340_),
    .B1(_3341_),
    .B2(_0323_),
    .C1(_0332_),
    .Y(_0333_));
 sky130_fd_sc_hd__and4_1 _3820_ (.A(_3305_),
    .B(_3321_),
    .C(_3337_),
    .D(_0333_),
    .X(_0334_));
 sky130_fd_sc_hd__nand2_1 _3821_ (.A(_3287_),
    .B(_0334_),
    .Y(_0335_));
 sky130_fd_sc_hd__nor2_1 _3822_ (.A(_3209_),
    .B(_0335_),
    .Y(_0336_));
 sky130_fd_sc_hd__clkbuf_4 _3823_ (.A(\egd_top.BitStream_buffer.BS_buffer[36] ),
    .X(_0337_));
 sky130_fd_sc_hd__and3_2 _3824_ (.A(_2932_),
    .B(_3211_),
    .C(\egd_top.BitStream_buffer.pc[5] ),
    .X(_0338_));
 sky130_fd_sc_hd__buf_2 _3825_ (.A(_0338_),
    .X(_0339_));
 sky130_fd_sc_hd__and2_1 _3826_ (.A(_3090_),
    .B(_0339_),
    .X(_0340_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _3827_ (.A(_0340_),
    .X(_0341_));
 sky130_fd_sc_hd__buf_2 _3828_ (.A(_0341_),
    .X(_0342_));
 sky130_fd_sc_hd__and2_1 _3829_ (.A(_3104_),
    .B(_0339_),
    .X(_0343_));
 sky130_fd_sc_hd__clkbuf_2 _3830_ (.A(_0343_),
    .X(_0344_));
 sky130_fd_sc_hd__buf_6 _3831_ (.A(_0344_),
    .X(_0345_));
 sky130_fd_sc_hd__clkbuf_4 _3832_ (.A(\egd_top.BitStream_buffer.BS_buffer[37] ),
    .X(_0346_));
 sky130_fd_sc_hd__clkbuf_4 _3833_ (.A(\egd_top.BitStream_buffer.BS_buffer[39] ),
    .X(_0347_));
 sky130_fd_sc_hd__clkinv_2 _3834_ (.A(_0347_),
    .Y(_0348_));
 sky130_fd_sc_hd__nand2_1 _3835_ (.A(_3087_),
    .B(_0339_),
    .Y(_0349_));
 sky130_fd_sc_hd__clkbuf_4 _3836_ (.A(_0349_),
    .X(_0350_));
 sky130_fd_sc_hd__nand2_1 _3837_ (.A(_3096_),
    .B(_0339_),
    .Y(_0351_));
 sky130_fd_sc_hd__inv_2 _3838_ (.A(_0351_),
    .Y(_0352_));
 sky130_fd_sc_hd__buf_2 _3839_ (.A(_0352_),
    .X(_0353_));
 sky130_fd_sc_hd__clkbuf_4 _3840_ (.A(\egd_top.BitStream_buffer.BS_buffer[38] ),
    .X(_0354_));
 sky130_fd_sc_hd__nand2_1 _3841_ (.A(_0353_),
    .B(_0354_),
    .Y(_0355_));
 sky130_fd_sc_hd__o21ai_1 _3842_ (.A1(_0348_),
    .A2(_0350_),
    .B1(_0355_),
    .Y(_0356_));
 sky130_fd_sc_hd__a221oi_1 _3843_ (.A1(_0337_),
    .A2(_0342_),
    .B1(_0345_),
    .B2(_0346_),
    .C1(_0356_),
    .Y(_0357_));
 sky130_fd_sc_hd__and2_1 _3844_ (.A(_3052_),
    .B(_0338_),
    .X(_0358_));
 sky130_fd_sc_hd__clkbuf_2 _3845_ (.A(_0358_),
    .X(_0359_));
 sky130_fd_sc_hd__buf_2 _3846_ (.A(_0359_),
    .X(_0360_));
 sky130_fd_sc_hd__and2_1 _3847_ (.A(_3058_),
    .B(_0338_),
    .X(_0361_));
 sky130_fd_sc_hd__clkbuf_2 _3848_ (.A(_0361_),
    .X(_0362_));
 sky130_fd_sc_hd__buf_2 _3849_ (.A(_0362_),
    .X(_0363_));
 sky130_fd_sc_hd__clkbuf_4 _3850_ (.A(\egd_top.BitStream_buffer.BS_buffer[35] ),
    .X(_0364_));
 sky130_fd_sc_hd__clkbuf_4 _3851_ (.A(\egd_top.BitStream_buffer.BS_buffer[33] ),
    .X(_0365_));
 sky130_fd_sc_hd__clkinv_2 _3852_ (.A(_0365_),
    .Y(_0366_));
 sky130_fd_sc_hd__nand2_2 _3853_ (.A(_3045_),
    .B(_0339_),
    .Y(_0367_));
 sky130_fd_sc_hd__buf_2 _3854_ (.A(_0367_),
    .X(_0368_));
 sky130_fd_sc_hd__and2_1 _3855_ (.A(_3033_),
    .B(_0338_),
    .X(_0369_));
 sky130_fd_sc_hd__clkbuf_2 _3856_ (.A(_0369_),
    .X(_0370_));
 sky130_fd_sc_hd__buf_2 _3857_ (.A(_0370_),
    .X(_0371_));
 sky130_fd_sc_hd__nand2_1 _3858_ (.A(_0371_),
    .B(\egd_top.BitStream_buffer.BS_buffer[32] ),
    .Y(_0372_));
 sky130_fd_sc_hd__o21ai_1 _3859_ (.A1(_0366_),
    .A2(_0368_),
    .B1(_0372_),
    .Y(_0373_));
 sky130_fd_sc_hd__a221oi_1 _3860_ (.A1(\egd_top.BitStream_buffer.BS_buffer[34] ),
    .A2(_0360_),
    .B1(_0363_),
    .B2(_0364_),
    .C1(_0373_),
    .Y(_0374_));
 sky130_fd_sc_hd__clkbuf_4 _3861_ (.A(\egd_top.BitStream_buffer.BS_buffer[40] ),
    .X(_0375_));
 sky130_fd_sc_hd__and2_1 _3862_ (.A(_3124_),
    .B(_0338_),
    .X(_0376_));
 sky130_fd_sc_hd__clkbuf_2 _3863_ (.A(_0376_),
    .X(_0377_));
 sky130_fd_sc_hd__clkbuf_4 _3864_ (.A(_0377_),
    .X(_0378_));
 sky130_fd_sc_hd__clkbuf_4 _3865_ (.A(\egd_top.BitStream_buffer.BS_buffer[41] ),
    .X(_0379_));
 sky130_fd_sc_hd__nand2_2 _3866_ (.A(_3121_),
    .B(_0338_),
    .Y(_0380_));
 sky130_fd_sc_hd__inv_2 _3867_ (.A(_0380_),
    .Y(_0381_));
 sky130_fd_sc_hd__buf_6 _3868_ (.A(_0381_),
    .X(_0382_));
 sky130_fd_sc_hd__clkinv_2 _3869_ (.A(\egd_top.BitStream_buffer.BS_buffer[43] ),
    .Y(_0383_));
 sky130_fd_sc_hd__nand2_1 _3870_ (.A(_3114_),
    .B(_0339_),
    .Y(_0384_));
 sky130_fd_sc_hd__clkbuf_4 _3871_ (.A(_0384_),
    .X(_0385_));
 sky130_fd_sc_hd__and2_1 _3872_ (.A(_3110_),
    .B(_0338_),
    .X(_0386_));
 sky130_fd_sc_hd__clkbuf_2 _3873_ (.A(_0386_),
    .X(_0387_));
 sky130_fd_sc_hd__buf_2 _3874_ (.A(_0387_),
    .X(_0388_));
 sky130_fd_sc_hd__buf_2 _3875_ (.A(\egd_top.BitStream_buffer.BS_buffer[42] ),
    .X(_0389_));
 sky130_fd_sc_hd__nand2_1 _3876_ (.A(_0388_),
    .B(_0389_),
    .Y(_0390_));
 sky130_fd_sc_hd__o21ai_1 _3877_ (.A1(_0383_),
    .A2(_0385_),
    .B1(_0390_),
    .Y(_0391_));
 sky130_fd_sc_hd__a221oi_1 _3878_ (.A1(_0375_),
    .A2(_0378_),
    .B1(_0379_),
    .B2(_0382_),
    .C1(_0391_),
    .Y(_0392_));
 sky130_fd_sc_hd__buf_2 _3879_ (.A(\egd_top.BitStream_buffer.BS_buffer[44] ),
    .X(_0393_));
 sky130_fd_sc_hd__and2_1 _3880_ (.A(_3067_),
    .B(_0338_),
    .X(_0394_));
 sky130_fd_sc_hd__clkbuf_2 _3881_ (.A(_0394_),
    .X(_0395_));
 sky130_fd_sc_hd__buf_2 _3882_ (.A(_0395_),
    .X(_0396_));
 sky130_fd_sc_hd__and2_1 _3883_ (.A(_3071_),
    .B(_0338_),
    .X(_0397_));
 sky130_fd_sc_hd__clkbuf_2 _3884_ (.A(_0397_),
    .X(_0398_));
 sky130_fd_sc_hd__buf_2 _3885_ (.A(_0398_),
    .X(_0399_));
 sky130_fd_sc_hd__clkbuf_4 _3886_ (.A(\egd_top.BitStream_buffer.BS_buffer[45] ),
    .X(_0400_));
 sky130_fd_sc_hd__clkinv_2 _3887_ (.A(\egd_top.BitStream_buffer.BS_buffer[47] ),
    .Y(_0401_));
 sky130_fd_sc_hd__nand2_2 _3888_ (.A(_2931_),
    .B(_0339_),
    .Y(_0402_));
 sky130_fd_sc_hd__clkbuf_4 _3889_ (.A(_0402_),
    .X(_0403_));
 sky130_fd_sc_hd__nand2_1 _3890_ (.A(_3076_),
    .B(_0339_),
    .Y(_0404_));
 sky130_fd_sc_hd__inv_2 _3891_ (.A(_0404_),
    .Y(_0405_));
 sky130_fd_sc_hd__buf_2 _3892_ (.A(_0405_),
    .X(_0406_));
 sky130_fd_sc_hd__buf_2 _3893_ (.A(\egd_top.BitStream_buffer.BS_buffer[46] ),
    .X(_0407_));
 sky130_fd_sc_hd__nand2_1 _3894_ (.A(_0406_),
    .B(_0407_),
    .Y(_0408_));
 sky130_fd_sc_hd__o21ai_1 _3895_ (.A1(_0401_),
    .A2(_0403_),
    .B1(_0408_),
    .Y(_0409_));
 sky130_fd_sc_hd__a221oi_1 _3896_ (.A1(_0393_),
    .A2(_0396_),
    .B1(_0399_),
    .B2(_0400_),
    .C1(_0409_),
    .Y(_0410_));
 sky130_fd_sc_hd__and4_1 _3897_ (.A(_0357_),
    .B(_0374_),
    .C(_0392_),
    .D(_0410_),
    .X(_0411_));
 sky130_fd_sc_hd__clkbuf_4 _3898_ (.A(\egd_top.BitStream_buffer.BS_buffer[50] ),
    .X(_0412_));
 sky130_fd_sc_hd__and2_1 _3899_ (.A(_3052_),
    .B(_2933_),
    .X(_0413_));
 sky130_fd_sc_hd__clkbuf_2 _3900_ (.A(_0413_),
    .X(_0414_));
 sky130_fd_sc_hd__buf_2 _3901_ (.A(_0414_),
    .X(_0415_));
 sky130_fd_sc_hd__buf_2 _3902_ (.A(\egd_top.BitStream_buffer.BS_buffer[51] ),
    .X(_0416_));
 sky130_fd_sc_hd__and2_1 _3903_ (.A(_3058_),
    .B(_2933_),
    .X(_0417_));
 sky130_fd_sc_hd__clkbuf_2 _3904_ (.A(_0417_),
    .X(_0418_));
 sky130_fd_sc_hd__buf_2 _3905_ (.A(_0418_),
    .X(_0419_));
 sky130_fd_sc_hd__clkinv_2 _3906_ (.A(\egd_top.BitStream_buffer.BS_buffer[49] ),
    .Y(_0420_));
 sky130_fd_sc_hd__nand2_2 _3907_ (.A(_3045_),
    .B(_2934_),
    .Y(_0421_));
 sky130_fd_sc_hd__buf_2 _3908_ (.A(_0421_),
    .X(_0422_));
 sky130_fd_sc_hd__inv_2 _3909_ (.A(\egd_top.BitStream_buffer.BS_buffer[48] ),
    .Y(_0423_));
 sky130_fd_sc_hd__nand2_1 _3910_ (.A(_3033_),
    .B(_2934_),
    .Y(_0424_));
 sky130_fd_sc_hd__clkbuf_2 _3911_ (.A(_0424_),
    .X(_0425_));
 sky130_fd_sc_hd__or2_1 _3912_ (.A(_0423_),
    .B(_0425_),
    .X(_0426_));
 sky130_fd_sc_hd__o21ai_1 _3913_ (.A1(_0420_),
    .A2(_0422_),
    .B1(_0426_),
    .Y(_0427_));
 sky130_fd_sc_hd__a221oi_1 _3914_ (.A1(_0412_),
    .A2(_0415_),
    .B1(_0416_),
    .B2(_0419_),
    .C1(_0427_),
    .Y(_0428_));
 sky130_fd_sc_hd__buf_2 _3915_ (.A(\egd_top.BitStream_buffer.BS_buffer[54] ),
    .X(_0429_));
 sky130_fd_sc_hd__and2_1 _3916_ (.A(_3096_),
    .B(_2933_),
    .X(_0430_));
 sky130_fd_sc_hd__clkbuf_2 _3917_ (.A(_0430_),
    .X(_0431_));
 sky130_fd_sc_hd__buf_2 _3918_ (.A(_0431_),
    .X(_0432_));
 sky130_fd_sc_hd__and2_1 _3919_ (.A(_3087_),
    .B(_2933_),
    .X(_0433_));
 sky130_fd_sc_hd__buf_6 _3920_ (.A(_0433_),
    .X(_0434_));
 sky130_fd_sc_hd__buf_6 _3921_ (.A(_0434_),
    .X(_0435_));
 sky130_fd_sc_hd__clkbuf_4 _3922_ (.A(\egd_top.BitStream_buffer.BS_buffer[55] ),
    .X(_0436_));
 sky130_fd_sc_hd__clkinv_2 _3923_ (.A(\egd_top.BitStream_buffer.BS_buffer[53] ),
    .Y(_0437_));
 sky130_fd_sc_hd__nand2_2 _3924_ (.A(_3104_),
    .B(_2934_),
    .Y(_0438_));
 sky130_fd_sc_hd__clkbuf_4 _3925_ (.A(_0438_),
    .X(_0439_));
 sky130_fd_sc_hd__and2_1 _3926_ (.A(_3090_),
    .B(_2933_),
    .X(_0440_));
 sky130_fd_sc_hd__clkbuf_2 _3927_ (.A(_0440_),
    .X(_0441_));
 sky130_fd_sc_hd__buf_2 _3928_ (.A(_0441_),
    .X(_0442_));
 sky130_fd_sc_hd__clkbuf_4 _3929_ (.A(\egd_top.BitStream_buffer.BS_buffer[52] ),
    .X(_0443_));
 sky130_fd_sc_hd__nand2_1 _3930_ (.A(_0442_),
    .B(_0443_),
    .Y(_0444_));
 sky130_fd_sc_hd__o21ai_1 _3931_ (.A1(_0437_),
    .A2(_0439_),
    .B1(_0444_),
    .Y(_0445_));
 sky130_fd_sc_hd__a221oi_1 _3932_ (.A1(_0429_),
    .A2(_0432_),
    .B1(_0435_),
    .B2(_0436_),
    .C1(_0445_),
    .Y(_0446_));
 sky130_fd_sc_hd__clkbuf_4 _3933_ (.A(\egd_top.BitStream_buffer.BS_buffer[59] ),
    .X(_0447_));
 sky130_fd_sc_hd__clkinv_2 _3934_ (.A(_0447_),
    .Y(_0448_));
 sky130_fd_sc_hd__nand2_2 _3935_ (.A(_3114_),
    .B(_2934_),
    .Y(_0449_));
 sky130_fd_sc_hd__buf_2 _3936_ (.A(_0449_),
    .X(_0450_));
 sky130_fd_sc_hd__nand2_1 _3937_ (.A(_3124_),
    .B(_2934_),
    .Y(_0451_));
 sky130_fd_sc_hd__clkinv_2 _3938_ (.A(_0451_),
    .Y(_0452_));
 sky130_fd_sc_hd__buf_2 _3939_ (.A(_0452_),
    .X(_0453_));
 sky130_fd_sc_hd__buf_2 _3940_ (.A(\egd_top.BitStream_buffer.BS_buffer[56] ),
    .X(_0454_));
 sky130_fd_sc_hd__nand2_1 _3941_ (.A(_0453_),
    .B(_0454_),
    .Y(_0455_));
 sky130_fd_sc_hd__nand2_1 _3942_ (.A(_3110_),
    .B(_2934_),
    .Y(_0456_));
 sky130_fd_sc_hd__clkinv_2 _3943_ (.A(_0456_),
    .Y(_0457_));
 sky130_fd_sc_hd__buf_2 _3944_ (.A(_0457_),
    .X(_0458_));
 sky130_fd_sc_hd__buf_2 _3945_ (.A(\egd_top.BitStream_buffer.BS_buffer[58] ),
    .X(_0459_));
 sky130_fd_sc_hd__nand2_1 _3946_ (.A(_0458_),
    .B(_0459_),
    .Y(_0460_));
 sky130_fd_sc_hd__clkbuf_4 _3947_ (.A(\egd_top.BitStream_buffer.BS_buffer[57] ),
    .X(_0461_));
 sky130_fd_sc_hd__clkinv_2 _3948_ (.A(_0461_),
    .Y(_0462_));
 sky130_fd_sc_hd__nand2_2 _3949_ (.A(_3121_),
    .B(_2933_),
    .Y(_0463_));
 sky130_fd_sc_hd__buf_2 _3950_ (.A(_0463_),
    .X(_0464_));
 sky130_fd_sc_hd__or2_1 _3951_ (.A(_0462_),
    .B(_0464_),
    .X(_0465_));
 sky130_fd_sc_hd__o2111a_1 _3952_ (.A1(_0448_),
    .A2(_0450_),
    .B1(_0455_),
    .C1(_0460_),
    .D1(_0465_),
    .X(_0466_));
 sky130_fd_sc_hd__clkbuf_4 _3953_ (.A(\egd_top.BitStream_buffer.BS_buffer[60] ),
    .X(_0467_));
 sky130_fd_sc_hd__nand2_1 _3954_ (.A(_3067_),
    .B(_2934_),
    .Y(_0468_));
 sky130_fd_sc_hd__inv_2 _3955_ (.A(_0468_),
    .Y(_0469_));
 sky130_fd_sc_hd__buf_2 _3956_ (.A(_0469_),
    .X(_0470_));
 sky130_fd_sc_hd__clkbuf_4 _3957_ (.A(\egd_top.BitStream_buffer.BS_buffer[61] ),
    .X(_0471_));
 sky130_fd_sc_hd__nand2_2 _3958_ (.A(_3071_),
    .B(_2934_),
    .Y(_0472_));
 sky130_fd_sc_hd__inv_2 _3959_ (.A(_0472_),
    .Y(_0473_));
 sky130_fd_sc_hd__clkinv_2 _3960_ (.A(\egd_top.BitStream_buffer.BS_buffer[63] ),
    .Y(_0474_));
 sky130_fd_sc_hd__and2_1 _3961_ (.A(_3076_),
    .B(_2933_),
    .X(_0475_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _3962_ (.A(_0475_),
    .X(_0476_));
 sky130_fd_sc_hd__buf_2 _3963_ (.A(_0476_),
    .X(_0477_));
 sky130_fd_sc_hd__buf_2 _3964_ (.A(\egd_top.BitStream_buffer.BS_buffer[62] ),
    .X(_0478_));
 sky130_fd_sc_hd__nand2_1 _3965_ (.A(_0477_),
    .B(_0478_),
    .Y(_0479_));
 sky130_fd_sc_hd__o21ai_1 _3966_ (.A1(_0474_),
    .A2(_2935_),
    .B1(_0479_),
    .Y(_0480_));
 sky130_fd_sc_hd__a221oi_1 _3967_ (.A1(_0467_),
    .A2(_0470_),
    .B1(_0471_),
    .B2(_0473_),
    .C1(_0480_),
    .Y(_0481_));
 sky130_fd_sc_hd__and4_1 _3968_ (.A(_0428_),
    .B(_0446_),
    .C(_0466_),
    .D(_0481_),
    .X(_0482_));
 sky130_fd_sc_hd__nand2_1 _3969_ (.A(_0411_),
    .B(_0482_),
    .Y(_0483_));
 sky130_fd_sc_hd__and3_2 _3970_ (.A(_2932_),
    .B(_3034_),
    .C(\egd_top.BitStream_buffer.pc[4] ),
    .X(_0484_));
 sky130_fd_sc_hd__and2_1 _3971_ (.A(_3033_),
    .B(_0484_),
    .X(_0485_));
 sky130_fd_sc_hd__clkbuf_2 _3972_ (.A(_0485_),
    .X(_0486_));
 sky130_fd_sc_hd__buf_2 _3973_ (.A(_0486_),
    .X(_0487_));
 sky130_fd_sc_hd__clkinv_4 _3974_ (.A(_0484_),
    .Y(_0488_));
 sky130_fd_sc_hd__nor2_2 _3975_ (.A(_0488_),
    .B(_3046_),
    .Y(_0489_));
 sky130_fd_sc_hd__buf_6 _3976_ (.A(_0489_),
    .X(_0490_));
 sky130_fd_sc_hd__clkbuf_4 _3977_ (.A(\egd_top.BitStream_buffer.BS_buffer[18] ),
    .X(_0491_));
 sky130_fd_sc_hd__clkinv_2 _3978_ (.A(_0491_),
    .Y(_0492_));
 sky130_fd_sc_hd__nor2_1 _3979_ (.A(_0488_),
    .B(_3053_),
    .Y(_0493_));
 sky130_fd_sc_hd__inv_2 _3980_ (.A(_0493_),
    .Y(_0494_));
 sky130_fd_sc_hd__buf_2 _3981_ (.A(_0494_),
    .X(_0495_));
 sky130_fd_sc_hd__nor2_2 _3982_ (.A(_0488_),
    .B(_3059_),
    .Y(_0496_));
 sky130_fd_sc_hd__buf_4 _3983_ (.A(_0496_),
    .X(_0497_));
 sky130_fd_sc_hd__clkbuf_4 _3984_ (.A(\egd_top.BitStream_buffer.BS_buffer[19] ),
    .X(_0498_));
 sky130_fd_sc_hd__nand2_1 _3985_ (.A(_0497_),
    .B(_0498_),
    .Y(_0499_));
 sky130_fd_sc_hd__o21ai_1 _3986_ (.A1(_0492_),
    .A2(_0495_),
    .B1(_0499_),
    .Y(_0500_));
 sky130_fd_sc_hd__a221oi_1 _3987_ (.A1(\egd_top.BitStream_buffer.BS_buffer[16] ),
    .A2(_0487_),
    .B1(\egd_top.BitStream_buffer.BS_buffer[17] ),
    .B2(_0490_),
    .C1(_0500_),
    .Y(_0501_));
 sky130_fd_sc_hd__clkbuf_4 _3988_ (.A(\egd_top.BitStream_buffer.BS_buffer[20] ),
    .X(_0502_));
 sky130_fd_sc_hd__nor2_2 _3989_ (.A(_0488_),
    .B(_3091_),
    .Y(_0503_));
 sky130_fd_sc_hd__buf_2 _3990_ (.A(_0503_),
    .X(_0504_));
 sky130_fd_sc_hd__clkbuf_4 _3991_ (.A(\egd_top.BitStream_buffer.BS_buffer[21] ),
    .X(_0505_));
 sky130_fd_sc_hd__nand2_1 _3992_ (.A(_3104_),
    .B(_0484_),
    .Y(_0506_));
 sky130_fd_sc_hd__inv_2 _3993_ (.A(_0506_),
    .Y(_0507_));
 sky130_fd_sc_hd__buf_6 _3994_ (.A(_0507_),
    .X(_0508_));
 sky130_fd_sc_hd__clkbuf_4 _3995_ (.A(\egd_top.BitStream_buffer.BS_buffer[23] ),
    .X(_0509_));
 sky130_fd_sc_hd__clkinv_2 _3996_ (.A(_0509_),
    .Y(_0510_));
 sky130_fd_sc_hd__nand2_1 _3997_ (.A(_3087_),
    .B(_0484_),
    .Y(_0511_));
 sky130_fd_sc_hd__clkbuf_4 _3998_ (.A(_0511_),
    .X(_0512_));
 sky130_fd_sc_hd__nor2_2 _3999_ (.A(_0488_),
    .B(_3097_),
    .Y(_0513_));
 sky130_fd_sc_hd__buf_4 _4000_ (.A(_0513_),
    .X(_0514_));
 sky130_fd_sc_hd__clkbuf_4 _4001_ (.A(\egd_top.BitStream_buffer.BS_buffer[22] ),
    .X(_0515_));
 sky130_fd_sc_hd__nand2_1 _4002_ (.A(_0514_),
    .B(_0515_),
    .Y(_0516_));
 sky130_fd_sc_hd__o21ai_1 _4003_ (.A1(_0510_),
    .A2(_0512_),
    .B1(_0516_),
    .Y(_0517_));
 sky130_fd_sc_hd__a221oi_1 _4004_ (.A1(_0502_),
    .A2(_0504_),
    .B1(_0505_),
    .B2(_0508_),
    .C1(_0517_),
    .Y(_0518_));
 sky130_fd_sc_hd__clkbuf_4 _4005_ (.A(\egd_top.BitStream_buffer.BS_buffer[24] ),
    .X(_0519_));
 sky130_fd_sc_hd__clkinv_2 _4006_ (.A(_0519_),
    .Y(_0520_));
 sky130_fd_sc_hd__and3_2 _4007_ (.A(_0484_),
    .B(_3031_),
    .C(\egd_top.BitStream_buffer.pc[3] ),
    .X(_0521_));
 sky130_fd_sc_hd__nand2_2 _4008_ (.A(_0521_),
    .B(_3030_),
    .Y(_0522_));
 sky130_fd_sc_hd__buf_2 _4009_ (.A(_0522_),
    .X(_0523_));
 sky130_fd_sc_hd__inv_2 _4010_ (.A(\egd_top.BitStream_buffer.BS_buffer[27] ),
    .Y(_0524_));
 sky130_fd_sc_hd__nand2_2 _4011_ (.A(_0521_),
    .B(_3057_),
    .Y(_0525_));
 sky130_fd_sc_hd__buf_2 _4012_ (.A(_0525_),
    .X(_0526_));
 sky130_fd_sc_hd__clkbuf_4 _4013_ (.A(\egd_top.BitStream_buffer.BS_buffer[25] ),
    .X(_0527_));
 sky130_fd_sc_hd__clkinv_2 _4014_ (.A(_0527_),
    .Y(_0528_));
 sky130_fd_sc_hd__nand2_2 _4015_ (.A(_0521_),
    .B(_3043_),
    .Y(_0529_));
 sky130_fd_sc_hd__buf_2 _4016_ (.A(_0529_),
    .X(_0530_));
 sky130_fd_sc_hd__clkbuf_4 _4017_ (.A(\egd_top.BitStream_buffer.BS_buffer[26] ),
    .X(_0531_));
 sky130_fd_sc_hd__clkinv_2 _4018_ (.A(_0531_),
    .Y(_0532_));
 sky130_fd_sc_hd__nand2_2 _4019_ (.A(_0521_),
    .B(_3051_),
    .Y(_0533_));
 sky130_fd_sc_hd__buf_2 _4020_ (.A(_0533_),
    .X(_0534_));
 sky130_fd_sc_hd__o22a_1 _4021_ (.A1(_0528_),
    .A2(_0530_),
    .B1(_0532_),
    .B2(_0534_),
    .X(_0535_));
 sky130_fd_sc_hd__o221a_1 _4022_ (.A1(_0520_),
    .A2(_0523_),
    .B1(_0524_),
    .B2(_0526_),
    .C1(_0535_),
    .X(_0536_));
 sky130_fd_sc_hd__clkbuf_4 _4023_ (.A(\egd_top.BitStream_buffer.BS_buffer[30] ),
    .X(_0537_));
 sky130_fd_sc_hd__nor2_2 _4024_ (.A(_0488_),
    .B(_3077_),
    .Y(_0538_));
 sky130_fd_sc_hd__buf_2 _4025_ (.A(_0538_),
    .X(_0539_));
 sky130_fd_sc_hd__clkbuf_4 _4026_ (.A(\egd_top.BitStream_buffer.BS_buffer[31] ),
    .X(_0540_));
 sky130_fd_sc_hd__nor2_2 _4027_ (.A(_0488_),
    .B(_3079_),
    .Y(_0541_));
 sky130_fd_sc_hd__buf_2 _4028_ (.A(_0541_),
    .X(_0542_));
 sky130_fd_sc_hd__inv_2 _4029_ (.A(\egd_top.BitStream_buffer.BS_buffer[29] ),
    .Y(_0543_));
 sky130_fd_sc_hd__nor2_1 _4030_ (.A(_0488_),
    .B(_3072_),
    .Y(_0544_));
 sky130_fd_sc_hd__inv_2 _4031_ (.A(_0544_),
    .Y(_0545_));
 sky130_fd_sc_hd__buf_2 _4032_ (.A(_0545_),
    .X(_0546_));
 sky130_fd_sc_hd__nor2_2 _4033_ (.A(_0488_),
    .B(_3068_),
    .Y(_0547_));
 sky130_fd_sc_hd__buf_4 _4034_ (.A(_0547_),
    .X(_0548_));
 sky130_fd_sc_hd__nand2_1 _4035_ (.A(_0548_),
    .B(\egd_top.BitStream_buffer.BS_buffer[28] ),
    .Y(_0549_));
 sky130_fd_sc_hd__o21ai_1 _4036_ (.A1(_0543_),
    .A2(_0546_),
    .B1(_0549_),
    .Y(_0550_));
 sky130_fd_sc_hd__a221oi_1 _4037_ (.A1(_0537_),
    .A2(_0539_),
    .B1(_0540_),
    .B2(_0542_),
    .C1(_0550_),
    .Y(_0551_));
 sky130_fd_sc_hd__and4_1 _4038_ (.A(_0501_),
    .B(_0518_),
    .C(_0536_),
    .D(_0551_),
    .X(_0552_));
 sky130_fd_sc_hd__clkbuf_4 _4039_ (.A(\egd_top.BitStream_buffer.BS_buffer[7] ),
    .X(_0553_));
 sky130_fd_sc_hd__clkinv_2 _4040_ (.A(_0553_),
    .Y(_0554_));
 sky130_fd_sc_hd__and3_1 _4041_ (.A(_2932_),
    .B(_3211_),
    .C(_3034_),
    .X(_0555_));
 sky130_fd_sc_hd__clkbuf_4 _4042_ (.A(_0555_),
    .X(_0556_));
 sky130_fd_sc_hd__nand2_2 _4043_ (.A(_3087_),
    .B(_0556_),
    .Y(_0557_));
 sky130_fd_sc_hd__buf_2 _4044_ (.A(_0557_),
    .X(_0558_));
 sky130_fd_sc_hd__inv_2 _4045_ (.A(_0556_),
    .Y(_0559_));
 sky130_fd_sc_hd__nor2_2 _4046_ (.A(_0559_),
    .B(_3097_),
    .Y(_0560_));
 sky130_fd_sc_hd__buf_2 _4047_ (.A(_0560_),
    .X(_0561_));
 sky130_fd_sc_hd__clkbuf_4 _4048_ (.A(\egd_top.BitStream_buffer.BS_buffer[6] ),
    .X(_0562_));
 sky130_fd_sc_hd__nand2_1 _4049_ (.A(_0561_),
    .B(_0562_),
    .Y(_0563_));
 sky130_fd_sc_hd__nor2_2 _4050_ (.A(_0559_),
    .B(_3091_),
    .Y(_0564_));
 sky130_fd_sc_hd__buf_2 _4051_ (.A(_0564_),
    .X(_0565_));
 sky130_fd_sc_hd__clkbuf_4 _4052_ (.A(\egd_top.BitStream_buffer.BS_buffer[4] ),
    .X(_0566_));
 sky130_fd_sc_hd__nand2_1 _4053_ (.A(_0565_),
    .B(_0566_),
    .Y(_0567_));
 sky130_fd_sc_hd__clkbuf_4 _4054_ (.A(\egd_top.BitStream_buffer.BS_buffer[5] ),
    .X(_0568_));
 sky130_fd_sc_hd__clkinv_2 _4055_ (.A(_0568_),
    .Y(_0569_));
 sky130_fd_sc_hd__nand2_1 _4056_ (.A(_3104_),
    .B(_0556_),
    .Y(_0570_));
 sky130_fd_sc_hd__buf_2 _4057_ (.A(_0570_),
    .X(_0571_));
 sky130_fd_sc_hd__or2_1 _4058_ (.A(_0569_),
    .B(_0571_),
    .X(_0572_));
 sky130_fd_sc_hd__o2111a_1 _4059_ (.A1(_0554_),
    .A2(_0558_),
    .B1(_0563_),
    .C1(_0567_),
    .D1(_0572_),
    .X(_0573_));
 sky130_fd_sc_hd__clkinv_2 _4060_ (.A(\egd_top.BitStream_buffer.BS_buffer[11] ),
    .Y(_0574_));
 sky130_fd_sc_hd__nand2_2 _4061_ (.A(_3114_),
    .B(_0556_),
    .Y(_0575_));
 sky130_fd_sc_hd__buf_2 _4062_ (.A(_0575_),
    .X(_0576_));
 sky130_fd_sc_hd__nor2_2 _4063_ (.A(_0559_),
    .B(_3125_),
    .Y(_0577_));
 sky130_fd_sc_hd__buf_4 _4064_ (.A(_0577_),
    .X(_0578_));
 sky130_fd_sc_hd__clkbuf_4 _4065_ (.A(\egd_top.BitStream_buffer.BS_buffer[8] ),
    .X(_0579_));
 sky130_fd_sc_hd__nand2_1 _4066_ (.A(_0578_),
    .B(_0579_),
    .Y(_0580_));
 sky130_fd_sc_hd__nor2_2 _4067_ (.A(_0559_),
    .B(_3111_),
    .Y(_0581_));
 sky130_fd_sc_hd__buf_4 _4068_ (.A(_0581_),
    .X(_0582_));
 sky130_fd_sc_hd__clkbuf_4 _4069_ (.A(\egd_top.BitStream_buffer.BS_buffer[10] ),
    .X(_0583_));
 sky130_fd_sc_hd__nand2_1 _4070_ (.A(_0582_),
    .B(_0583_),
    .Y(_0584_));
 sky130_fd_sc_hd__clkbuf_4 _4071_ (.A(\egd_top.BitStream_buffer.BS_buffer[9] ),
    .X(_0585_));
 sky130_fd_sc_hd__clkinv_2 _4072_ (.A(_0585_),
    .Y(_0586_));
 sky130_fd_sc_hd__nand2_2 _4073_ (.A(_3121_),
    .B(_0556_),
    .Y(_0587_));
 sky130_fd_sc_hd__buf_2 _4074_ (.A(_0587_),
    .X(_0588_));
 sky130_fd_sc_hd__or2_1 _4075_ (.A(_0586_),
    .B(_0588_),
    .X(_0589_));
 sky130_fd_sc_hd__o2111a_1 _4076_ (.A1(_0574_),
    .A2(_0576_),
    .B1(_0580_),
    .C1(_0584_),
    .D1(_0589_),
    .X(_0590_));
 sky130_fd_sc_hd__clkinv_2 _4077_ (.A(\egd_top.BitStream_buffer.BS_buffer[2] ),
    .Y(_0591_));
 sky130_fd_sc_hd__nand2_2 _4078_ (.A(_3052_),
    .B(_0556_),
    .Y(_0592_));
 sky130_fd_sc_hd__buf_2 _4079_ (.A(_0592_),
    .X(_0593_));
 sky130_fd_sc_hd__inv_2 _4080_ (.A(\egd_top.BitStream_buffer.BS_buffer[1] ),
    .Y(_0594_));
 sky130_fd_sc_hd__nand2_1 _4081_ (.A(_3045_),
    .B(_0556_),
    .Y(_0595_));
 sky130_fd_sc_hd__buf_2 _4082_ (.A(_0595_),
    .X(_0596_));
 sky130_fd_sc_hd__clkinv_2 _4083_ (.A(\egd_top.BitStream_buffer.BS_buffer[3] ),
    .Y(_0597_));
 sky130_fd_sc_hd__nand2_1 _4084_ (.A(_3058_),
    .B(_0556_),
    .Y(_0598_));
 sky130_fd_sc_hd__clkbuf_2 _4085_ (.A(_0598_),
    .X(_0599_));
 sky130_fd_sc_hd__or2_1 _4086_ (.A(_0597_),
    .B(_0599_),
    .X(_0600_));
 sky130_fd_sc_hd__o221a_1 _4087_ (.A1(_0591_),
    .A2(_0593_),
    .B1(_0594_),
    .B2(_0596_),
    .C1(_0600_),
    .X(_0601_));
 sky130_fd_sc_hd__inv_2 _4088_ (.A(\egd_top.BitStream_buffer.BS_buffer[15] ),
    .Y(_0602_));
 sky130_fd_sc_hd__nand2_2 _4089_ (.A(_2931_),
    .B(_0556_),
    .Y(_0603_));
 sky130_fd_sc_hd__buf_2 _4090_ (.A(_0603_),
    .X(_0604_));
 sky130_fd_sc_hd__nor2_2 _4091_ (.A(_0559_),
    .B(_3068_),
    .Y(_0605_));
 sky130_fd_sc_hd__buf_2 _4092_ (.A(_0605_),
    .X(_0606_));
 sky130_fd_sc_hd__nand2_1 _4093_ (.A(_0606_),
    .B(\egd_top.BitStream_buffer.BS_buffer[12] ),
    .Y(_0607_));
 sky130_fd_sc_hd__nor2_2 _4094_ (.A(_0559_),
    .B(_3077_),
    .Y(_0608_));
 sky130_fd_sc_hd__buf_2 _4095_ (.A(_0608_),
    .X(_0609_));
 sky130_fd_sc_hd__nand2_1 _4096_ (.A(_0609_),
    .B(\egd_top.BitStream_buffer.BS_buffer[14] ),
    .Y(_0610_));
 sky130_fd_sc_hd__clkinv_2 _4097_ (.A(\egd_top.BitStream_buffer.BS_buffer[13] ),
    .Y(_0611_));
 sky130_fd_sc_hd__nand2_2 _4098_ (.A(_3071_),
    .B(_0556_),
    .Y(_0612_));
 sky130_fd_sc_hd__clkbuf_2 _4099_ (.A(_0612_),
    .X(_0613_));
 sky130_fd_sc_hd__or2_1 _4100_ (.A(_0611_),
    .B(_0613_),
    .X(_0614_));
 sky130_fd_sc_hd__o2111a_1 _4101_ (.A1(_0602_),
    .A2(_0604_),
    .B1(_0607_),
    .C1(_0610_),
    .D1(_0614_),
    .X(_0615_));
 sky130_fd_sc_hd__and4_1 _4102_ (.A(_0573_),
    .B(_0590_),
    .C(_0601_),
    .D(_0615_),
    .X(_0616_));
 sky130_fd_sc_hd__nand2_1 _4103_ (.A(_0552_),
    .B(_0616_),
    .Y(_0617_));
 sky130_fd_sc_hd__nor2_1 _4104_ (.A(_0483_),
    .B(_0617_),
    .Y(_0618_));
 sky130_fd_sc_hd__a41o_1 _4105_ (.A1(_2929_),
    .A2(_3031_),
    .A3(_3032_),
    .A4(_2921_),
    .B1(_0559_),
    .X(_0619_));
 sky130_fd_sc_hd__and4_1 _4106_ (.A(_0619_),
    .B(_2932_),
    .C(_3211_),
    .D(_3034_),
    .X(_0620_));
 sky130_fd_sc_hd__clkbuf_2 _4107_ (.A(_0620_),
    .X(_0621_));
 sky130_fd_sc_hd__buf_2 _4108_ (.A(_0621_),
    .X(_0622_));
 sky130_fd_sc_hd__clkbuf_4 _4109_ (.A(\egd_top.BitStream_buffer.BS_buffer[0] ),
    .X(_0623_));
 sky130_fd_sc_hd__nand2_1 _4110_ (.A(_0622_),
    .B(_0623_),
    .Y(_0624_));
 sky130_fd_sc_hd__nand3_1 _4111_ (.A(_0336_),
    .B(_0618_),
    .C(_0624_),
    .Y(_0625_));
 sky130_fd_sc_hd__o21a_1 _4112_ (.A1(\egd_top.BitStream_buffer.BitStream_buffer_output[15] ),
    .A2(_2964_),
    .B1(_2901_),
    .X(_0626_));
 sky130_fd_sc_hd__o21a_1 _4113_ (.A1(_3027_),
    .A2(_0625_),
    .B1(_0626_),
    .X(_0297_));
 sky130_fd_sc_hd__buf_2 _4114_ (.A(_2904_),
    .X(_0627_));
 sky130_fd_sc_hd__o21ai_1 _4115_ (.A1(\egd_top.BitStream_buffer.BitStream_buffer_output[14] ),
    .A2(_2965_),
    .B1(_0627_),
    .Y(_0628_));
 sky130_fd_sc_hd__clkinv_2 _4116_ (.A(\egd_top.BitStream_buffer.BS_buffer[40] ),
    .Y(_0629_));
 sky130_fd_sc_hd__nand2_1 _4117_ (.A(_0352_),
    .B(_0347_),
    .Y(_0630_));
 sky130_fd_sc_hd__o21ai_1 _4118_ (.A1(_0629_),
    .A2(_0349_),
    .B1(_0630_),
    .Y(_0631_));
 sky130_fd_sc_hd__a221oi_1 _4119_ (.A1(_0346_),
    .A2(_0341_),
    .B1(_0344_),
    .B2(_0354_),
    .C1(_0631_),
    .Y(_0632_));
 sky130_fd_sc_hd__inv_2 _4120_ (.A(\egd_top.BitStream_buffer.BS_buffer[34] ),
    .Y(_0633_));
 sky130_fd_sc_hd__nand2_1 _4121_ (.A(_0370_),
    .B(_0365_),
    .Y(_0634_));
 sky130_fd_sc_hd__o21ai_1 _4122_ (.A1(_0633_),
    .A2(_0367_),
    .B1(_0634_),
    .Y(_0635_));
 sky130_fd_sc_hd__a221oi_1 _4123_ (.A1(_0364_),
    .A2(_0359_),
    .B1(_0362_),
    .B2(_0337_),
    .C1(_0635_),
    .Y(_0636_));
 sky130_fd_sc_hd__clkinv_2 _4124_ (.A(\egd_top.BitStream_buffer.BS_buffer[44] ),
    .Y(_0637_));
 sky130_fd_sc_hd__nand2_1 _4125_ (.A(_0377_),
    .B(\egd_top.BitStream_buffer.BS_buffer[41] ),
    .Y(_0638_));
 sky130_fd_sc_hd__nand2_1 _4126_ (.A(_0387_),
    .B(\egd_top.BitStream_buffer.BS_buffer[43] ),
    .Y(_0639_));
 sky130_fd_sc_hd__nand2_1 _4127_ (.A(_0382_),
    .B(\egd_top.BitStream_buffer.BS_buffer[42] ),
    .Y(_0640_));
 sky130_fd_sc_hd__o2111a_1 _4128_ (.A1(_0637_),
    .A2(_0384_),
    .B1(_0638_),
    .C1(_0639_),
    .D1(_0640_),
    .X(_0641_));
 sky130_fd_sc_hd__clkbuf_4 _4129_ (.A(\egd_top.BitStream_buffer.BS_buffer[47] ),
    .X(_0642_));
 sky130_fd_sc_hd__nand2_1 _4130_ (.A(_0405_),
    .B(_0642_),
    .Y(_0643_));
 sky130_fd_sc_hd__o21ai_1 _4131_ (.A1(_0423_),
    .A2(_0402_),
    .B1(_0643_),
    .Y(_0644_));
 sky130_fd_sc_hd__a221oi_1 _4132_ (.A1(\egd_top.BitStream_buffer.BS_buffer[45] ),
    .A2(_0395_),
    .B1(_0398_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[46] ),
    .C1(_0644_),
    .Y(_0645_));
 sky130_fd_sc_hd__and4_1 _4133_ (.A(_0632_),
    .B(_0636_),
    .C(_0641_),
    .D(_0645_),
    .X(_0646_));
 sky130_fd_sc_hd__clkinv_2 _4134_ (.A(_0467_),
    .Y(_0647_));
 sky130_fd_sc_hd__nand2_1 _4135_ (.A(_0457_),
    .B(_0447_),
    .Y(_0648_));
 sky130_fd_sc_hd__nand2_1 _4136_ (.A(_0452_),
    .B(_0461_),
    .Y(_0649_));
 sky130_fd_sc_hd__inv_2 _4137_ (.A(\egd_top.BitStream_buffer.BS_buffer[58] ),
    .Y(_0650_));
 sky130_fd_sc_hd__or2_1 _4138_ (.A(_0650_),
    .B(_0463_),
    .X(_0651_));
 sky130_fd_sc_hd__o2111a_1 _4139_ (.A1(_0647_),
    .A2(_0449_),
    .B1(_0648_),
    .C1(_0649_),
    .D1(_0651_),
    .X(_0652_));
 sky130_fd_sc_hd__inv_2 _4140_ (.A(\egd_top.BitStream_buffer.BS_buffer[54] ),
    .Y(_0653_));
 sky130_fd_sc_hd__nand2_1 _4141_ (.A(_0431_),
    .B(_0436_),
    .Y(_0654_));
 sky130_fd_sc_hd__buf_2 _4142_ (.A(\egd_top.BitStream_buffer.BS_buffer[53] ),
    .X(_0655_));
 sky130_fd_sc_hd__nand2_1 _4143_ (.A(_0441_),
    .B(_0655_),
    .Y(_0656_));
 sky130_fd_sc_hd__nand2_1 _4144_ (.A(_0434_),
    .B(_0454_),
    .Y(_0657_));
 sky130_fd_sc_hd__o2111a_1 _4145_ (.A1(_0653_),
    .A2(_0438_),
    .B1(_0654_),
    .C1(_0656_),
    .D1(_0657_),
    .X(_0658_));
 sky130_fd_sc_hd__clkinv_2 _4146_ (.A(\egd_top.BitStream_buffer.BS_buffer[50] ),
    .Y(_0659_));
 sky130_fd_sc_hd__o22ai_1 _4147_ (.A1(_0420_),
    .A2(_0425_),
    .B1(_0659_),
    .B2(_0421_),
    .Y(_0660_));
 sky130_fd_sc_hd__a22o_1 _4148_ (.A1(_0416_),
    .A2(_0414_),
    .B1(_0418_),
    .B2(_0443_),
    .X(_0661_));
 sky130_fd_sc_hd__nor2_1 _4149_ (.A(_0660_),
    .B(_0661_),
    .Y(_0662_));
 sky130_fd_sc_hd__clkinv_2 _4150_ (.A(\egd_top.BitStream_buffer.BS_buffer[64] ),
    .Y(_0663_));
 sky130_fd_sc_hd__buf_2 _4151_ (.A(\egd_top.BitStream_buffer.BS_buffer[63] ),
    .X(_0664_));
 sky130_fd_sc_hd__nand2_1 _4152_ (.A(_0476_),
    .B(_0664_),
    .Y(_0665_));
 sky130_fd_sc_hd__o21ai_1 _4153_ (.A1(_0663_),
    .A2(_2935_),
    .B1(_0665_),
    .Y(_0666_));
 sky130_fd_sc_hd__a221oi_1 _4154_ (.A1(_0471_),
    .A2(_0469_),
    .B1(_0478_),
    .B2(_0473_),
    .C1(_0666_),
    .Y(_0667_));
 sky130_fd_sc_hd__and4_1 _4155_ (.A(_0652_),
    .B(_0658_),
    .C(_0662_),
    .D(_0667_),
    .X(_0668_));
 sky130_fd_sc_hd__and2_1 _4156_ (.A(_0646_),
    .B(_0668_),
    .X(_0669_));
 sky130_fd_sc_hd__clkinv_2 _4157_ (.A(\egd_top.BitStream_buffer.BS_buffer[8] ),
    .Y(_0670_));
 sky130_fd_sc_hd__nand2_1 _4158_ (.A(_0565_),
    .B(_0568_),
    .Y(_0671_));
 sky130_fd_sc_hd__nand2_1 _4159_ (.A(_0561_),
    .B(_0553_),
    .Y(_0672_));
 sky130_fd_sc_hd__clkinv_2 _4160_ (.A(\egd_top.BitStream_buffer.BS_buffer[6] ),
    .Y(_0673_));
 sky130_fd_sc_hd__or2_1 _4161_ (.A(_0673_),
    .B(_0571_),
    .X(_0674_));
 sky130_fd_sc_hd__o2111a_1 _4162_ (.A1(_0670_),
    .A2(_0558_),
    .B1(_0671_),
    .C1(_0672_),
    .D1(_0674_),
    .X(_0675_));
 sky130_fd_sc_hd__inv_2 _4163_ (.A(\egd_top.BitStream_buffer.BS_buffer[12] ),
    .Y(_0676_));
 sky130_fd_sc_hd__nand2_1 _4164_ (.A(_0578_),
    .B(_0585_),
    .Y(_0677_));
 sky130_fd_sc_hd__nand2_1 _4165_ (.A(_0582_),
    .B(\egd_top.BitStream_buffer.BS_buffer[11] ),
    .Y(_0678_));
 sky130_fd_sc_hd__clkinv_2 _4166_ (.A(_0583_),
    .Y(_0679_));
 sky130_fd_sc_hd__or2_1 _4167_ (.A(_0679_),
    .B(_0587_),
    .X(_0680_));
 sky130_fd_sc_hd__o2111a_1 _4168_ (.A1(_0676_),
    .A2(_0576_),
    .B1(_0677_),
    .C1(_0678_),
    .D1(_0680_),
    .X(_0681_));
 sky130_fd_sc_hd__clkinv_2 _4169_ (.A(\egd_top.BitStream_buffer.BS_buffer[4] ),
    .Y(_0682_));
 sky130_fd_sc_hd__or2_1 _4170_ (.A(_0591_),
    .B(_0595_),
    .X(_0683_));
 sky130_fd_sc_hd__o221a_1 _4171_ (.A1(_0597_),
    .A2(_0593_),
    .B1(_0682_),
    .B2(_0599_),
    .C1(_0683_),
    .X(_0684_));
 sky130_fd_sc_hd__clkinv_2 _4172_ (.A(\egd_top.BitStream_buffer.BS_buffer[16] ),
    .Y(_0685_));
 sky130_fd_sc_hd__nand2_1 _4173_ (.A(_0609_),
    .B(\egd_top.BitStream_buffer.BS_buffer[15] ),
    .Y(_0686_));
 sky130_fd_sc_hd__nand2_1 _4174_ (.A(_0606_),
    .B(\egd_top.BitStream_buffer.BS_buffer[13] ),
    .Y(_0687_));
 sky130_fd_sc_hd__inv_2 _4175_ (.A(\egd_top.BitStream_buffer.BS_buffer[14] ),
    .Y(_0688_));
 sky130_fd_sc_hd__or2_1 _4176_ (.A(_0688_),
    .B(_0613_),
    .X(_0689_));
 sky130_fd_sc_hd__o2111a_1 _4177_ (.A1(_0685_),
    .A2(_0604_),
    .B1(_0686_),
    .C1(_0687_),
    .D1(_0689_),
    .X(_0690_));
 sky130_fd_sc_hd__and4_1 _4178_ (.A(_0675_),
    .B(_0681_),
    .C(_0684_),
    .D(_0690_),
    .X(_0691_));
 sky130_fd_sc_hd__clkinv_2 _4179_ (.A(_0498_),
    .Y(_0692_));
 sky130_fd_sc_hd__nand2_1 _4180_ (.A(_0497_),
    .B(_0502_),
    .Y(_0693_));
 sky130_fd_sc_hd__o21ai_1 _4181_ (.A1(_0692_),
    .A2(_0495_),
    .B1(_0693_),
    .Y(_0694_));
 sky130_fd_sc_hd__a221oi_1 _4182_ (.A1(\egd_top.BitStream_buffer.BS_buffer[17] ),
    .A2(_0487_),
    .B1(_0491_),
    .B2(_0490_),
    .C1(_0694_),
    .Y(_0695_));
 sky130_fd_sc_hd__nand2_1 _4183_ (.A(_0514_),
    .B(_0509_),
    .Y(_0696_));
 sky130_fd_sc_hd__o21ai_1 _4184_ (.A1(_0520_),
    .A2(_0512_),
    .B1(_0696_),
    .Y(_0697_));
 sky130_fd_sc_hd__a221oi_1 _4185_ (.A1(_0505_),
    .A2(_0504_),
    .B1(_0515_),
    .B2(_0508_),
    .C1(_0697_),
    .Y(_0698_));
 sky130_fd_sc_hd__inv_2 _4186_ (.A(\egd_top.BitStream_buffer.BS_buffer[28] ),
    .Y(_0699_));
 sky130_fd_sc_hd__o22a_1 _4187_ (.A1(_0532_),
    .A2(_0530_),
    .B1(_0524_),
    .B2(_0533_),
    .X(_0700_));
 sky130_fd_sc_hd__o221a_1 _4188_ (.A1(_0528_),
    .A2(_0523_),
    .B1(_0699_),
    .B2(_0526_),
    .C1(_0700_),
    .X(_0701_));
 sky130_fd_sc_hd__clkinv_2 _4189_ (.A(_0537_),
    .Y(_0702_));
 sky130_fd_sc_hd__nand2_1 _4190_ (.A(_0548_),
    .B(\egd_top.BitStream_buffer.BS_buffer[29] ),
    .Y(_0703_));
 sky130_fd_sc_hd__o21ai_1 _4191_ (.A1(_0702_),
    .A2(_0546_),
    .B1(_0703_),
    .Y(_0704_));
 sky130_fd_sc_hd__a221oi_1 _4192_ (.A1(_0540_),
    .A2(_0539_),
    .B1(\egd_top.BitStream_buffer.BS_buffer[32] ),
    .B2(_0542_),
    .C1(_0704_),
    .Y(_0705_));
 sky130_fd_sc_hd__and4_1 _4193_ (.A(_0695_),
    .B(_0698_),
    .C(_0701_),
    .D(_0705_),
    .X(_0706_));
 sky130_fd_sc_hd__and3_1 _4194_ (.A(_0669_),
    .B(_0691_),
    .C(_0706_),
    .X(_0707_));
 sky130_fd_sc_hd__clkbuf_4 _4195_ (.A(\egd_top.BitStream_buffer.BS_buffer[98] ),
    .X(_0708_));
 sky130_fd_sc_hd__clkinv_2 _4196_ (.A(\egd_top.BitStream_buffer.BS_buffer[99] ),
    .Y(_0709_));
 sky130_fd_sc_hd__nand2_1 _4197_ (.A(_3061_),
    .B(_3094_),
    .Y(_0710_));
 sky130_fd_sc_hd__o21ai_1 _4198_ (.A1(_0709_),
    .A2(_3056_),
    .B1(_0710_),
    .Y(_0711_));
 sky130_fd_sc_hd__a221oi_1 _4199_ (.A1(_3040_),
    .A2(_3039_),
    .B1(_0708_),
    .B2(_3048_),
    .C1(_0711_),
    .Y(_0712_));
 sky130_fd_sc_hd__inv_2 _4200_ (.A(\egd_top.BitStream_buffer.BS_buffer[102] ),
    .Y(_0713_));
 sky130_fd_sc_hd__clkbuf_4 _4201_ (.A(\egd_top.BitStream_buffer.BS_buffer[103] ),
    .X(_0714_));
 sky130_fd_sc_hd__nand2_1 _4202_ (.A(_3099_),
    .B(_0714_),
    .Y(_0715_));
 sky130_fd_sc_hd__buf_2 _4203_ (.A(\egd_top.BitStream_buffer.BS_buffer[101] ),
    .X(_0716_));
 sky130_fd_sc_hd__nand2_1 _4204_ (.A(_3093_),
    .B(_0716_),
    .Y(_0717_));
 sky130_fd_sc_hd__inv_2 _4205_ (.A(\egd_top.BitStream_buffer.BS_buffer[104] ),
    .Y(_0718_));
 sky130_fd_sc_hd__or2_1 _4206_ (.A(_0718_),
    .B(_3088_),
    .X(_0719_));
 sky130_fd_sc_hd__o2111a_1 _4207_ (.A1(_0713_),
    .A2(_3106_),
    .B1(_0715_),
    .C1(_0717_),
    .D1(_0719_),
    .X(_0720_));
 sky130_fd_sc_hd__clkinv_2 _4208_ (.A(\egd_top.BitStream_buffer.BS_buffer[106] ),
    .Y(_0721_));
 sky130_fd_sc_hd__clkbuf_4 _4209_ (.A(\egd_top.BitStream_buffer.BS_buffer[105] ),
    .X(_0722_));
 sky130_fd_sc_hd__nand2_1 _4210_ (.A(_3127_),
    .B(_0722_),
    .Y(_0723_));
 sky130_fd_sc_hd__o21ai_1 _4211_ (.A1(_0721_),
    .A2(_3123_),
    .B1(_0723_),
    .Y(_0724_));
 sky130_fd_sc_hd__a221oi_1 _4212_ (.A1(_3118_),
    .A2(_3113_),
    .B1(_3117_),
    .B2(_3066_),
    .C1(_0724_),
    .Y(_0725_));
 sky130_fd_sc_hd__buf_2 _4213_ (.A(_3078_),
    .X(_0726_));
 sky130_fd_sc_hd__clkinv_2 _4214_ (.A(\egd_top.BitStream_buffer.BS_buffer[109] ),
    .Y(_0727_));
 sky130_fd_sc_hd__inv_2 _4215_ (.A(_3069_),
    .Y(_0728_));
 sky130_fd_sc_hd__clkbuf_4 _4216_ (.A(_0728_),
    .X(_0729_));
 sky130_fd_sc_hd__nand2_1 _4217_ (.A(_3074_),
    .B(_3075_),
    .Y(_0730_));
 sky130_fd_sc_hd__o21ai_1 _4218_ (.A1(_0727_),
    .A2(_0729_),
    .B1(_0730_),
    .Y(_0731_));
 sky130_fd_sc_hd__a221oi_1 _4219_ (.A1(_3169_),
    .A2(_3081_),
    .B1(_3082_),
    .B2(_0726_),
    .C1(_0731_),
    .Y(_0732_));
 sky130_fd_sc_hd__and4_1 _4220_ (.A(_0712_),
    .B(_0720_),
    .C(_0725_),
    .D(_0732_),
    .X(_0733_));
 sky130_fd_sc_hd__nand2_1 _4221_ (.A(_3148_),
    .B(_3133_),
    .Y(_0734_));
 sky130_fd_sc_hd__o21ai_1 _4222_ (.A1(_3006_),
    .A2(_3145_),
    .B1(_0734_),
    .Y(_0735_));
 sky130_fd_sc_hd__a221oi_2 _4223_ (.A1(_3138_),
    .A2(_3137_),
    .B1(_3173_),
    .B2(_3141_),
    .C1(_0735_),
    .Y(_0736_));
 sky130_fd_sc_hd__nand2_1 _4224_ (.A(_3163_),
    .B(_3153_),
    .Y(_0737_));
 sky130_fd_sc_hd__nand2_1 _4225_ (.A(_3168_),
    .B(_3164_),
    .Y(_0738_));
 sky130_fd_sc_hd__nand2_1 _4226_ (.A(_0737_),
    .B(_0738_),
    .Y(_0739_));
 sky130_fd_sc_hd__a221oi_1 _4227_ (.A1(_3157_),
    .A2(_3156_),
    .B1(_3204_),
    .B2(_3160_),
    .C1(_0739_),
    .Y(_0740_));
 sky130_fd_sc_hd__clkbuf_4 _4228_ (.A(\egd_top.BitStream_buffer.BS_buffer[126] ),
    .X(_0741_));
 sky130_fd_sc_hd__a22o_1 _4229_ (.A1(_3181_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[127] ),
    .B1(\egd_top.BitStream_buffer.BS_buffer[125] ),
    .B2(_3175_),
    .X(_0742_));
 sky130_fd_sc_hd__a221oi_4 _4230_ (.A1(_0741_),
    .A2(_3180_),
    .B1(_0623_),
    .B2(_3186_),
    .C1(_0742_),
    .Y(_0743_));
 sky130_fd_sc_hd__clkbuf_4 _4231_ (.A(\egd_top.BitStream_buffer.BS_buffer[120] ),
    .X(_0744_));
 sky130_fd_sc_hd__a22o_1 _4232_ (.A1(_3198_),
    .A2(_3193_),
    .B1(_3196_),
    .B2(_0744_),
    .X(_0745_));
 sky130_fd_sc_hd__clkbuf_4 _4233_ (.A(\egd_top.BitStream_buffer.BS_buffer[117] ),
    .X(_0746_));
 sky130_fd_sc_hd__a32o_1 _4234_ (.A1(_3104_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[118] ),
    .A3(_3142_),
    .B1(_0746_),
    .B2(_3202_),
    .X(_0747_));
 sky130_fd_sc_hd__nor2_1 _4235_ (.A(_0745_),
    .B(_0747_),
    .Y(_0748_));
 sky130_fd_sc_hd__and4_1 _4236_ (.A(_0736_),
    .B(_0740_),
    .C(_0743_),
    .D(_0748_),
    .X(_0749_));
 sky130_fd_sc_hd__nand2_1 _4237_ (.A(_0733_),
    .B(_0749_),
    .Y(_0750_));
 sky130_fd_sc_hd__clkbuf_4 _4238_ (.A(\egd_top.BitStream_buffer.BS_buffer[65] ),
    .X(_0751_));
 sky130_fd_sc_hd__inv_2 _4239_ (.A(_3239_),
    .Y(_0752_));
 sky130_fd_sc_hd__a22o_1 _4240_ (.A1(_0751_),
    .A2(_3243_),
    .B1(_0752_),
    .B2(_3230_),
    .X(_0753_));
 sky130_fd_sc_hd__a221oi_1 _4241_ (.A1(_3237_),
    .A2(_3233_),
    .B1(_3210_),
    .B2(_3236_),
    .C1(_0753_),
    .Y(_0754_));
 sky130_fd_sc_hd__inv_2 _4242_ (.A(\egd_top.BitStream_buffer.BS_buffer[70] ),
    .Y(_0755_));
 sky130_fd_sc_hd__nand2_1 _4243_ (.A(_3216_),
    .B(_3217_),
    .Y(_0756_));
 sky130_fd_sc_hd__o21ai_1 _4244_ (.A1(_0755_),
    .A2(_3218_),
    .B1(_0756_),
    .Y(_0757_));
 sky130_fd_sc_hd__a221oi_1 _4245_ (.A1(_3227_),
    .A2(_3224_),
    .B1(_3256_),
    .B2(_3226_),
    .C1(_0757_),
    .Y(_0758_));
 sky130_fd_sc_hd__clkinv_2 _4246_ (.A(\egd_top.BitStream_buffer.BS_buffer[73] ),
    .Y(_0759_));
 sky130_fd_sc_hd__nand2_1 _4247_ (.A(_3263_),
    .B(_3248_),
    .Y(_0760_));
 sky130_fd_sc_hd__o21ai_1 _4248_ (.A1(_0759_),
    .A2(_3260_),
    .B1(_0760_),
    .Y(_0761_));
 sky130_fd_sc_hd__a221oi_1 _4249_ (.A1(_3252_),
    .A2(_3251_),
    .B1(_3268_),
    .B2(_3255_),
    .C1(_0761_),
    .Y(_0762_));
 sky130_fd_sc_hd__nand2_1 _4250_ (.A(_3282_),
    .B(_3276_),
    .Y(_0763_));
 sky130_fd_sc_hd__o21ai_1 _4251_ (.A1(_3296_),
    .A2(_3279_),
    .B1(_0763_),
    .Y(_0764_));
 sky130_fd_sc_hd__a221oi_1 _4252_ (.A1(_3272_),
    .A2(_3271_),
    .B1(_3283_),
    .B2(_3275_),
    .C1(_0764_),
    .Y(_0765_));
 sky130_fd_sc_hd__and4_1 _4253_ (.A(_0754_),
    .B(_0758_),
    .C(_0762_),
    .D(_0765_),
    .X(_0766_));
 sky130_fd_sc_hd__clkinv_2 _4254_ (.A(\egd_top.BitStream_buffer.BS_buffer[81] ),
    .Y(_0767_));
 sky130_fd_sc_hd__nand2_1 _4255_ (.A(_3301_),
    .B(_3288_),
    .Y(_0768_));
 sky130_fd_sc_hd__o21ai_1 _4256_ (.A1(_0767_),
    .A2(_3299_),
    .B1(_0768_),
    .Y(_0769_));
 sky130_fd_sc_hd__a221oi_1 _4257_ (.A1(_3293_),
    .A2(_3292_),
    .B1(_3315_),
    .B2(_3295_),
    .C1(_0769_),
    .Y(_0770_));
 sky130_fd_sc_hd__clkinv_2 _4258_ (.A(\egd_top.BitStream_buffer.BS_buffer[86] ),
    .Y(_0771_));
 sky130_fd_sc_hd__buf_2 _4259_ (.A(\egd_top.BitStream_buffer.BS_buffer[87] ),
    .X(_0772_));
 sky130_fd_sc_hd__nand2_1 _4260_ (.A(_3310_),
    .B(_0772_),
    .Y(_0773_));
 sky130_fd_sc_hd__buf_2 _4261_ (.A(\egd_top.BitStream_buffer.BS_buffer[85] ),
    .X(_0774_));
 sky130_fd_sc_hd__nand2_1 _4262_ (.A(_3314_),
    .B(_0774_),
    .Y(_0775_));
 sky130_fd_sc_hd__inv_2 _4263_ (.A(\egd_top.BitStream_buffer.BS_buffer[88] ),
    .Y(_0776_));
 sky130_fd_sc_hd__or2_1 _4264_ (.A(_0776_),
    .B(_3307_),
    .X(_0777_));
 sky130_fd_sc_hd__o2111a_1 _4265_ (.A1(_0771_),
    .A2(_3319_),
    .B1(_0773_),
    .C1(_0775_),
    .D1(_0777_),
    .X(_0778_));
 sky130_fd_sc_hd__clkinv_2 _4266_ (.A(\egd_top.BitStream_buffer.BS_buffer[90] ),
    .Y(_0779_));
 sky130_fd_sc_hd__clkbuf_4 _4267_ (.A(\egd_top.BitStream_buffer.BS_buffer[89] ),
    .X(_0780_));
 sky130_fd_sc_hd__nand2_1 _4268_ (.A(_3333_),
    .B(_0780_),
    .Y(_0781_));
 sky130_fd_sc_hd__o21ai_1 _4269_ (.A1(_0779_),
    .A2(_3330_),
    .B1(_0781_),
    .Y(_0782_));
 sky130_fd_sc_hd__a221oi_1 _4270_ (.A1(_3327_),
    .A2(_3324_),
    .B1(_3326_),
    .B2(_0330_),
    .C1(_0782_),
    .Y(_0783_));
 sky130_fd_sc_hd__clkinv_2 _4271_ (.A(\egd_top.BitStream_buffer.BS_buffer[94] ),
    .Y(_0784_));
 sky130_fd_sc_hd__clkbuf_4 _4272_ (.A(\egd_top.BitStream_buffer.BS_buffer[93] ),
    .X(_0785_));
 sky130_fd_sc_hd__nand2_1 _4273_ (.A(_0329_),
    .B(_0785_),
    .Y(_0786_));
 sky130_fd_sc_hd__o21ai_1 _4274_ (.A1(_0784_),
    .A2(_0327_),
    .B1(_0786_),
    .Y(_0787_));
 sky130_fd_sc_hd__a221oi_1 _4275_ (.A1(_3028_),
    .A2(_0323_),
    .B1(_3341_),
    .B2(_3340_),
    .C1(_0787_),
    .Y(_0788_));
 sky130_fd_sc_hd__and4_1 _4276_ (.A(_0770_),
    .B(_0778_),
    .C(_0783_),
    .D(_0788_),
    .X(_0789_));
 sky130_fd_sc_hd__nand2_1 _4277_ (.A(_0766_),
    .B(_0789_),
    .Y(_0790_));
 sky130_fd_sc_hd__nor2_1 _4278_ (.A(_0750_),
    .B(_0790_),
    .Y(_0791_));
 sky130_fd_sc_hd__clkbuf_4 _4279_ (.A(\egd_top.BitStream_buffer.BS_buffer[1] ),
    .X(_0792_));
 sky130_fd_sc_hd__nand2_1 _4280_ (.A(_0622_),
    .B(_0792_),
    .Y(_0793_));
 sky130_fd_sc_hd__nand3_1 _4281_ (.A(_0707_),
    .B(_0791_),
    .C(_0793_),
    .Y(_0794_));
 sky130_fd_sc_hd__nor2_1 _4282_ (.A(_3027_),
    .B(_0794_),
    .Y(_0795_));
 sky130_fd_sc_hd__nor2_1 _4283_ (.A(_0628_),
    .B(_0795_),
    .Y(_0296_));
 sky130_fd_sc_hd__clkinv_2 _4284_ (.A(\egd_top.BitStream_buffer.BS_buffer[100] ),
    .Y(_0796_));
 sky130_fd_sc_hd__nand2_1 _4285_ (.A(_3061_),
    .B(_0716_),
    .Y(_0797_));
 sky130_fd_sc_hd__o21ai_1 _4286_ (.A1(_0796_),
    .A2(_3056_),
    .B1(_0797_),
    .Y(_0798_));
 sky130_fd_sc_hd__a221oi_1 _4287_ (.A1(_0708_),
    .A2(_3039_),
    .B1(_3062_),
    .B2(_3048_),
    .C1(_0798_),
    .Y(_0799_));
 sky130_fd_sc_hd__nand2_1 _4288_ (.A(_3093_),
    .B(_3100_),
    .Y(_0800_));
 sky130_fd_sc_hd__nand2_1 _4289_ (.A(_3099_),
    .B(_3128_),
    .Y(_0801_));
 sky130_fd_sc_hd__or2_1 _4290_ (.A(_3085_),
    .B(_3106_),
    .X(_0802_));
 sky130_fd_sc_hd__o2111a_1 _4291_ (.A1(_3119_),
    .A2(_3089_),
    .B1(_0800_),
    .C1(_0801_),
    .D1(_0802_),
    .X(_0803_));
 sky130_fd_sc_hd__clkinv_2 _4292_ (.A(\egd_top.BitStream_buffer.BS_buffer[107] ),
    .Y(_0804_));
 sky130_fd_sc_hd__nand2_1 _4293_ (.A(_3127_),
    .B(_3109_),
    .Y(_0805_));
 sky130_fd_sc_hd__o21ai_1 _4294_ (.A1(_0804_),
    .A2(_3123_),
    .B1(_0805_),
    .Y(_0806_));
 sky130_fd_sc_hd__a221oi_1 _4295_ (.A1(_3066_),
    .A2(_3113_),
    .B1(_3117_),
    .B2(_3070_),
    .C1(_0806_),
    .Y(_0807_));
 sky130_fd_sc_hd__clkinv_2 _4296_ (.A(\egd_top.BitStream_buffer.BS_buffer[110] ),
    .Y(_0808_));
 sky130_fd_sc_hd__nand2_1 _4297_ (.A(_3074_),
    .B(_3082_),
    .Y(_0809_));
 sky130_fd_sc_hd__o21ai_1 _4298_ (.A1(_0808_),
    .A2(_0729_),
    .B1(_0809_),
    .Y(_0810_));
 sky130_fd_sc_hd__a221oi_1 _4299_ (.A1(_3169_),
    .A2(_0726_),
    .B1(_3164_),
    .B2(_3081_),
    .C1(_0810_),
    .Y(_0811_));
 sky130_fd_sc_hd__and4_1 _4300_ (.A(_0799_),
    .B(_0803_),
    .C(_0807_),
    .D(_0811_),
    .X(_0812_));
 sky130_fd_sc_hd__nand2_1 _4301_ (.A(_3148_),
    .B(_3138_),
    .Y(_0813_));
 sky130_fd_sc_hd__o21ai_1 _4302_ (.A1(_3009_),
    .A2(_3145_),
    .B1(_0813_),
    .Y(_0814_));
 sky130_fd_sc_hd__a221oi_1 _4303_ (.A1(_3173_),
    .A2(_3137_),
    .B1(_3177_),
    .B2(_3141_),
    .C1(_0814_),
    .Y(_0815_));
 sky130_fd_sc_hd__nand2_1 _4304_ (.A(_3163_),
    .B(_3157_),
    .Y(_0816_));
 sky130_fd_sc_hd__nand2_1 _4305_ (.A(_3168_),
    .B(_3153_),
    .Y(_0817_));
 sky130_fd_sc_hd__nand2_1 _4306_ (.A(_0816_),
    .B(_0817_),
    .Y(_0818_));
 sky130_fd_sc_hd__a221oi_2 _4307_ (.A1(_3204_),
    .A2(_3156_),
    .B1(_0746_),
    .B2(_3160_),
    .C1(_0818_),
    .Y(_0819_));
 sky130_fd_sc_hd__a22o_1 _4308_ (.A1(_3181_),
    .A2(_0623_),
    .B1(_0741_),
    .B2(_3176_),
    .X(_0820_));
 sky130_fd_sc_hd__a221oi_1 _4309_ (.A1(_3187_),
    .A2(_3180_),
    .B1(_0792_),
    .B2(_3186_),
    .C1(_0820_),
    .Y(_0821_));
 sky130_fd_sc_hd__nand2_1 _4310_ (.A(_3203_),
    .B(_3191_),
    .Y(_0822_));
 sky130_fd_sc_hd__o21ai_1 _4311_ (.A1(_2999_),
    .A2(_3200_),
    .B1(_0822_),
    .Y(_0823_));
 sky130_fd_sc_hd__a221oi_1 _4312_ (.A1(_0744_),
    .A2(_3194_),
    .B1(_3197_),
    .B2(_3149_),
    .C1(_0823_),
    .Y(_0824_));
 sky130_fd_sc_hd__and4_1 _4313_ (.A(_0815_),
    .B(_0819_),
    .C(_0821_),
    .D(_0824_),
    .X(_0825_));
 sky130_fd_sc_hd__nand2_1 _4314_ (.A(_0812_),
    .B(_0825_),
    .Y(_0826_));
 sky130_fd_sc_hd__a22o_1 _4315_ (.A1(_3256_),
    .A2(_3224_),
    .B1(_3226_),
    .B2(_3264_),
    .X(_0827_));
 sky130_fd_sc_hd__a221oi_1 _4316_ (.A1(_3221_),
    .A2(_3216_),
    .B1(_3227_),
    .B2(_3220_),
    .C1(_0827_),
    .Y(_0828_));
 sky130_fd_sc_hd__clkinv_2 _4317_ (.A(\egd_top.BitStream_buffer.BS_buffer[67] ),
    .Y(_0829_));
 sky130_fd_sc_hd__nand2_1 _4318_ (.A(_3243_),
    .B(_3230_),
    .Y(_0830_));
 sky130_fd_sc_hd__o21ai_1 _4319_ (.A1(_0829_),
    .A2(_3240_),
    .B1(_0830_),
    .Y(_0831_));
 sky130_fd_sc_hd__a221oi_1 _4320_ (.A1(_3210_),
    .A2(_3233_),
    .B1(_3236_),
    .B2(_3217_),
    .C1(_0831_),
    .Y(_0832_));
 sky130_fd_sc_hd__inv_2 _4321_ (.A(\egd_top.BitStream_buffer.BS_buffer[74] ),
    .Y(_0833_));
 sky130_fd_sc_hd__nand2_1 _4322_ (.A(_3263_),
    .B(_3252_),
    .Y(_0834_));
 sky130_fd_sc_hd__o21ai_1 _4323_ (.A1(_0833_),
    .A2(_3260_),
    .B1(_0834_),
    .Y(_0835_));
 sky130_fd_sc_hd__a221oi_1 _4324_ (.A1(_3268_),
    .A2(_3251_),
    .B1(_3272_),
    .B2(_3255_),
    .C1(_0835_),
    .Y(_0836_));
 sky130_fd_sc_hd__buf_2 _4325_ (.A(\egd_top.BitStream_buffer.BS_buffer[80] ),
    .X(_0837_));
 sky130_fd_sc_hd__nand2_1 _4326_ (.A(_3282_),
    .B(_0837_),
    .Y(_0838_));
 sky130_fd_sc_hd__o21ai_1 _4327_ (.A1(_0767_),
    .A2(_3279_),
    .B1(_0838_),
    .Y(_0839_));
 sky130_fd_sc_hd__a221oi_1 _4328_ (.A1(_3283_),
    .A2(_3271_),
    .B1(_3276_),
    .B2(_3275_),
    .C1(_0839_),
    .Y(_0840_));
 sky130_fd_sc_hd__and4_1 _4329_ (.A(_0828_),
    .B(_0832_),
    .C(_0836_),
    .D(_0840_),
    .X(_0841_));
 sky130_fd_sc_hd__clkinv_2 _4330_ (.A(\egd_top.BitStream_buffer.BS_buffer[82] ),
    .Y(_0842_));
 sky130_fd_sc_hd__nand2_1 _4331_ (.A(_3301_),
    .B(_3293_),
    .Y(_0843_));
 sky130_fd_sc_hd__o21ai_1 _4332_ (.A1(_0842_),
    .A2(_3299_),
    .B1(_0843_),
    .Y(_0844_));
 sky130_fd_sc_hd__a221oi_1 _4333_ (.A1(_3315_),
    .A2(_3292_),
    .B1(_0774_),
    .B2(_3295_),
    .C1(_0844_),
    .Y(_0845_));
 sky130_fd_sc_hd__nand2_1 _4334_ (.A(_3310_),
    .B(_3334_),
    .Y(_0846_));
 sky130_fd_sc_hd__nand2_1 _4335_ (.A(_3314_),
    .B(_3311_),
    .Y(_0847_));
 sky130_fd_sc_hd__or2_1 _4336_ (.A(_3306_),
    .B(_3319_),
    .X(_0848_));
 sky130_fd_sc_hd__o2111a_1 _4337_ (.A1(_3328_),
    .A2(_3308_),
    .B1(_0846_),
    .C1(_0847_),
    .D1(_0848_),
    .X(_0849_));
 sky130_fd_sc_hd__clkinv_2 _4338_ (.A(\egd_top.BitStream_buffer.BS_buffer[91] ),
    .Y(_0850_));
 sky130_fd_sc_hd__nand2_1 _4339_ (.A(_3333_),
    .B(_3322_),
    .Y(_0851_));
 sky130_fd_sc_hd__o21ai_1 _4340_ (.A1(_0850_),
    .A2(_3330_),
    .B1(_0851_),
    .Y(_0852_));
 sky130_fd_sc_hd__a221oi_1 _4341_ (.A1(_0330_),
    .A2(_3324_),
    .B1(_3326_),
    .B2(_0785_),
    .C1(_0852_),
    .Y(_0853_));
 sky130_fd_sc_hd__inv_2 _4342_ (.A(\egd_top.BitStream_buffer.BS_buffer[95] ),
    .Y(_0854_));
 sky130_fd_sc_hd__nand2_1 _4343_ (.A(_0329_),
    .B(_3338_),
    .Y(_0855_));
 sky130_fd_sc_hd__o21ai_1 _4344_ (.A1(_0854_),
    .A2(_0327_),
    .B1(_0855_),
    .Y(_0856_));
 sky130_fd_sc_hd__a221oi_1 _4345_ (.A1(_3028_),
    .A2(_3340_),
    .B1(_3040_),
    .B2(_0323_),
    .C1(_0856_),
    .Y(_0857_));
 sky130_fd_sc_hd__and4_1 _4346_ (.A(_0845_),
    .B(_0849_),
    .C(_0853_),
    .D(_0857_),
    .X(_0858_));
 sky130_fd_sc_hd__nand2_2 _4347_ (.A(_0841_),
    .B(_0858_),
    .Y(_0859_));
 sky130_fd_sc_hd__nor2_1 _4348_ (.A(_0826_),
    .B(_0859_),
    .Y(_0860_));
 sky130_fd_sc_hd__clkinv_2 _4349_ (.A(\egd_top.BitStream_buffer.BS_buffer[41] ),
    .Y(_0861_));
 sky130_fd_sc_hd__nand2_1 _4350_ (.A(_0353_),
    .B(_0375_),
    .Y(_0862_));
 sky130_fd_sc_hd__o21ai_1 _4351_ (.A1(_0861_),
    .A2(_0350_),
    .B1(_0862_),
    .Y(_0863_));
 sky130_fd_sc_hd__a221oi_1 _4352_ (.A1(_0354_),
    .A2(_0342_),
    .B1(_0345_),
    .B2(_0347_),
    .C1(_0863_),
    .Y(_0864_));
 sky130_fd_sc_hd__clkinv_2 _4353_ (.A(_0364_),
    .Y(_0865_));
 sky130_fd_sc_hd__nand2_1 _4354_ (.A(_0371_),
    .B(\egd_top.BitStream_buffer.BS_buffer[34] ),
    .Y(_0866_));
 sky130_fd_sc_hd__o21ai_1 _4355_ (.A1(_0865_),
    .A2(_0368_),
    .B1(_0866_),
    .Y(_0867_));
 sky130_fd_sc_hd__a221oi_1 _4356_ (.A1(_0337_),
    .A2(_0360_),
    .B1(_0363_),
    .B2(_0346_),
    .C1(_0867_),
    .Y(_0868_));
 sky130_fd_sc_hd__clkbuf_4 _4357_ (.A(\egd_top.BitStream_buffer.BS_buffer[43] ),
    .X(_0869_));
 sky130_fd_sc_hd__inv_2 _4358_ (.A(\egd_top.BitStream_buffer.BS_buffer[45] ),
    .Y(_0870_));
 sky130_fd_sc_hd__nand2_1 _4359_ (.A(_0388_),
    .B(_0393_),
    .Y(_0871_));
 sky130_fd_sc_hd__o21ai_1 _4360_ (.A1(_0870_),
    .A2(_0385_),
    .B1(_0871_),
    .Y(_0872_));
 sky130_fd_sc_hd__a221oi_1 _4361_ (.A1(_0389_),
    .A2(_0378_),
    .B1(_0869_),
    .B2(_0382_),
    .C1(_0872_),
    .Y(_0873_));
 sky130_fd_sc_hd__buf_2 _4362_ (.A(\egd_top.BitStream_buffer.BS_buffer[48] ),
    .X(_0874_));
 sky130_fd_sc_hd__nand2_1 _4363_ (.A(_0406_),
    .B(_0874_),
    .Y(_0875_));
 sky130_fd_sc_hd__o21ai_1 _4364_ (.A1(_0420_),
    .A2(_0403_),
    .B1(_0875_),
    .Y(_0876_));
 sky130_fd_sc_hd__a221oi_1 _4365_ (.A1(_0407_),
    .A2(_0396_),
    .B1(_0399_),
    .B2(_0642_),
    .C1(_0876_),
    .Y(_0877_));
 sky130_fd_sc_hd__and4_1 _4366_ (.A(_0864_),
    .B(_0868_),
    .C(_0873_),
    .D(_0877_),
    .X(_0878_));
 sky130_fd_sc_hd__clkinv_2 _4367_ (.A(\egd_top.BitStream_buffer.BS_buffer[51] ),
    .Y(_0879_));
 sky130_fd_sc_hd__or2_1 _4368_ (.A(_0659_),
    .B(_0425_),
    .X(_0880_));
 sky130_fd_sc_hd__o21ai_1 _4369_ (.A1(_0879_),
    .A2(_0422_),
    .B1(_0880_),
    .Y(_0881_));
 sky130_fd_sc_hd__a221oi_1 _4370_ (.A1(_0443_),
    .A2(_0415_),
    .B1(_0655_),
    .B2(_0419_),
    .C1(_0881_),
    .Y(_0882_));
 sky130_fd_sc_hd__clkinv_2 _4371_ (.A(_0436_),
    .Y(_0883_));
 sky130_fd_sc_hd__nand2_1 _4372_ (.A(_0442_),
    .B(_0429_),
    .Y(_0884_));
 sky130_fd_sc_hd__o21ai_1 _4373_ (.A1(_0883_),
    .A2(_0439_),
    .B1(_0884_),
    .Y(_0885_));
 sky130_fd_sc_hd__a221oi_1 _4374_ (.A1(_0454_),
    .A2(_0432_),
    .B1(_0435_),
    .B2(_0461_),
    .C1(_0885_),
    .Y(_0886_));
 sky130_fd_sc_hd__clkinv_2 _4375_ (.A(_0471_),
    .Y(_0887_));
 sky130_fd_sc_hd__nand2_1 _4376_ (.A(_0453_),
    .B(_0459_),
    .Y(_0888_));
 sky130_fd_sc_hd__nand2_1 _4377_ (.A(_0458_),
    .B(_0467_),
    .Y(_0889_));
 sky130_fd_sc_hd__or2_1 _4378_ (.A(_0448_),
    .B(_0464_),
    .X(_0890_));
 sky130_fd_sc_hd__o2111a_1 _4379_ (.A1(_0887_),
    .A2(_0450_),
    .B1(_0888_),
    .C1(_0889_),
    .D1(_0890_),
    .X(_0891_));
 sky130_fd_sc_hd__nand2_1 _4380_ (.A(_0477_),
    .B(_3244_),
    .Y(_0892_));
 sky130_fd_sc_hd__o21ai_1 _4381_ (.A1(_3238_),
    .A2(_2935_),
    .B1(_0892_),
    .Y(_0893_));
 sky130_fd_sc_hd__a221oi_1 _4382_ (.A1(_0478_),
    .A2(_0470_),
    .B1(_0664_),
    .B2(_0473_),
    .C1(_0893_),
    .Y(_0894_));
 sky130_fd_sc_hd__and4_1 _4383_ (.A(_0882_),
    .B(_0886_),
    .C(_0891_),
    .D(_0894_),
    .X(_0895_));
 sky130_fd_sc_hd__nand2_1 _4384_ (.A(_0878_),
    .B(_0895_),
    .Y(_0896_));
 sky130_fd_sc_hd__clkinv_2 _4385_ (.A(_0502_),
    .Y(_0897_));
 sky130_fd_sc_hd__nand2_1 _4386_ (.A(_0497_),
    .B(_0505_),
    .Y(_0898_));
 sky130_fd_sc_hd__o21ai_1 _4387_ (.A1(_0897_),
    .A2(_0495_),
    .B1(_0898_),
    .Y(_0899_));
 sky130_fd_sc_hd__a221oi_1 _4388_ (.A1(_0491_),
    .A2(_0487_),
    .B1(_0498_),
    .B2(_0490_),
    .C1(_0899_),
    .Y(_0900_));
 sky130_fd_sc_hd__inv_2 _4389_ (.A(_0511_),
    .Y(_0901_));
 sky130_fd_sc_hd__nand2_1 _4390_ (.A(_0504_),
    .B(_0515_),
    .Y(_0902_));
 sky130_fd_sc_hd__o21ai_1 _4391_ (.A1(_0510_),
    .A2(_0506_),
    .B1(_0902_),
    .Y(_0903_));
 sky130_fd_sc_hd__a221oi_1 _4392_ (.A1(_0519_),
    .A2(_0514_),
    .B1(_0527_),
    .B2(_0901_),
    .C1(_0903_),
    .Y(_0904_));
 sky130_fd_sc_hd__o22a_1 _4393_ (.A1(_0524_),
    .A2(_0530_),
    .B1(_0532_),
    .B2(_0523_),
    .X(_0905_));
 sky130_fd_sc_hd__o221a_1 _4394_ (.A1(_0699_),
    .A2(_0534_),
    .B1(_0543_),
    .B2(_0526_),
    .C1(_0905_),
    .X(_0906_));
 sky130_fd_sc_hd__inv_2 _4395_ (.A(_0540_),
    .Y(_0907_));
 sky130_fd_sc_hd__nand2_1 _4396_ (.A(_0548_),
    .B(_0537_),
    .Y(_0908_));
 sky130_fd_sc_hd__o21ai_1 _4397_ (.A1(_0907_),
    .A2(_0546_),
    .B1(_0908_),
    .Y(_0909_));
 sky130_fd_sc_hd__a221oi_1 _4398_ (.A1(\egd_top.BitStream_buffer.BS_buffer[32] ),
    .A2(_0539_),
    .B1(_0365_),
    .B2(_0542_),
    .C1(_0909_),
    .Y(_0910_));
 sky130_fd_sc_hd__and4_1 _4399_ (.A(_0900_),
    .B(_0904_),
    .C(_0906_),
    .D(_0910_),
    .X(_0911_));
 sky130_fd_sc_hd__nand2_1 _4400_ (.A(_0565_),
    .B(_0562_),
    .Y(_0912_));
 sky130_fd_sc_hd__nand2_1 _4401_ (.A(_0561_),
    .B(_0579_),
    .Y(_0913_));
 sky130_fd_sc_hd__or2_1 _4402_ (.A(_0554_),
    .B(_0571_),
    .X(_0914_));
 sky130_fd_sc_hd__o2111a_1 _4403_ (.A1(_0586_),
    .A2(_0558_),
    .B1(_0912_),
    .C1(_0913_),
    .D1(_0914_),
    .X(_0915_));
 sky130_fd_sc_hd__nand2_1 _4404_ (.A(_0578_),
    .B(_0583_),
    .Y(_0916_));
 sky130_fd_sc_hd__nand2_1 _4405_ (.A(_0582_),
    .B(\egd_top.BitStream_buffer.BS_buffer[12] ),
    .Y(_0917_));
 sky130_fd_sc_hd__or2_1 _4406_ (.A(_0574_),
    .B(_0588_),
    .X(_0918_));
 sky130_fd_sc_hd__o2111a_1 _4407_ (.A1(_0611_),
    .A2(_0576_),
    .B1(_0916_),
    .C1(_0917_),
    .D1(_0918_),
    .X(_0919_));
 sky130_fd_sc_hd__or2_1 _4408_ (.A(_0597_),
    .B(_0595_),
    .X(_0920_));
 sky130_fd_sc_hd__o221a_1 _4409_ (.A1(_0682_),
    .A2(_0593_),
    .B1(_0569_),
    .B2(_0599_),
    .C1(_0920_),
    .X(_0921_));
 sky130_fd_sc_hd__clkinv_2 _4410_ (.A(\egd_top.BitStream_buffer.BS_buffer[17] ),
    .Y(_0922_));
 sky130_fd_sc_hd__nand2_1 _4411_ (.A(_0606_),
    .B(\egd_top.BitStream_buffer.BS_buffer[14] ),
    .Y(_0923_));
 sky130_fd_sc_hd__nand2_1 _4412_ (.A(_0609_),
    .B(\egd_top.BitStream_buffer.BS_buffer[16] ),
    .Y(_0924_));
 sky130_fd_sc_hd__or2_1 _4413_ (.A(_0602_),
    .B(_0613_),
    .X(_0925_));
 sky130_fd_sc_hd__o2111a_1 _4414_ (.A1(_0922_),
    .A2(_0604_),
    .B1(_0923_),
    .C1(_0924_),
    .D1(_0925_),
    .X(_0926_));
 sky130_fd_sc_hd__and4_1 _4415_ (.A(_0915_),
    .B(_0919_),
    .C(_0921_),
    .D(_0926_),
    .X(_0927_));
 sky130_fd_sc_hd__nand2_1 _4416_ (.A(_0911_),
    .B(_0927_),
    .Y(_0928_));
 sky130_fd_sc_hd__nor2_1 _4417_ (.A(_0896_),
    .B(_0928_),
    .Y(_0929_));
 sky130_fd_sc_hd__clkbuf_4 _4418_ (.A(\egd_top.BitStream_buffer.BS_buffer[2] ),
    .X(_0930_));
 sky130_fd_sc_hd__nand2_1 _4419_ (.A(_0622_),
    .B(_0930_),
    .Y(_0931_));
 sky130_fd_sc_hd__nand3_1 _4420_ (.A(_0860_),
    .B(_0929_),
    .C(_0931_),
    .Y(_0932_));
 sky130_fd_sc_hd__inv_2 _4421_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[13] ),
    .Y(_0933_));
 sky130_fd_sc_hd__a21oi_1 _4422_ (.A1(_0933_),
    .A2(_3027_),
    .B1(_2905_),
    .Y(_0934_));
 sky130_fd_sc_hd__o21a_1 _4423_ (.A1(_3027_),
    .A2(_0932_),
    .B1(_0934_),
    .X(_0295_));
 sky130_fd_sc_hd__o21ai_1 _4424_ (.A1(\egd_top.BitStream_buffer.BitStream_buffer_output[12] ),
    .A2(_2965_),
    .B1(_0627_),
    .Y(_0935_));
 sky130_fd_sc_hd__inv_2 _4425_ (.A(\egd_top.BitStream_buffer.BS_buffer[42] ),
    .Y(_0936_));
 sky130_fd_sc_hd__nand2_1 _4426_ (.A(_0353_),
    .B(_0379_),
    .Y(_0937_));
 sky130_fd_sc_hd__o21ai_1 _4427_ (.A1(_0936_),
    .A2(_0350_),
    .B1(_0937_),
    .Y(_0938_));
 sky130_fd_sc_hd__a221oi_1 _4428_ (.A1(_0347_),
    .A2(_0342_),
    .B1(_0345_),
    .B2(_0375_),
    .C1(_0938_),
    .Y(_0939_));
 sky130_fd_sc_hd__clkinv_2 _4429_ (.A(_0337_),
    .Y(_0940_));
 sky130_fd_sc_hd__nand2_1 _4430_ (.A(_0370_),
    .B(_0364_),
    .Y(_0941_));
 sky130_fd_sc_hd__o21ai_1 _4431_ (.A1(_0940_),
    .A2(_0367_),
    .B1(_0941_),
    .Y(_0942_));
 sky130_fd_sc_hd__a221oi_1 _4432_ (.A1(_0346_),
    .A2(_0359_),
    .B1(_0362_),
    .B2(_0354_),
    .C1(_0942_),
    .Y(_0943_));
 sky130_fd_sc_hd__inv_2 _4433_ (.A(_0385_),
    .Y(_0944_));
 sky130_fd_sc_hd__nand2_1 _4434_ (.A(_0377_),
    .B(_0869_),
    .Y(_0945_));
 sky130_fd_sc_hd__o21ai_1 _4435_ (.A1(_0637_),
    .A2(_0380_),
    .B1(_0945_),
    .Y(_0946_));
 sky130_fd_sc_hd__a221oi_1 _4436_ (.A1(_0400_),
    .A2(_0388_),
    .B1(_0407_),
    .B2(_0944_),
    .C1(_0946_),
    .Y(_0947_));
 sky130_fd_sc_hd__buf_2 _4437_ (.A(\egd_top.BitStream_buffer.BS_buffer[49] ),
    .X(_0948_));
 sky130_fd_sc_hd__nand2_1 _4438_ (.A(_0406_),
    .B(_0948_),
    .Y(_0949_));
 sky130_fd_sc_hd__o21ai_1 _4439_ (.A1(_0659_),
    .A2(_0403_),
    .B1(_0949_),
    .Y(_0950_));
 sky130_fd_sc_hd__a221oi_1 _4440_ (.A1(_0642_),
    .A2(_0396_),
    .B1(_0399_),
    .B2(_0874_),
    .C1(_0950_),
    .Y(_0951_));
 sky130_fd_sc_hd__and4_1 _4441_ (.A(_0939_),
    .B(_0943_),
    .C(_0947_),
    .D(_0951_),
    .X(_0952_));
 sky130_fd_sc_hd__a22o_1 _4442_ (.A1(_0751_),
    .A2(_0476_),
    .B1(_2936_),
    .B2(_3230_),
    .X(_0953_));
 sky130_fd_sc_hd__a221oi_1 _4443_ (.A1(_0664_),
    .A2(_0470_),
    .B1(_3244_),
    .B2(_0473_),
    .C1(_0953_),
    .Y(_0954_));
 sky130_fd_sc_hd__inv_2 _4444_ (.A(\egd_top.BitStream_buffer.BS_buffer[62] ),
    .Y(_0955_));
 sky130_fd_sc_hd__nand2_1 _4445_ (.A(_0452_),
    .B(_0447_),
    .Y(_0956_));
 sky130_fd_sc_hd__nand2_1 _4446_ (.A(_0458_),
    .B(_0471_),
    .Y(_0957_));
 sky130_fd_sc_hd__or2_1 _4447_ (.A(_0647_),
    .B(_0463_),
    .X(_0958_));
 sky130_fd_sc_hd__o2111a_1 _4448_ (.A1(_0955_),
    .A2(_0450_),
    .B1(_0956_),
    .C1(_0957_),
    .D1(_0958_),
    .X(_0959_));
 sky130_fd_sc_hd__clkinv_2 _4449_ (.A(_0443_),
    .Y(_0960_));
 sky130_fd_sc_hd__or2_1 _4450_ (.A(_0879_),
    .B(_0424_),
    .X(_0961_));
 sky130_fd_sc_hd__nand2_1 _4451_ (.A(_0414_),
    .B(_0655_),
    .Y(_0962_));
 sky130_fd_sc_hd__nand2_1 _4452_ (.A(_0418_),
    .B(_0429_),
    .Y(_0963_));
 sky130_fd_sc_hd__o2111a_1 _4453_ (.A1(_0960_),
    .A2(_0421_),
    .B1(_0961_),
    .C1(_0962_),
    .D1(_0963_),
    .X(_0964_));
 sky130_fd_sc_hd__clkinv_2 _4454_ (.A(\egd_top.BitStream_buffer.BS_buffer[56] ),
    .Y(_0965_));
 sky130_fd_sc_hd__nand2_1 _4455_ (.A(_0431_),
    .B(_0461_),
    .Y(_0966_));
 sky130_fd_sc_hd__nand2_1 _4456_ (.A(_0441_),
    .B(_0436_),
    .Y(_0967_));
 sky130_fd_sc_hd__nand2_1 _4457_ (.A(_0434_),
    .B(_0459_),
    .Y(_0968_));
 sky130_fd_sc_hd__o2111a_1 _4458_ (.A1(_0965_),
    .A2(_0438_),
    .B1(_0966_),
    .C1(_0967_),
    .D1(_0968_),
    .X(_0969_));
 sky130_fd_sc_hd__and4_1 _4459_ (.A(_0954_),
    .B(_0959_),
    .C(_0964_),
    .D(_0969_),
    .X(_0970_));
 sky130_fd_sc_hd__nand2_1 _4460_ (.A(_0564_),
    .B(_0553_),
    .Y(_0971_));
 sky130_fd_sc_hd__nand2_1 _4461_ (.A(_0560_),
    .B(_0585_),
    .Y(_0972_));
 sky130_fd_sc_hd__or2_1 _4462_ (.A(_0670_),
    .B(_0570_),
    .X(_0973_));
 sky130_fd_sc_hd__o2111a_1 _4463_ (.A1(_0679_),
    .A2(_0557_),
    .B1(_0971_),
    .C1(_0972_),
    .D1(_0973_),
    .X(_0974_));
 sky130_fd_sc_hd__nand2_1 _4464_ (.A(_0577_),
    .B(\egd_top.BitStream_buffer.BS_buffer[11] ),
    .Y(_0975_));
 sky130_fd_sc_hd__nand2_1 _4465_ (.A(_0581_),
    .B(\egd_top.BitStream_buffer.BS_buffer[13] ),
    .Y(_0976_));
 sky130_fd_sc_hd__or2_1 _4466_ (.A(_0676_),
    .B(_0587_),
    .X(_0977_));
 sky130_fd_sc_hd__o2111a_1 _4467_ (.A1(_0688_),
    .A2(_0575_),
    .B1(_0975_),
    .C1(_0976_),
    .D1(_0977_),
    .X(_0978_));
 sky130_fd_sc_hd__or2_1 _4468_ (.A(_0673_),
    .B(_0598_),
    .X(_0979_));
 sky130_fd_sc_hd__o221a_1 _4469_ (.A1(_0569_),
    .A2(_0592_),
    .B1(_0682_),
    .B2(_0596_),
    .C1(_0979_),
    .X(_0980_));
 sky130_fd_sc_hd__nand2_1 _4470_ (.A(_0608_),
    .B(\egd_top.BitStream_buffer.BS_buffer[17] ),
    .Y(_0981_));
 sky130_fd_sc_hd__nand2_1 _4471_ (.A(_0605_),
    .B(\egd_top.BitStream_buffer.BS_buffer[15] ),
    .Y(_0982_));
 sky130_fd_sc_hd__or2_1 _4472_ (.A(_0685_),
    .B(_0612_),
    .X(_0983_));
 sky130_fd_sc_hd__o2111a_1 _4473_ (.A1(_0492_),
    .A2(_0603_),
    .B1(_0981_),
    .C1(_0982_),
    .D1(_0983_),
    .X(_0984_));
 sky130_fd_sc_hd__and4_1 _4474_ (.A(_0974_),
    .B(_0978_),
    .C(_0980_),
    .D(_0984_),
    .X(_0985_));
 sky130_fd_sc_hd__clkinv_2 _4475_ (.A(_0505_),
    .Y(_0986_));
 sky130_fd_sc_hd__nand2_1 _4476_ (.A(_0486_),
    .B(_0498_),
    .Y(_0987_));
 sky130_fd_sc_hd__nand2_1 _4477_ (.A(_0496_),
    .B(_0515_),
    .Y(_0988_));
 sky130_fd_sc_hd__nand2_1 _4478_ (.A(_0489_),
    .B(_0502_),
    .Y(_0989_));
 sky130_fd_sc_hd__o2111a_1 _4479_ (.A1(_0986_),
    .A2(_0494_),
    .B1(_0987_),
    .C1(_0988_),
    .D1(_0989_),
    .X(_0990_));
 sky130_fd_sc_hd__nand2_1 _4480_ (.A(_0513_),
    .B(_0527_),
    .Y(_0991_));
 sky130_fd_sc_hd__nand2_1 _4481_ (.A(_0503_),
    .B(_0509_),
    .Y(_0992_));
 sky130_fd_sc_hd__nand2_1 _4482_ (.A(_0507_),
    .B(_0519_),
    .Y(_0993_));
 sky130_fd_sc_hd__o2111a_1 _4483_ (.A1(_0532_),
    .A2(_0512_),
    .B1(_0991_),
    .C1(_0992_),
    .D1(_0993_),
    .X(_0994_));
 sky130_fd_sc_hd__clkinv_2 _4484_ (.A(\egd_top.BitStream_buffer.BS_buffer[32] ),
    .Y(_0995_));
 sky130_fd_sc_hd__nand2_1 _4485_ (.A(_0547_),
    .B(_0540_),
    .Y(_0996_));
 sky130_fd_sc_hd__o21ai_1 _4486_ (.A1(_0995_),
    .A2(_0545_),
    .B1(_0996_),
    .Y(_0997_));
 sky130_fd_sc_hd__a221oi_1 _4487_ (.A1(_0365_),
    .A2(_0538_),
    .B1(\egd_top.BitStream_buffer.BS_buffer[34] ),
    .B2(_0541_),
    .C1(_0997_),
    .Y(_0998_));
 sky130_fd_sc_hd__o22a_1 _4488_ (.A1(_0699_),
    .A2(_0529_),
    .B1(_0543_),
    .B2(_0533_),
    .X(_0999_));
 sky130_fd_sc_hd__o221a_1 _4489_ (.A1(_0524_),
    .A2(_0522_),
    .B1(_0702_),
    .B2(_0525_),
    .C1(_0999_),
    .X(_1000_));
 sky130_fd_sc_hd__and4_1 _4490_ (.A(_0990_),
    .B(_0994_),
    .C(_0998_),
    .D(_1000_),
    .X(_1001_));
 sky130_fd_sc_hd__and4_1 _4491_ (.A(_0952_),
    .B(_0970_),
    .C(_0985_),
    .D(_1001_),
    .X(_1002_));
 sky130_fd_sc_hd__clkinv_2 _4492_ (.A(\egd_top.BitStream_buffer.BS_buffer[92] ),
    .Y(_1003_));
 sky130_fd_sc_hd__nand2_1 _4493_ (.A(_3332_),
    .B(_3327_),
    .Y(_1004_));
 sky130_fd_sc_hd__o21ai_1 _4494_ (.A1(_1003_),
    .A2(_3329_),
    .B1(_1004_),
    .Y(_1005_));
 sky130_fd_sc_hd__a221oi_1 _4495_ (.A1(_0785_),
    .A2(_3324_),
    .B1(_3326_),
    .B2(_3338_),
    .C1(_1005_),
    .Y(_1006_));
 sky130_fd_sc_hd__inv_2 _4496_ (.A(\egd_top.BitStream_buffer.BS_buffer[83] ),
    .Y(_1007_));
 sky130_fd_sc_hd__nand2_1 _4497_ (.A(_3291_),
    .B(_0774_),
    .Y(_1008_));
 sky130_fd_sc_hd__nand2_1 _4498_ (.A(_3294_),
    .B(_3311_),
    .Y(_1009_));
 sky130_fd_sc_hd__nand2_1 _4499_ (.A(_3300_),
    .B(_3315_),
    .Y(_1010_));
 sky130_fd_sc_hd__o2111a_1 _4500_ (.A1(_1007_),
    .A2(_3298_),
    .B1(_1008_),
    .C1(_1009_),
    .D1(_1010_),
    .X(_1011_));
 sky130_fd_sc_hd__nand2_1 _4501_ (.A(_3313_),
    .B(\egd_top.BitStream_buffer.BS_buffer[87] ),
    .Y(_1012_));
 sky130_fd_sc_hd__nand2_1 _4502_ (.A(_3309_),
    .B(_0780_),
    .Y(_1013_));
 sky130_fd_sc_hd__or2_1 _4503_ (.A(_0776_),
    .B(_3318_),
    .X(_1014_));
 sky130_fd_sc_hd__o2111a_1 _4504_ (.A1(_0779_),
    .A2(_3307_),
    .B1(_1012_),
    .C1(_1013_),
    .D1(_1014_),
    .X(_1015_));
 sky130_fd_sc_hd__inv_2 _4505_ (.A(\egd_top.BitStream_buffer.BS_buffer[96] ),
    .Y(_1016_));
 sky130_fd_sc_hd__nand2_1 _4506_ (.A(_0328_),
    .B(_3341_),
    .Y(_1017_));
 sky130_fd_sc_hd__o21ai_1 _4507_ (.A1(_1016_),
    .A2(_0326_),
    .B1(_1017_),
    .Y(_1018_));
 sky130_fd_sc_hd__a221oi_1 _4508_ (.A1(_3040_),
    .A2(_3339_),
    .B1(_0708_),
    .B2(_0322_),
    .C1(_1018_),
    .Y(_1019_));
 sky130_fd_sc_hd__and4_1 _4509_ (.A(_1006_),
    .B(_1011_),
    .C(_1015_),
    .D(_1019_),
    .X(_1020_));
 sky130_fd_sc_hd__nand2_1 _4510_ (.A(_3098_),
    .B(_0722_),
    .Y(_1021_));
 sky130_fd_sc_hd__nand2_1 _4511_ (.A(_3093_),
    .B(_0714_),
    .Y(_1022_));
 sky130_fd_sc_hd__or2_1 _4512_ (.A(_0721_),
    .B(_3088_),
    .X(_1023_));
 sky130_fd_sc_hd__o2111a_1 _4513_ (.A1(_0718_),
    .A2(_3106_),
    .B1(_1021_),
    .C1(_1022_),
    .D1(_1023_),
    .X(_1024_));
 sky130_fd_sc_hd__inv_2 _4514_ (.A(\egd_top.BitStream_buffer.BS_buffer[108] ),
    .Y(_1025_));
 sky130_fd_sc_hd__nand2_1 _4515_ (.A(_3126_),
    .B(_3118_),
    .Y(_1026_));
 sky130_fd_sc_hd__nand2_1 _4516_ (.A(_3112_),
    .B(_3070_),
    .Y(_1027_));
 sky130_fd_sc_hd__nand2_1 _4517_ (.A(_3116_),
    .B(_3075_),
    .Y(_1028_));
 sky130_fd_sc_hd__o2111a_1 _4518_ (.A1(_1025_),
    .A2(_3122_),
    .B1(_1026_),
    .C1(_1027_),
    .D1(_1028_),
    .X(_1029_));
 sky130_fd_sc_hd__nand2_1 _4519_ (.A(_3060_),
    .B(\egd_top.BitStream_buffer.BS_buffer[102] ),
    .Y(_1030_));
 sky130_fd_sc_hd__nand2_1 _4520_ (.A(_3047_),
    .B(\egd_top.BitStream_buffer.BS_buffer[100] ),
    .Y(_1031_));
 sky130_fd_sc_hd__nand2_1 _4521_ (.A(_3054_),
    .B(\egd_top.BitStream_buffer.BS_buffer[101] ),
    .Y(_1032_));
 sky130_fd_sc_hd__nand2_1 _4522_ (.A(_3038_),
    .B(_3062_),
    .Y(_1033_));
 sky130_fd_sc_hd__and4_1 _4523_ (.A(_1030_),
    .B(_1031_),
    .C(_1032_),
    .D(_1033_),
    .X(_1034_));
 sky130_fd_sc_hd__clkinv_2 _4524_ (.A(\egd_top.BitStream_buffer.BS_buffer[111] ),
    .Y(_1035_));
 sky130_fd_sc_hd__nand2_1 _4525_ (.A(_3073_),
    .B(_3169_),
    .Y(_1036_));
 sky130_fd_sc_hd__o21ai_1 _4526_ (.A1(_1035_),
    .A2(_0728_),
    .B1(_1036_),
    .Y(_1037_));
 sky130_fd_sc_hd__a221oi_1 _4527_ (.A1(_3164_),
    .A2(_3078_),
    .B1(_3153_),
    .B2(_3080_),
    .C1(_1037_),
    .Y(_1038_));
 sky130_fd_sc_hd__and4_1 _4528_ (.A(_1024_),
    .B(_1029_),
    .C(_1034_),
    .D(_1038_),
    .X(_1039_));
 sky130_fd_sc_hd__nand2_1 _4529_ (.A(_3215_),
    .B(_3227_),
    .Y(_1040_));
 sky130_fd_sc_hd__o21ai_1 _4530_ (.A1(_3257_),
    .A2(_3218_),
    .B1(_1040_),
    .Y(_1041_));
 sky130_fd_sc_hd__a221oi_2 _4531_ (.A1(_3264_),
    .A2(_3224_),
    .B1(_3248_),
    .B2(_3226_),
    .C1(_1041_),
    .Y(_1042_));
 sky130_fd_sc_hd__inv_2 _4532_ (.A(\egd_top.BitStream_buffer.BS_buffer[68] ),
    .Y(_1043_));
 sky130_fd_sc_hd__nand2_1 _4533_ (.A(_3232_),
    .B(\egd_top.BitStream_buffer.BS_buffer[69] ),
    .Y(_1044_));
 sky130_fd_sc_hd__nand2_1 _4534_ (.A(_3242_),
    .B(_3237_),
    .Y(_1045_));
 sky130_fd_sc_hd__nand2_1 _4535_ (.A(_3235_),
    .B(_3221_),
    .Y(_1046_));
 sky130_fd_sc_hd__o2111a_1 _4536_ (.A1(_1043_),
    .A2(_3239_),
    .B1(_1044_),
    .C1(_1045_),
    .D1(_1046_),
    .X(_1047_));
 sky130_fd_sc_hd__nand2_1 _4537_ (.A(_3262_),
    .B(\egd_top.BitStream_buffer.BS_buffer[76] ),
    .Y(_1048_));
 sky130_fd_sc_hd__nand2_1 _4538_ (.A(_3254_),
    .B(\egd_top.BitStream_buffer.BS_buffer[78] ),
    .Y(_1049_));
 sky130_fd_sc_hd__nand2_1 _4539_ (.A(_3250_),
    .B(\egd_top.BitStream_buffer.BS_buffer[77] ),
    .Y(_1050_));
 sky130_fd_sc_hd__nand2_1 _4540_ (.A(_3259_),
    .B(\egd_top.BitStream_buffer.BS_buffer[75] ),
    .Y(_1051_));
 sky130_fd_sc_hd__and4_1 _4541_ (.A(_1048_),
    .B(_1049_),
    .C(_1050_),
    .D(_1051_),
    .X(_1052_));
 sky130_fd_sc_hd__nand2_1 _4542_ (.A(_3281_),
    .B(_3302_),
    .Y(_1053_));
 sky130_fd_sc_hd__o21ai_1 _4543_ (.A1(_0842_),
    .A2(_3279_),
    .B1(_1053_),
    .Y(_1054_));
 sky130_fd_sc_hd__a221oi_1 _4544_ (.A1(_3276_),
    .A2(_3270_),
    .B1(_0837_),
    .B2(_3274_),
    .C1(_1054_),
    .Y(_1055_));
 sky130_fd_sc_hd__and4_1 _4545_ (.A(_1042_),
    .B(_1047_),
    .C(_1052_),
    .D(_1055_),
    .X(_1056_));
 sky130_fd_sc_hd__nand2_1 _4546_ (.A(_3202_),
    .B(_3198_),
    .Y(_1057_));
 sky130_fd_sc_hd__nand2_1 _4547_ (.A(_3193_),
    .B(\egd_top.BitStream_buffer.BS_buffer[121] ),
    .Y(_1058_));
 sky130_fd_sc_hd__nand2_1 _4548_ (.A(_3196_),
    .B(\egd_top.BitStream_buffer.BS_buffer[122] ),
    .Y(_1059_));
 sky130_fd_sc_hd__o2111a_1 _4549_ (.A1(_3003_),
    .A2(_3199_),
    .B1(_1057_),
    .C1(_1058_),
    .D1(_1059_),
    .X(_1060_));
 sky130_fd_sc_hd__nand2_1 _4550_ (.A(_3162_),
    .B(\egd_top.BitStream_buffer.BS_buffer[116] ),
    .Y(_1061_));
 sky130_fd_sc_hd__nand2_1 _4551_ (.A(_3159_),
    .B(\egd_top.BitStream_buffer.BS_buffer[118] ),
    .Y(_1062_));
 sky130_fd_sc_hd__nand2_1 _4552_ (.A(_3167_),
    .B(\egd_top.BitStream_buffer.BS_buffer[115] ),
    .Y(_1063_));
 sky130_fd_sc_hd__nand2_1 _4553_ (.A(_3155_),
    .B(\egd_top.BitStream_buffer.BS_buffer[117] ),
    .Y(_1064_));
 sky130_fd_sc_hd__and4_1 _4554_ (.A(_1061_),
    .B(_1062_),
    .C(_1063_),
    .D(_1064_),
    .X(_1065_));
 sky130_fd_sc_hd__nand2_1 _4555_ (.A(_3140_),
    .B(_0741_),
    .Y(_1066_));
 sky130_fd_sc_hd__nand2_1 _4556_ (.A(_3147_),
    .B(\egd_top.BitStream_buffer.BS_buffer[124] ),
    .Y(_1067_));
 sky130_fd_sc_hd__nand2_1 _4557_ (.A(_3144_),
    .B(\egd_top.BitStream_buffer.BS_buffer[123] ),
    .Y(_1068_));
 sky130_fd_sc_hd__nand2_1 _4558_ (.A(_3136_),
    .B(\egd_top.BitStream_buffer.BS_buffer[125] ),
    .Y(_1069_));
 sky130_fd_sc_hd__and4_1 _4559_ (.A(_1066_),
    .B(_1067_),
    .C(_1068_),
    .D(_1069_),
    .X(_1070_));
 sky130_fd_sc_hd__nand2_1 _4560_ (.A(_3185_),
    .B(_0930_),
    .Y(_1071_));
 sky130_fd_sc_hd__o21ai_1 _4561_ (.A1(_0594_),
    .A2(_3183_),
    .B1(_1071_),
    .Y(_1072_));
 sky130_fd_sc_hd__a221oi_1 _4562_ (.A1(_3187_),
    .A2(_3176_),
    .B1(_0623_),
    .B2(_3179_),
    .C1(_1072_),
    .Y(_1073_));
 sky130_fd_sc_hd__and4_1 _4563_ (.A(_1060_),
    .B(_1065_),
    .C(_1070_),
    .D(_1073_),
    .X(_1074_));
 sky130_fd_sc_hd__and4_1 _4564_ (.A(_1020_),
    .B(_1039_),
    .C(_1056_),
    .D(_1074_),
    .X(_1075_));
 sky130_fd_sc_hd__clkbuf_4 _4565_ (.A(\egd_top.BitStream_buffer.BS_buffer[3] ),
    .X(_1076_));
 sky130_fd_sc_hd__nand2_1 _4566_ (.A(_0622_),
    .B(_1076_),
    .Y(_1077_));
 sky130_fd_sc_hd__nand3_1 _4567_ (.A(_1002_),
    .B(_1075_),
    .C(_1077_),
    .Y(_1078_));
 sky130_fd_sc_hd__nor2_1 _4568_ (.A(_3026_),
    .B(_1078_),
    .Y(_1079_));
 sky130_fd_sc_hd__nor2_1 _4569_ (.A(_0935_),
    .B(_1079_),
    .Y(_0294_));
 sky130_fd_sc_hd__o21ai_1 _4570_ (.A1(\egd_top.BitStream_buffer.BitStream_buffer_output[11] ),
    .A2(_2965_),
    .B1(_0627_),
    .Y(_1080_));
 sky130_fd_sc_hd__nand2_1 _4571_ (.A(_0352_),
    .B(\egd_top.BitStream_buffer.BS_buffer[42] ),
    .Y(_1081_));
 sky130_fd_sc_hd__o21ai_1 _4572_ (.A1(_0383_),
    .A2(_0349_),
    .B1(_1081_),
    .Y(_1082_));
 sky130_fd_sc_hd__a221oi_1 _4573_ (.A1(_0375_),
    .A2(_0341_),
    .B1(_0344_),
    .B2(_0379_),
    .C1(_1082_),
    .Y(_1083_));
 sky130_fd_sc_hd__clkinv_2 _4574_ (.A(_0346_),
    .Y(_1084_));
 sky130_fd_sc_hd__nand2_1 _4575_ (.A(_0370_),
    .B(_0337_),
    .Y(_1085_));
 sky130_fd_sc_hd__nand2_1 _4576_ (.A(_0359_),
    .B(_0354_),
    .Y(_1086_));
 sky130_fd_sc_hd__nand2_1 _4577_ (.A(_0362_),
    .B(_0347_),
    .Y(_1087_));
 sky130_fd_sc_hd__o2111a_1 _4578_ (.A1(_1084_),
    .A2(_0367_),
    .B1(_1085_),
    .C1(_1086_),
    .D1(_1087_),
    .X(_1088_));
 sky130_fd_sc_hd__nand2_1 _4579_ (.A(_0387_),
    .B(\egd_top.BitStream_buffer.BS_buffer[46] ),
    .Y(_1089_));
 sky130_fd_sc_hd__nand2_1 _4580_ (.A(_0377_),
    .B(\egd_top.BitStream_buffer.BS_buffer[44] ),
    .Y(_1090_));
 sky130_fd_sc_hd__nand2_1 _4581_ (.A(_0381_),
    .B(\egd_top.BitStream_buffer.BS_buffer[45] ),
    .Y(_1091_));
 sky130_fd_sc_hd__o2111a_1 _4582_ (.A1(_0401_),
    .A2(_0384_),
    .B1(_1089_),
    .C1(_1090_),
    .D1(_1091_),
    .X(_1092_));
 sky130_fd_sc_hd__nand2_1 _4583_ (.A(_0405_),
    .B(_0412_),
    .Y(_1093_));
 sky130_fd_sc_hd__o21ai_1 _4584_ (.A1(_0879_),
    .A2(_0402_),
    .B1(_1093_),
    .Y(_1094_));
 sky130_fd_sc_hd__a221oi_1 _4585_ (.A1(\egd_top.BitStream_buffer.BS_buffer[48] ),
    .A2(_0395_),
    .B1(_0398_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[49] ),
    .C1(_1094_),
    .Y(_1095_));
 sky130_fd_sc_hd__and4_1 _4586_ (.A(_1083_),
    .B(_1088_),
    .C(_1092_),
    .D(_1095_),
    .X(_1096_));
 sky130_fd_sc_hd__nand2_1 _4587_ (.A(_0457_),
    .B(_0478_),
    .Y(_1097_));
 sky130_fd_sc_hd__nand2_1 _4588_ (.A(_0452_),
    .B(_0467_),
    .Y(_1098_));
 sky130_fd_sc_hd__or2_1 _4589_ (.A(_0887_),
    .B(_0463_),
    .X(_1099_));
 sky130_fd_sc_hd__o2111a_1 _4590_ (.A1(_0474_),
    .A2(_0449_),
    .B1(_1097_),
    .C1(_1098_),
    .D1(_1099_),
    .X(_1100_));
 sky130_fd_sc_hd__nand2_1 _4591_ (.A(_0431_),
    .B(\egd_top.BitStream_buffer.BS_buffer[58] ),
    .Y(_1101_));
 sky130_fd_sc_hd__nand2_1 _4592_ (.A(_0441_),
    .B(_0454_),
    .Y(_1102_));
 sky130_fd_sc_hd__nand2_1 _4593_ (.A(_0434_),
    .B(_0447_),
    .Y(_1103_));
 sky130_fd_sc_hd__o2111a_1 _4594_ (.A1(_0462_),
    .A2(_0438_),
    .B1(_1101_),
    .C1(_1102_),
    .D1(_1103_),
    .X(_1104_));
 sky130_fd_sc_hd__o22ai_1 _4595_ (.A1(_0960_),
    .A2(_0424_),
    .B1(_0437_),
    .B2(_0421_),
    .Y(_1105_));
 sky130_fd_sc_hd__a22o_1 _4596_ (.A1(\egd_top.BitStream_buffer.BS_buffer[54] ),
    .A2(_0414_),
    .B1(_0418_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[55] ),
    .X(_1106_));
 sky130_fd_sc_hd__nor2_1 _4597_ (.A(_1105_),
    .B(_1106_),
    .Y(_1107_));
 sky130_fd_sc_hd__nand2_1 _4598_ (.A(_0476_),
    .B(\egd_top.BitStream_buffer.BS_buffer[66] ),
    .Y(_1108_));
 sky130_fd_sc_hd__o21ai_1 _4599_ (.A1(_0829_),
    .A2(_2935_),
    .B1(_1108_),
    .Y(_1109_));
 sky130_fd_sc_hd__a221oi_1 _4600_ (.A1(\egd_top.BitStream_buffer.BS_buffer[64] ),
    .A2(_0469_),
    .B1(_0751_),
    .B2(_0473_),
    .C1(_1109_),
    .Y(_1110_));
 sky130_fd_sc_hd__and4_1 _4601_ (.A(_1100_),
    .B(_1104_),
    .C(_1107_),
    .D(_1110_),
    .X(_1111_));
 sky130_fd_sc_hd__and2_1 _4602_ (.A(_1096_),
    .B(_1111_),
    .X(_1112_));
 sky130_fd_sc_hd__nand2_1 _4603_ (.A(_0564_),
    .B(_0579_),
    .Y(_1113_));
 sky130_fd_sc_hd__nand2_1 _4604_ (.A(_0560_),
    .B(_0583_),
    .Y(_1114_));
 sky130_fd_sc_hd__or2_1 _4605_ (.A(_0586_),
    .B(_0570_),
    .X(_1115_));
 sky130_fd_sc_hd__o2111a_1 _4606_ (.A1(_0574_),
    .A2(_0558_),
    .B1(_1113_),
    .C1(_1114_),
    .D1(_1115_),
    .X(_1116_));
 sky130_fd_sc_hd__nand2_1 _4607_ (.A(_0577_),
    .B(\egd_top.BitStream_buffer.BS_buffer[12] ),
    .Y(_1117_));
 sky130_fd_sc_hd__nand2_1 _4608_ (.A(_0581_),
    .B(\egd_top.BitStream_buffer.BS_buffer[14] ),
    .Y(_1118_));
 sky130_fd_sc_hd__or2_1 _4609_ (.A(_0611_),
    .B(_0587_),
    .X(_1119_));
 sky130_fd_sc_hd__o2111a_1 _4610_ (.A1(_0602_),
    .A2(_0576_),
    .B1(_1117_),
    .C1(_1118_),
    .D1(_1119_),
    .X(_1120_));
 sky130_fd_sc_hd__or2_1 _4611_ (.A(_0554_),
    .B(_0598_),
    .X(_1121_));
 sky130_fd_sc_hd__o221a_1 _4612_ (.A1(_0673_),
    .A2(_0592_),
    .B1(_0569_),
    .B2(_0596_),
    .C1(_1121_),
    .X(_1122_));
 sky130_fd_sc_hd__nand2_1 _4613_ (.A(_0608_),
    .B(_0491_),
    .Y(_1123_));
 sky130_fd_sc_hd__nand2_1 _4614_ (.A(_0605_),
    .B(\egd_top.BitStream_buffer.BS_buffer[16] ),
    .Y(_1124_));
 sky130_fd_sc_hd__or2_1 _4615_ (.A(_0922_),
    .B(_0612_),
    .X(_1125_));
 sky130_fd_sc_hd__o2111a_1 _4616_ (.A1(_0692_),
    .A2(_0604_),
    .B1(_1123_),
    .C1(_1124_),
    .D1(_1125_),
    .X(_1126_));
 sky130_fd_sc_hd__and4_1 _4617_ (.A(_1116_),
    .B(_1120_),
    .C(_1122_),
    .D(_1126_),
    .X(_1127_));
 sky130_fd_sc_hd__clkinv_2 _4618_ (.A(\egd_top.BitStream_buffer.BS_buffer[22] ),
    .Y(_1128_));
 sky130_fd_sc_hd__nand2_1 _4619_ (.A(_0496_),
    .B(_0509_),
    .Y(_1129_));
 sky130_fd_sc_hd__o21ai_1 _4620_ (.A1(_1128_),
    .A2(_0494_),
    .B1(_1129_),
    .Y(_1130_));
 sky130_fd_sc_hd__a221oi_1 _4621_ (.A1(_0502_),
    .A2(_0486_),
    .B1(_0505_),
    .B2(_0489_),
    .C1(_1130_),
    .Y(_1131_));
 sky130_fd_sc_hd__nand2_1 _4622_ (.A(_0513_),
    .B(_0531_),
    .Y(_1132_));
 sky130_fd_sc_hd__o21ai_1 _4623_ (.A1(_0524_),
    .A2(_0512_),
    .B1(_1132_),
    .Y(_1133_));
 sky130_fd_sc_hd__a221oi_1 _4624_ (.A1(_0519_),
    .A2(_0504_),
    .B1(_0527_),
    .B2(_0508_),
    .C1(_1133_),
    .Y(_1134_));
 sky130_fd_sc_hd__o22a_1 _4625_ (.A1(_0543_),
    .A2(_0529_),
    .B1(_0907_),
    .B2(_0525_),
    .X(_1135_));
 sky130_fd_sc_hd__o221a_1 _4626_ (.A1(_0699_),
    .A2(_0522_),
    .B1(_0702_),
    .B2(_0534_),
    .C1(_1135_),
    .X(_1136_));
 sky130_fd_sc_hd__nand2_1 _4627_ (.A(_0547_),
    .B(\egd_top.BitStream_buffer.BS_buffer[32] ),
    .Y(_1137_));
 sky130_fd_sc_hd__o21ai_1 _4628_ (.A1(_0366_),
    .A2(_0545_),
    .B1(_1137_),
    .Y(_1138_));
 sky130_fd_sc_hd__a221oi_1 _4629_ (.A1(\egd_top.BitStream_buffer.BS_buffer[34] ),
    .A2(_0538_),
    .B1(_0364_),
    .B2(_0541_),
    .C1(_1138_),
    .Y(_1139_));
 sky130_fd_sc_hd__and4_1 _4630_ (.A(_1131_),
    .B(_1134_),
    .C(_1136_),
    .D(_1139_),
    .X(_1140_));
 sky130_fd_sc_hd__and3_1 _4631_ (.A(_1112_),
    .B(_1127_),
    .C(_1140_),
    .X(_1141_));
 sky130_fd_sc_hd__a22o_1 _4632_ (.A1(_3210_),
    .A2(_3242_),
    .B1(_0752_),
    .B2(_3217_),
    .X(_1142_));
 sky130_fd_sc_hd__a221oi_1 _4633_ (.A1(_3221_),
    .A2(_3233_),
    .B1(_3227_),
    .B2(_3236_),
    .C1(_1142_),
    .Y(_1143_));
 sky130_fd_sc_hd__inv_2 _4634_ (.A(\egd_top.BitStream_buffer.BS_buffer[75] ),
    .Y(_1144_));
 sky130_fd_sc_hd__buf_2 _4635_ (.A(_3225_),
    .X(_1145_));
 sky130_fd_sc_hd__nand2_1 _4636_ (.A(_3224_),
    .B(\egd_top.BitStream_buffer.BS_buffer[74] ),
    .Y(_1146_));
 sky130_fd_sc_hd__o21ai_1 _4637_ (.A1(_1144_),
    .A2(_1145_),
    .B1(_1146_),
    .Y(_1147_));
 sky130_fd_sc_hd__a221oi_1 _4638_ (.A1(_3256_),
    .A2(_3216_),
    .B1(_3264_),
    .B2(_3220_),
    .C1(_1147_),
    .Y(_1148_));
 sky130_fd_sc_hd__inv_2 _4639_ (.A(\egd_top.BitStream_buffer.BS_buffer[76] ),
    .Y(_1149_));
 sky130_fd_sc_hd__nand2_1 _4640_ (.A(_3263_),
    .B(_3272_),
    .Y(_1150_));
 sky130_fd_sc_hd__o21ai_1 _4641_ (.A1(_1149_),
    .A2(_3260_),
    .B1(_1150_),
    .Y(_1151_));
 sky130_fd_sc_hd__a221oi_1 _4642_ (.A1(_3283_),
    .A2(_3251_),
    .B1(_3276_),
    .B2(_3255_),
    .C1(_1151_),
    .Y(_1152_));
 sky130_fd_sc_hd__inv_2 _4643_ (.A(_3278_),
    .Y(_1153_));
 sky130_fd_sc_hd__nand2_1 _4644_ (.A(_3271_),
    .B(_0837_),
    .Y(_1154_));
 sky130_fd_sc_hd__o21ai_1 _4645_ (.A1(_0767_),
    .A2(_3273_),
    .B1(_1154_),
    .Y(_1155_));
 sky130_fd_sc_hd__a221oi_1 _4646_ (.A1(_3288_),
    .A2(_3282_),
    .B1(_3293_),
    .B2(_1153_),
    .C1(_1155_),
    .Y(_1156_));
 sky130_fd_sc_hd__and4_1 _4647_ (.A(_1143_),
    .B(_1148_),
    .C(_1152_),
    .D(_1156_),
    .X(_1157_));
 sky130_fd_sc_hd__inv_2 _4648_ (.A(\egd_top.BitStream_buffer.BS_buffer[84] ),
    .Y(_1158_));
 sky130_fd_sc_hd__nand2_1 _4649_ (.A(_3301_),
    .B(_0774_),
    .Y(_1159_));
 sky130_fd_sc_hd__o21ai_1 _4650_ (.A1(_1158_),
    .A2(_3299_),
    .B1(_1159_),
    .Y(_1160_));
 sky130_fd_sc_hd__a221oi_1 _4651_ (.A1(_3311_),
    .A2(_3292_),
    .B1(_0772_),
    .B2(_3295_),
    .C1(_1160_),
    .Y(_1161_));
 sky130_fd_sc_hd__nand2_1 _4652_ (.A(_3314_),
    .B(_3334_),
    .Y(_1162_));
 sky130_fd_sc_hd__nand2_1 _4653_ (.A(_3310_),
    .B(_3322_),
    .Y(_1163_));
 sky130_fd_sc_hd__or2_1 _4654_ (.A(_3328_),
    .B(_3318_),
    .X(_1164_));
 sky130_fd_sc_hd__o2111a_1 _4655_ (.A1(_0850_),
    .A2(_3308_),
    .B1(_1162_),
    .C1(_1163_),
    .D1(_1164_),
    .X(_1165_));
 sky130_fd_sc_hd__nand2_1 _4656_ (.A(_3332_),
    .B(_0330_),
    .Y(_1166_));
 sky130_fd_sc_hd__o21ai_1 _4657_ (.A1(_0324_),
    .A2(_3330_),
    .B1(_1166_),
    .Y(_1167_));
 sky130_fd_sc_hd__a221oi_1 _4658_ (.A1(_3338_),
    .A2(_3324_),
    .B1(_3326_),
    .B2(_3341_),
    .C1(_1167_),
    .Y(_1168_));
 sky130_fd_sc_hd__inv_2 _4659_ (.A(\egd_top.BitStream_buffer.BS_buffer[97] ),
    .Y(_1169_));
 sky130_fd_sc_hd__nand2_1 _4660_ (.A(_0329_),
    .B(\egd_top.BitStream_buffer.BS_buffer[96] ),
    .Y(_1170_));
 sky130_fd_sc_hd__o21ai_1 _4661_ (.A1(_1169_),
    .A2(_0327_),
    .B1(_1170_),
    .Y(_1171_));
 sky130_fd_sc_hd__a221oi_1 _4662_ (.A1(_0708_),
    .A2(_3340_),
    .B1(_3062_),
    .B2(_0323_),
    .C1(_1171_),
    .Y(_1172_));
 sky130_fd_sc_hd__and4_1 _4663_ (.A(_1161_),
    .B(_1165_),
    .C(_1168_),
    .D(_1172_),
    .X(_1173_));
 sky130_fd_sc_hd__nand2_1 _4664_ (.A(_1157_),
    .B(_1173_),
    .Y(_1174_));
 sky130_fd_sc_hd__a22o_1 _4665_ (.A1(_3100_),
    .A2(_3054_),
    .B1(_3061_),
    .B2(_0714_),
    .X(_1175_));
 sky130_fd_sc_hd__a221oi_1 _4666_ (.A1(_3094_),
    .A2(_3039_),
    .B1(_0716_),
    .B2(_3048_),
    .C1(_1175_),
    .Y(_1176_));
 sky130_fd_sc_hd__nand2_1 _4667_ (.A(_3093_),
    .B(_3128_),
    .Y(_1177_));
 sky130_fd_sc_hd__nand2_1 _4668_ (.A(_3099_),
    .B(_3109_),
    .Y(_1178_));
 sky130_fd_sc_hd__or2_1 _4669_ (.A(_3119_),
    .B(_3105_),
    .X(_1179_));
 sky130_fd_sc_hd__o2111a_1 _4670_ (.A1(_0804_),
    .A2(_3089_),
    .B1(_1177_),
    .C1(_1178_),
    .D1(_1179_),
    .X(_1180_));
 sky130_fd_sc_hd__nand2_1 _4671_ (.A(_3127_),
    .B(_3066_),
    .Y(_1181_));
 sky130_fd_sc_hd__o21ai_1 _4672_ (.A1(_0727_),
    .A2(_3123_),
    .B1(_1181_),
    .Y(_1182_));
 sky130_fd_sc_hd__a221oi_1 _4673_ (.A1(_3075_),
    .A2(_3113_),
    .B1(_3117_),
    .B2(_3082_),
    .C1(_1182_),
    .Y(_1183_));
 sky130_fd_sc_hd__nand2_1 _4674_ (.A(_3074_),
    .B(_3164_),
    .Y(_1184_));
 sky130_fd_sc_hd__o21ai_1 _4675_ (.A1(_2977_),
    .A2(_0729_),
    .B1(_1184_),
    .Y(_1185_));
 sky130_fd_sc_hd__a221oi_1 _4676_ (.A1(_3153_),
    .A2(_0726_),
    .B1(_3157_),
    .B2(_3081_),
    .C1(_1185_),
    .Y(_1186_));
 sky130_fd_sc_hd__and4_1 _4677_ (.A(_1176_),
    .B(_1180_),
    .C(_1183_),
    .D(_1186_),
    .X(_1187_));
 sky130_fd_sc_hd__nand2_1 _4678_ (.A(_3148_),
    .B(_3177_),
    .Y(_1188_));
 sky130_fd_sc_hd__o21ai_1 _4679_ (.A1(_3015_),
    .A2(_3145_),
    .B1(_1188_),
    .Y(_1189_));
 sky130_fd_sc_hd__a221oi_1 _4680_ (.A1(_0741_),
    .A2(_3137_),
    .B1(_3187_),
    .B2(_3141_),
    .C1(_1189_),
    .Y(_1190_));
 sky130_fd_sc_hd__nand2_1 _4681_ (.A(_3163_),
    .B(_0746_),
    .Y(_1191_));
 sky130_fd_sc_hd__nand2_1 _4682_ (.A(_3168_),
    .B(_3204_),
    .Y(_1192_));
 sky130_fd_sc_hd__nand2_1 _4683_ (.A(_1191_),
    .B(_1192_),
    .Y(_1193_));
 sky130_fd_sc_hd__a221oi_1 _4684_ (.A1(_3191_),
    .A2(_3156_),
    .B1(_3198_),
    .B2(_3160_),
    .C1(_1193_),
    .Y(_1194_));
 sky130_fd_sc_hd__nand2_1 _4685_ (.A(_3203_),
    .B(_0744_),
    .Y(_1195_));
 sky130_fd_sc_hd__o21ai_1 _4686_ (.A1(_3006_),
    .A2(_3200_),
    .B1(_1195_),
    .Y(_1196_));
 sky130_fd_sc_hd__a221oi_1 _4687_ (.A1(_3133_),
    .A2(_3194_),
    .B1(_3197_),
    .B2(_3138_),
    .C1(_1196_),
    .Y(_1197_));
 sky130_fd_sc_hd__nand2_1 _4688_ (.A(_3186_),
    .B(_1076_),
    .Y(_1198_));
 sky130_fd_sc_hd__o21ai_1 _4689_ (.A1(_0591_),
    .A2(_3183_),
    .B1(_1198_),
    .Y(_1199_));
 sky130_fd_sc_hd__a221oi_1 _4690_ (.A1(_0623_),
    .A2(_3176_),
    .B1(_0792_),
    .B2(_3180_),
    .C1(_1199_),
    .Y(_1200_));
 sky130_fd_sc_hd__and4_1 _4691_ (.A(_1190_),
    .B(_1194_),
    .C(_1197_),
    .D(_1200_),
    .X(_1201_));
 sky130_fd_sc_hd__nand2_1 _4692_ (.A(_1187_),
    .B(_1201_),
    .Y(_1202_));
 sky130_fd_sc_hd__nor2_1 _4693_ (.A(_1174_),
    .B(_1202_),
    .Y(_1203_));
 sky130_fd_sc_hd__nand2_1 _4694_ (.A(_0622_),
    .B(_0566_),
    .Y(_1204_));
 sky130_fd_sc_hd__nand3_1 _4695_ (.A(_1141_),
    .B(_1203_),
    .C(_1204_),
    .Y(_1205_));
 sky130_fd_sc_hd__nor2_1 _4696_ (.A(_3026_),
    .B(_1205_),
    .Y(_1206_));
 sky130_fd_sc_hd__nor2_1 _4697_ (.A(_1080_),
    .B(_1206_),
    .Y(_0293_));
 sky130_fd_sc_hd__o21ai_1 _4698_ (.A1(\egd_top.BitStream_buffer.BitStream_buffer_output[10] ),
    .A2(_2965_),
    .B1(_0627_),
    .Y(_1207_));
 sky130_fd_sc_hd__nand2_1 _4699_ (.A(_3333_),
    .B(_0785_),
    .Y(_1208_));
 sky130_fd_sc_hd__o21ai_1 _4700_ (.A1(_0784_),
    .A2(_3330_),
    .B1(_1208_),
    .Y(_1209_));
 sky130_fd_sc_hd__a221oi_1 _4701_ (.A1(_3341_),
    .A2(_3324_),
    .B1(_3326_),
    .B2(_3028_),
    .C1(_1209_),
    .Y(_1210_));
 sky130_fd_sc_hd__nand2_1 _4702_ (.A(_3292_),
    .B(_0772_),
    .Y(_1211_));
 sky130_fd_sc_hd__nand2_1 _4703_ (.A(_3294_),
    .B(_3334_),
    .Y(_1212_));
 sky130_fd_sc_hd__nand2_1 _4704_ (.A(_3301_),
    .B(_3311_),
    .Y(_1213_));
 sky130_fd_sc_hd__o2111a_1 _4705_ (.A1(_3317_),
    .A2(_3299_),
    .B1(_1211_),
    .C1(_1212_),
    .D1(_1213_),
    .X(_1214_));
 sky130_fd_sc_hd__nand2_1 _4706_ (.A(_3314_),
    .B(_0780_),
    .Y(_1215_));
 sky130_fd_sc_hd__nand2_1 _4707_ (.A(_3310_),
    .B(_3327_),
    .Y(_1216_));
 sky130_fd_sc_hd__or2_1 _4708_ (.A(_0779_),
    .B(_3318_),
    .X(_1217_));
 sky130_fd_sc_hd__o2111a_1 _4709_ (.A1(_1003_),
    .A2(_3308_),
    .B1(_1215_),
    .C1(_1216_),
    .D1(_1217_),
    .X(_1218_));
 sky130_fd_sc_hd__nand2_1 _4710_ (.A(_0329_),
    .B(_3040_),
    .Y(_1219_));
 sky130_fd_sc_hd__o21ai_1 _4711_ (.A1(_3049_),
    .A2(_0327_),
    .B1(_1219_),
    .Y(_1220_));
 sky130_fd_sc_hd__a221oi_1 _4712_ (.A1(_3062_),
    .A2(_3340_),
    .B1(_3094_),
    .B2(_0323_),
    .C1(_1220_),
    .Y(_1221_));
 sky130_fd_sc_hd__and4_1 _4713_ (.A(_1210_),
    .B(_1214_),
    .C(_1218_),
    .D(_1221_),
    .X(_1222_));
 sky130_fd_sc_hd__nand2_1 _4714_ (.A(_3039_),
    .B(_0716_),
    .Y(_1223_));
 sky130_fd_sc_hd__nand2_1 _4715_ (.A(_3060_),
    .B(\egd_top.BitStream_buffer.BS_buffer[104] ),
    .Y(_1224_));
 sky130_fd_sc_hd__nand2_1 _4716_ (.A(_3048_),
    .B(_3100_),
    .Y(_1225_));
 sky130_fd_sc_hd__o2111a_1 _4717_ (.A1(_3085_),
    .A2(_3056_),
    .B1(_1223_),
    .C1(_1224_),
    .D1(_1225_),
    .X(_1226_));
 sky130_fd_sc_hd__nand2_1 _4718_ (.A(_3098_),
    .B(_3118_),
    .Y(_1227_));
 sky130_fd_sc_hd__nand2_1 _4719_ (.A(_3092_),
    .B(_0722_),
    .Y(_1228_));
 sky130_fd_sc_hd__or2_1 _4720_ (.A(_1025_),
    .B(_3088_),
    .X(_1229_));
 sky130_fd_sc_hd__o2111a_1 _4721_ (.A1(_0721_),
    .A2(_3106_),
    .B1(_1227_),
    .C1(_1228_),
    .D1(_1229_),
    .X(_1230_));
 sky130_fd_sc_hd__nand2_1 _4722_ (.A(_3126_),
    .B(_3070_),
    .Y(_1231_));
 sky130_fd_sc_hd__nand2_1 _4723_ (.A(_3112_),
    .B(_3082_),
    .Y(_1232_));
 sky130_fd_sc_hd__nand2_1 _4724_ (.A(_3116_),
    .B(_3169_),
    .Y(_1233_));
 sky130_fd_sc_hd__o2111a_1 _4725_ (.A1(_0808_),
    .A2(_3122_),
    .B1(_1231_),
    .C1(_1232_),
    .D1(_1233_),
    .X(_1234_));
 sky130_fd_sc_hd__nand2_1 _4726_ (.A(_3073_),
    .B(\egd_top.BitStream_buffer.BS_buffer[114] ),
    .Y(_1235_));
 sky130_fd_sc_hd__o21ai_1 _4727_ (.A1(_2980_),
    .A2(_0729_),
    .B1(_1235_),
    .Y(_1236_));
 sky130_fd_sc_hd__a221oi_1 _4728_ (.A1(_3157_),
    .A2(_0726_),
    .B1(_3204_),
    .B2(_3081_),
    .C1(_1236_),
    .Y(_1237_));
 sky130_fd_sc_hd__and4_1 _4729_ (.A(_1226_),
    .B(_1230_),
    .C(_1234_),
    .D(_1237_),
    .X(_1238_));
 sky130_fd_sc_hd__nand2_1 _4730_ (.A(_3175_),
    .B(\egd_top.BitStream_buffer.BS_buffer[1] ),
    .Y(_1239_));
 sky130_fd_sc_hd__nand2_1 _4731_ (.A(_3179_),
    .B(_0930_),
    .Y(_1240_));
 sky130_fd_sc_hd__nand2_1 _4732_ (.A(_3185_),
    .B(\egd_top.BitStream_buffer.BS_buffer[4] ),
    .Y(_1241_));
 sky130_fd_sc_hd__o2111a_1 _4733_ (.A1(_0597_),
    .A2(_3182_),
    .B1(_1239_),
    .C1(_1240_),
    .D1(_1241_),
    .X(_1242_));
 sky130_fd_sc_hd__nand2_1 _4734_ (.A(_3140_),
    .B(\egd_top.BitStream_buffer.BS_buffer[0] ),
    .Y(_1243_));
 sky130_fd_sc_hd__nand2_1 _4735_ (.A(_3147_),
    .B(\egd_top.BitStream_buffer.BS_buffer[126] ),
    .Y(_1244_));
 sky130_fd_sc_hd__nand2_1 _4736_ (.A(_3136_),
    .B(\egd_top.BitStream_buffer.BS_buffer[127] ),
    .Y(_1245_));
 sky130_fd_sc_hd__and3_1 _4737_ (.A(_1243_),
    .B(_1244_),
    .C(_1245_),
    .X(_1246_));
 sky130_fd_sc_hd__o211a_1 _4738_ (.A1(_3018_),
    .A2(_3145_),
    .B1(_1242_),
    .C1(_1246_),
    .X(_1247_));
 sky130_fd_sc_hd__nand2_1 _4739_ (.A(_3163_),
    .B(_3191_),
    .Y(_1248_));
 sky130_fd_sc_hd__nand2_1 _4740_ (.A(_3168_),
    .B(\egd_top.BitStream_buffer.BS_buffer[117] ),
    .Y(_1249_));
 sky130_fd_sc_hd__nand2_1 _4741_ (.A(_1248_),
    .B(_1249_),
    .Y(_1250_));
 sky130_fd_sc_hd__a221oi_2 _4742_ (.A1(_3198_),
    .A2(_3156_),
    .B1(_0744_),
    .B2(_3160_),
    .C1(_1250_),
    .Y(_1251_));
 sky130_fd_sc_hd__nand2_1 _4743_ (.A(_3203_),
    .B(_3149_),
    .Y(_1252_));
 sky130_fd_sc_hd__o21ai_1 _4744_ (.A1(_3009_),
    .A2(_3200_),
    .B1(_1252_),
    .Y(_1253_));
 sky130_fd_sc_hd__a221oi_1 _4745_ (.A1(\egd_top.BitStream_buffer.BS_buffer[123] ),
    .A2(_3194_),
    .B1(_3197_),
    .B2(_3173_),
    .C1(_1253_),
    .Y(_1254_));
 sky130_fd_sc_hd__and3_1 _4746_ (.A(_1247_),
    .B(_1251_),
    .C(_1254_),
    .X(_1255_));
 sky130_fd_sc_hd__nand2_1 _4747_ (.A(_3223_),
    .B(_3252_),
    .Y(_1256_));
 sky130_fd_sc_hd__o21ai_1 _4748_ (.A1(_1149_),
    .A2(_1145_),
    .B1(_1256_),
    .Y(_1257_));
 sky130_fd_sc_hd__a221oi_1 _4749_ (.A1(_3264_),
    .A2(_3215_),
    .B1(_3248_),
    .B2(_3220_),
    .C1(_1257_),
    .Y(_1258_));
 sky130_fd_sc_hd__nand2_1 _4750_ (.A(_3242_),
    .B(_3217_),
    .Y(_1259_));
 sky130_fd_sc_hd__nand2_1 _4751_ (.A(_3232_),
    .B(\egd_top.BitStream_buffer.BS_buffer[71] ),
    .Y(_1260_));
 sky130_fd_sc_hd__nand2_1 _4752_ (.A(_3235_),
    .B(_3256_),
    .Y(_1261_));
 sky130_fd_sc_hd__o2111a_1 _4753_ (.A1(_0755_),
    .A2(_3239_),
    .B1(_1259_),
    .C1(_1260_),
    .D1(_1261_),
    .X(_1262_));
 sky130_fd_sc_hd__nand2_1 _4754_ (.A(_3254_),
    .B(\egd_top.BitStream_buffer.BS_buffer[80] ),
    .Y(_1263_));
 sky130_fd_sc_hd__nand2_1 _4755_ (.A(_3262_),
    .B(\egd_top.BitStream_buffer.BS_buffer[78] ),
    .Y(_1264_));
 sky130_fd_sc_hd__nand2_1 _4756_ (.A(_3250_),
    .B(\egd_top.BitStream_buffer.BS_buffer[79] ),
    .Y(_1265_));
 sky130_fd_sc_hd__nand2_1 _4757_ (.A(_3259_),
    .B(\egd_top.BitStream_buffer.BS_buffer[77] ),
    .Y(_1266_));
 sky130_fd_sc_hd__and4_1 _4758_ (.A(_1263_),
    .B(_1264_),
    .C(_1265_),
    .D(_1266_),
    .X(_1267_));
 sky130_fd_sc_hd__nand2_1 _4759_ (.A(_3281_),
    .B(\egd_top.BitStream_buffer.BS_buffer[83] ),
    .Y(_1268_));
 sky130_fd_sc_hd__o21ai_1 _4760_ (.A1(_1158_),
    .A2(_3279_),
    .B1(_1268_),
    .Y(_1269_));
 sky130_fd_sc_hd__a221oi_1 _4761_ (.A1(_3302_),
    .A2(_3270_),
    .B1(_3288_),
    .B2(_3274_),
    .C1(_1269_),
    .Y(_1270_));
 sky130_fd_sc_hd__and4_1 _4762_ (.A(_1258_),
    .B(_1262_),
    .C(_1267_),
    .D(_1270_),
    .X(_1271_));
 sky130_fd_sc_hd__and4_1 _4763_ (.A(_1222_),
    .B(_1238_),
    .C(_1255_),
    .D(_1271_),
    .X(_1272_));
 sky130_fd_sc_hd__nand2_1 _4764_ (.A(_0353_),
    .B(_0869_),
    .Y(_1273_));
 sky130_fd_sc_hd__o21ai_1 _4765_ (.A1(_0637_),
    .A2(_0350_),
    .B1(_1273_),
    .Y(_1274_));
 sky130_fd_sc_hd__a221oi_1 _4766_ (.A1(_0379_),
    .A2(_0342_),
    .B1(_0345_),
    .B2(_0389_),
    .C1(_1274_),
    .Y(_1275_));
 sky130_fd_sc_hd__clkinv_2 _4767_ (.A(_0354_),
    .Y(_1276_));
 sky130_fd_sc_hd__nand2_1 _4768_ (.A(_0371_),
    .B(_0346_),
    .Y(_1277_));
 sky130_fd_sc_hd__o21ai_1 _4769_ (.A1(_1276_),
    .A2(_0368_),
    .B1(_1277_),
    .Y(_1278_));
 sky130_fd_sc_hd__a221oi_1 _4770_ (.A1(_0347_),
    .A2(_0360_),
    .B1(_0363_),
    .B2(_0375_),
    .C1(_1278_),
    .Y(_1279_));
 sky130_fd_sc_hd__nand2_1 _4771_ (.A(_0387_),
    .B(_0642_),
    .Y(_1280_));
 sky130_fd_sc_hd__o21ai_1 _4772_ (.A1(_0423_),
    .A2(_0385_),
    .B1(_1280_),
    .Y(_1281_));
 sky130_fd_sc_hd__a221oi_1 _4773_ (.A1(_0400_),
    .A2(_0378_),
    .B1(_0407_),
    .B2(_0382_),
    .C1(_1281_),
    .Y(_1282_));
 sky130_fd_sc_hd__nand2_1 _4774_ (.A(_0406_),
    .B(_0416_),
    .Y(_1283_));
 sky130_fd_sc_hd__o21ai_1 _4775_ (.A1(_0960_),
    .A2(_0403_),
    .B1(_1283_),
    .Y(_1284_));
 sky130_fd_sc_hd__a221oi_1 _4776_ (.A1(_0948_),
    .A2(_0396_),
    .B1(_0399_),
    .B2(_0412_),
    .C1(_1284_),
    .Y(_1285_));
 sky130_fd_sc_hd__and4_1 _4777_ (.A(_1275_),
    .B(_1279_),
    .C(_1282_),
    .D(_1285_),
    .X(_1286_));
 sky130_fd_sc_hd__or2_1 _4778_ (.A(_0437_),
    .B(_0425_),
    .X(_1287_));
 sky130_fd_sc_hd__o21ai_1 _4779_ (.A1(_0653_),
    .A2(_0422_),
    .B1(_1287_),
    .Y(_1288_));
 sky130_fd_sc_hd__a221oi_1 _4780_ (.A1(_0436_),
    .A2(_0415_),
    .B1(_0454_),
    .B2(_0419_),
    .C1(_1288_),
    .Y(_1289_));
 sky130_fd_sc_hd__nand2_1 _4781_ (.A(_0453_),
    .B(_0471_),
    .Y(_1290_));
 sky130_fd_sc_hd__nand2_1 _4782_ (.A(_0458_),
    .B(_0664_),
    .Y(_1291_));
 sky130_fd_sc_hd__or2_1 _4783_ (.A(_0955_),
    .B(_0464_),
    .X(_1292_));
 sky130_fd_sc_hd__o2111a_1 _4784_ (.A1(_0663_),
    .A2(_0450_),
    .B1(_1290_),
    .C1(_1291_),
    .D1(_1292_),
    .X(_1293_));
 sky130_fd_sc_hd__a22o_1 _4785_ (.A1(_0447_),
    .A2(_0431_),
    .B1(_0435_),
    .B2(_0467_),
    .X(_1294_));
 sky130_fd_sc_hd__a32o_1 _4786_ (.A1(_3104_),
    .A2(_0459_),
    .A3(_2934_),
    .B1(_0461_),
    .B2(_0442_),
    .X(_1295_));
 sky130_fd_sc_hd__nor2_1 _4787_ (.A(_1294_),
    .B(_1295_),
    .Y(_1296_));
 sky130_fd_sc_hd__clkinv_2 _4788_ (.A(\egd_top.BitStream_buffer.BS_buffer[66] ),
    .Y(_1297_));
 sky130_fd_sc_hd__nand2_1 _4789_ (.A(_0469_),
    .B(_0751_),
    .Y(_1298_));
 sky130_fd_sc_hd__o21ai_1 _4790_ (.A1(_1297_),
    .A2(_0472_),
    .B1(_1298_),
    .Y(_1299_));
 sky130_fd_sc_hd__a221oi_1 _4791_ (.A1(_3237_),
    .A2(_0477_),
    .B1(_3210_),
    .B2(_2936_),
    .C1(_1299_),
    .Y(_1300_));
 sky130_fd_sc_hd__and4_1 _4792_ (.A(_1289_),
    .B(_1293_),
    .C(_1296_),
    .D(_1300_),
    .X(_1301_));
 sky130_fd_sc_hd__nand2_1 _4793_ (.A(_1286_),
    .B(_1301_),
    .Y(_1302_));
 sky130_fd_sc_hd__nand2_1 _4794_ (.A(_0497_),
    .B(_0519_),
    .Y(_1303_));
 sky130_fd_sc_hd__o21ai_1 _4795_ (.A1(_0510_),
    .A2(_0495_),
    .B1(_1303_),
    .Y(_1304_));
 sky130_fd_sc_hd__a221oi_1 _4796_ (.A1(_0505_),
    .A2(_0487_),
    .B1(_0515_),
    .B2(_0490_),
    .C1(_1304_),
    .Y(_1305_));
 sky130_fd_sc_hd__nand2_1 _4797_ (.A(_0514_),
    .B(\egd_top.BitStream_buffer.BS_buffer[27] ),
    .Y(_1306_));
 sky130_fd_sc_hd__o21ai_1 _4798_ (.A1(_0699_),
    .A2(_0512_),
    .B1(_1306_),
    .Y(_1307_));
 sky130_fd_sc_hd__a221oi_1 _4799_ (.A1(_0527_),
    .A2(_0504_),
    .B1(_0531_),
    .B2(_0508_),
    .C1(_1307_),
    .Y(_1308_));
 sky130_fd_sc_hd__o22a_1 _4800_ (.A1(_0702_),
    .A2(_0530_),
    .B1(_0995_),
    .B2(_0526_),
    .X(_1309_));
 sky130_fd_sc_hd__o221a_1 _4801_ (.A1(_0543_),
    .A2(_0523_),
    .B1(_0907_),
    .B2(_0534_),
    .C1(_1309_),
    .X(_1310_));
 sky130_fd_sc_hd__nand2_1 _4802_ (.A(_0548_),
    .B(_0365_),
    .Y(_1311_));
 sky130_fd_sc_hd__o21ai_1 _4803_ (.A1(_0633_),
    .A2(_0546_),
    .B1(_1311_),
    .Y(_1312_));
 sky130_fd_sc_hd__a221oi_1 _4804_ (.A1(_0364_),
    .A2(_0539_),
    .B1(_0337_),
    .B2(_0542_),
    .C1(_1312_),
    .Y(_1313_));
 sky130_fd_sc_hd__and4_1 _4805_ (.A(_1305_),
    .B(_1308_),
    .C(_1310_),
    .D(_1313_),
    .X(_1314_));
 sky130_fd_sc_hd__nand2_1 _4806_ (.A(_0561_),
    .B(\egd_top.BitStream_buffer.BS_buffer[11] ),
    .Y(_1315_));
 sky130_fd_sc_hd__nand2_1 _4807_ (.A(_0565_),
    .B(_0585_),
    .Y(_1316_));
 sky130_fd_sc_hd__or2_1 _4808_ (.A(_0679_),
    .B(_0571_),
    .X(_1317_));
 sky130_fd_sc_hd__o2111a_1 _4809_ (.A1(_0676_),
    .A2(_0558_),
    .B1(_1315_),
    .C1(_1316_),
    .D1(_1317_),
    .X(_1318_));
 sky130_fd_sc_hd__nand2_1 _4810_ (.A(_0582_),
    .B(\egd_top.BitStream_buffer.BS_buffer[15] ),
    .Y(_1319_));
 sky130_fd_sc_hd__nand2_1 _4811_ (.A(_0578_),
    .B(\egd_top.BitStream_buffer.BS_buffer[13] ),
    .Y(_1320_));
 sky130_fd_sc_hd__or2_1 _4812_ (.A(_0685_),
    .B(_0575_),
    .X(_1321_));
 sky130_fd_sc_hd__o2111a_1 _4813_ (.A1(_0688_),
    .A2(_0588_),
    .B1(_1319_),
    .C1(_1320_),
    .D1(_1321_),
    .X(_1322_));
 sky130_fd_sc_hd__or2_1 _4814_ (.A(_0670_),
    .B(_0599_),
    .X(_1323_));
 sky130_fd_sc_hd__o221a_1 _4815_ (.A1(_0554_),
    .A2(_0593_),
    .B1(_0673_),
    .B2(_0596_),
    .C1(_1323_),
    .X(_1324_));
 sky130_fd_sc_hd__nand2_1 _4816_ (.A(_0606_),
    .B(\egd_top.BitStream_buffer.BS_buffer[17] ),
    .Y(_1325_));
 sky130_fd_sc_hd__nand2_1 _4817_ (.A(_0609_),
    .B(_0498_),
    .Y(_1326_));
 sky130_fd_sc_hd__or2_1 _4818_ (.A(_0897_),
    .B(_0603_),
    .X(_1327_));
 sky130_fd_sc_hd__o2111a_1 _4819_ (.A1(_0492_),
    .A2(_0613_),
    .B1(_1325_),
    .C1(_1326_),
    .D1(_1327_),
    .X(_1328_));
 sky130_fd_sc_hd__and4_1 _4820_ (.A(_1318_),
    .B(_1322_),
    .C(_1324_),
    .D(_1328_),
    .X(_1329_));
 sky130_fd_sc_hd__nand2_1 _4821_ (.A(_1314_),
    .B(_1329_),
    .Y(_1330_));
 sky130_fd_sc_hd__nor2_1 _4822_ (.A(_1302_),
    .B(_1330_),
    .Y(_1331_));
 sky130_fd_sc_hd__nand2_1 _4823_ (.A(_0622_),
    .B(_0568_),
    .Y(_1332_));
 sky130_fd_sc_hd__nand3_1 _4824_ (.A(_1272_),
    .B(_1331_),
    .C(_1332_),
    .Y(_1333_));
 sky130_fd_sc_hd__nor2_1 _4825_ (.A(_3026_),
    .B(_1333_),
    .Y(_1334_));
 sky130_fd_sc_hd__nor2_1 _4826_ (.A(_1207_),
    .B(_1334_),
    .Y(_0292_));
 sky130_fd_sc_hd__o21ai_1 _4827_ (.A1(\egd_top.BitStream_buffer.BitStream_buffer_output[9] ),
    .A2(_2965_),
    .B1(_0627_),
    .Y(_1335_));
 sky130_fd_sc_hd__nand2_1 _4828_ (.A(_0353_),
    .B(_0393_),
    .Y(_1336_));
 sky130_fd_sc_hd__o21ai_1 _4829_ (.A1(_0870_),
    .A2(_0350_),
    .B1(_1336_),
    .Y(_1337_));
 sky130_fd_sc_hd__a221oi_1 _4830_ (.A1(_0389_),
    .A2(_0342_),
    .B1(_0345_),
    .B2(_0869_),
    .C1(_1337_),
    .Y(_1338_));
 sky130_fd_sc_hd__nand2_1 _4831_ (.A(_0370_),
    .B(_0354_),
    .Y(_1339_));
 sky130_fd_sc_hd__o21ai_1 _4832_ (.A1(_0348_),
    .A2(_0367_),
    .B1(_1339_),
    .Y(_1340_));
 sky130_fd_sc_hd__a221oi_1 _4833_ (.A1(_0375_),
    .A2(_0359_),
    .B1(_0362_),
    .B2(_0379_),
    .C1(_1340_),
    .Y(_1341_));
 sky130_fd_sc_hd__nand2_1 _4834_ (.A(_0377_),
    .B(_0407_),
    .Y(_1342_));
 sky130_fd_sc_hd__o21ai_1 _4835_ (.A1(_0401_),
    .A2(_0380_),
    .B1(_1342_),
    .Y(_1343_));
 sky130_fd_sc_hd__a221oi_1 _4836_ (.A1(_0874_),
    .A2(_0388_),
    .B1(_0948_),
    .B2(_0944_),
    .C1(_1343_),
    .Y(_1344_));
 sky130_fd_sc_hd__nand2_1 _4837_ (.A(_0405_),
    .B(_0443_),
    .Y(_1345_));
 sky130_fd_sc_hd__o21ai_1 _4838_ (.A1(_0437_),
    .A2(_0402_),
    .B1(_1345_),
    .Y(_1346_));
 sky130_fd_sc_hd__a221oi_1 _4839_ (.A1(_0412_),
    .A2(_0396_),
    .B1(_0399_),
    .B2(_0416_),
    .C1(_1346_),
    .Y(_1347_));
 sky130_fd_sc_hd__and4_1 _4840_ (.A(_1338_),
    .B(_1341_),
    .C(_1344_),
    .D(_1347_),
    .X(_1348_));
 sky130_fd_sc_hd__or2_1 _4841_ (.A(_0653_),
    .B(_0424_),
    .X(_1349_));
 sky130_fd_sc_hd__o21ai_1 _4842_ (.A1(_0883_),
    .A2(_0422_),
    .B1(_1349_),
    .Y(_1350_));
 sky130_fd_sc_hd__a221oi_1 _4843_ (.A1(_0454_),
    .A2(_0415_),
    .B1(_0461_),
    .B2(_0419_),
    .C1(_1350_),
    .Y(_1351_));
 sky130_fd_sc_hd__nand2_1 _4844_ (.A(_0452_),
    .B(_0478_),
    .Y(_1352_));
 sky130_fd_sc_hd__nand2_1 _4845_ (.A(_0457_),
    .B(_3244_),
    .Y(_1353_));
 sky130_fd_sc_hd__or2_1 _4846_ (.A(_0474_),
    .B(_0463_),
    .X(_1354_));
 sky130_fd_sc_hd__o2111a_1 _4847_ (.A1(_3238_),
    .A2(_0450_),
    .B1(_1352_),
    .C1(_1353_),
    .D1(_1354_),
    .X(_1355_));
 sky130_fd_sc_hd__nand2_1 _4848_ (.A(_0441_),
    .B(_0459_),
    .Y(_1356_));
 sky130_fd_sc_hd__nand2_1 _4849_ (.A(_0432_),
    .B(_0467_),
    .Y(_1357_));
 sky130_fd_sc_hd__nand2_1 _4850_ (.A(_0435_),
    .B(_0471_),
    .Y(_1358_));
 sky130_fd_sc_hd__o2111a_1 _4851_ (.A1(_0448_),
    .A2(_0439_),
    .B1(_1356_),
    .C1(_1357_),
    .D1(_1358_),
    .X(_1359_));
 sky130_fd_sc_hd__inv_2 _4852_ (.A(\egd_top.BitStream_buffer.BS_buffer[69] ),
    .Y(_1360_));
 sky130_fd_sc_hd__nand2_1 _4853_ (.A(_0476_),
    .B(\egd_top.BitStream_buffer.BS_buffer[68] ),
    .Y(_1361_));
 sky130_fd_sc_hd__o21ai_1 _4854_ (.A1(_1360_),
    .A2(_2935_),
    .B1(_1361_),
    .Y(_1362_));
 sky130_fd_sc_hd__a221oi_1 _4855_ (.A1(_3230_),
    .A2(_0470_),
    .B1(_3237_),
    .B2(_0473_),
    .C1(_1362_),
    .Y(_1363_));
 sky130_fd_sc_hd__and4_1 _4856_ (.A(_1351_),
    .B(_1355_),
    .C(_1359_),
    .D(_1363_),
    .X(_1364_));
 sky130_fd_sc_hd__nand2_1 _4857_ (.A(_0564_),
    .B(_0583_),
    .Y(_1365_));
 sky130_fd_sc_hd__nand2_1 _4858_ (.A(_0560_),
    .B(\egd_top.BitStream_buffer.BS_buffer[12] ),
    .Y(_1366_));
 sky130_fd_sc_hd__or2_1 _4859_ (.A(_0574_),
    .B(_0570_),
    .X(_1367_));
 sky130_fd_sc_hd__o2111a_1 _4860_ (.A1(_0611_),
    .A2(_0557_),
    .B1(_1365_),
    .C1(_1366_),
    .D1(_1367_),
    .X(_1368_));
 sky130_fd_sc_hd__nand2_1 _4861_ (.A(_0581_),
    .B(\egd_top.BitStream_buffer.BS_buffer[16] ),
    .Y(_1369_));
 sky130_fd_sc_hd__nand2_1 _4862_ (.A(_0577_),
    .B(\egd_top.BitStream_buffer.BS_buffer[14] ),
    .Y(_1370_));
 sky130_fd_sc_hd__or2_1 _4863_ (.A(_0602_),
    .B(_0587_),
    .X(_1371_));
 sky130_fd_sc_hd__o2111a_1 _4864_ (.A1(_0922_),
    .A2(_0575_),
    .B1(_1369_),
    .C1(_1370_),
    .D1(_1371_),
    .X(_1372_));
 sky130_fd_sc_hd__or2_1 _4865_ (.A(_0586_),
    .B(_0598_),
    .X(_1373_));
 sky130_fd_sc_hd__o221a_1 _4866_ (.A1(_0670_),
    .A2(_0592_),
    .B1(_0554_),
    .B2(_0596_),
    .C1(_1373_),
    .X(_1374_));
 sky130_fd_sc_hd__nand2_1 _4867_ (.A(_0608_),
    .B(_0502_),
    .Y(_1375_));
 sky130_fd_sc_hd__nand2_1 _4868_ (.A(_0605_),
    .B(_0491_),
    .Y(_1376_));
 sky130_fd_sc_hd__or2_1 _4869_ (.A(_0692_),
    .B(_0612_),
    .X(_1377_));
 sky130_fd_sc_hd__o2111a_1 _4870_ (.A1(_0986_),
    .A2(_0603_),
    .B1(_1375_),
    .C1(_1376_),
    .D1(_1377_),
    .X(_1378_));
 sky130_fd_sc_hd__and4_1 _4871_ (.A(_1368_),
    .B(_1372_),
    .C(_1374_),
    .D(_1378_),
    .X(_1379_));
 sky130_fd_sc_hd__nand2_1 _4872_ (.A(_0486_),
    .B(_0515_),
    .Y(_1380_));
 sky130_fd_sc_hd__nand2_1 _4873_ (.A(_0489_),
    .B(_0509_),
    .Y(_1381_));
 sky130_fd_sc_hd__nand2_1 _4874_ (.A(_0496_),
    .B(_0527_),
    .Y(_1382_));
 sky130_fd_sc_hd__o2111a_1 _4875_ (.A1(_0520_),
    .A2(_0494_),
    .B1(_1380_),
    .C1(_1381_),
    .D1(_1382_),
    .X(_1383_));
 sky130_fd_sc_hd__nand2_1 _4876_ (.A(_0503_),
    .B(_0531_),
    .Y(_1384_));
 sky130_fd_sc_hd__nand2_1 _4877_ (.A(_0513_),
    .B(\egd_top.BitStream_buffer.BS_buffer[28] ),
    .Y(_1385_));
 sky130_fd_sc_hd__nand2_1 _4878_ (.A(_0507_),
    .B(\egd_top.BitStream_buffer.BS_buffer[27] ),
    .Y(_1386_));
 sky130_fd_sc_hd__o2111a_1 _4879_ (.A1(_0543_),
    .A2(_0512_),
    .B1(_1384_),
    .C1(_1385_),
    .D1(_1386_),
    .X(_1387_));
 sky130_fd_sc_hd__nand2_1 _4880_ (.A(_0547_),
    .B(\egd_top.BitStream_buffer.BS_buffer[34] ),
    .Y(_1388_));
 sky130_fd_sc_hd__o21ai_1 _4881_ (.A1(_0865_),
    .A2(_0545_),
    .B1(_1388_),
    .Y(_1389_));
 sky130_fd_sc_hd__a221oi_1 _4882_ (.A1(_0337_),
    .A2(_0538_),
    .B1(_0346_),
    .B2(_0541_),
    .C1(_1389_),
    .Y(_1390_));
 sky130_fd_sc_hd__o22a_1 _4883_ (.A1(_0907_),
    .A2(_0529_),
    .B1(_0995_),
    .B2(_0533_),
    .X(_1391_));
 sky130_fd_sc_hd__o221a_1 _4884_ (.A1(_0702_),
    .A2(_0522_),
    .B1(_0366_),
    .B2(_0525_),
    .C1(_1391_),
    .X(_1392_));
 sky130_fd_sc_hd__and4_1 _4885_ (.A(_1383_),
    .B(_1387_),
    .C(_1390_),
    .D(_1392_),
    .X(_1393_));
 sky130_fd_sc_hd__and4_1 _4886_ (.A(_1348_),
    .B(_1364_),
    .C(_1379_),
    .D(_1393_),
    .X(_1394_));
 sky130_fd_sc_hd__nand2_1 _4887_ (.A(_3332_),
    .B(_3338_),
    .Y(_1395_));
 sky130_fd_sc_hd__o21ai_1 _4888_ (.A1(_0854_),
    .A2(_3329_),
    .B1(_1395_),
    .Y(_1396_));
 sky130_fd_sc_hd__a221oi_1 _4889_ (.A1(_3028_),
    .A2(_3323_),
    .B1(_3325_),
    .B2(_3040_),
    .C1(_1396_),
    .Y(_1397_));
 sky130_fd_sc_hd__nand2_1 _4890_ (.A(_3291_),
    .B(\egd_top.BitStream_buffer.BS_buffer[88] ),
    .Y(_1398_));
 sky130_fd_sc_hd__nand2_1 _4891_ (.A(_3300_),
    .B(_0772_),
    .Y(_1399_));
 sky130_fd_sc_hd__nand2_1 _4892_ (.A(_3294_),
    .B(_0780_),
    .Y(_1400_));
 sky130_fd_sc_hd__o2111a_1 _4893_ (.A1(_0771_),
    .A2(_3298_),
    .B1(_1398_),
    .C1(_1399_),
    .D1(_1400_),
    .X(_1401_));
 sky130_fd_sc_hd__nand2_1 _4894_ (.A(_3313_),
    .B(_3322_),
    .Y(_1402_));
 sky130_fd_sc_hd__nand2_1 _4895_ (.A(_3309_),
    .B(_0330_),
    .Y(_1403_));
 sky130_fd_sc_hd__or2_1 _4896_ (.A(_0324_),
    .B(_3307_),
    .X(_1404_));
 sky130_fd_sc_hd__o2111a_1 _4897_ (.A1(_0850_),
    .A2(_3319_),
    .B1(_1402_),
    .C1(_1403_),
    .D1(_1404_),
    .X(_1405_));
 sky130_fd_sc_hd__nand2_1 _4898_ (.A(_0328_),
    .B(_0708_),
    .Y(_1406_));
 sky130_fd_sc_hd__o21ai_1 _4899_ (.A1(_0709_),
    .A2(_0326_),
    .B1(_1406_),
    .Y(_1407_));
 sky130_fd_sc_hd__a221oi_1 _4900_ (.A1(_3094_),
    .A2(_3339_),
    .B1(_0716_),
    .B2(_0322_),
    .C1(_1407_),
    .Y(_1408_));
 sky130_fd_sc_hd__and4_1 _4901_ (.A(_1397_),
    .B(_1401_),
    .C(_1405_),
    .D(_1408_),
    .X(_1409_));
 sky130_fd_sc_hd__nand2_1 _4902_ (.A(_3038_),
    .B(\egd_top.BitStream_buffer.BS_buffer[102] ),
    .Y(_1410_));
 sky130_fd_sc_hd__nand2_1 _4903_ (.A(_3047_),
    .B(_0714_),
    .Y(_1411_));
 sky130_fd_sc_hd__nand2_1 _4904_ (.A(_3060_),
    .B(_0722_),
    .Y(_1412_));
 sky130_fd_sc_hd__o2111a_1 _4905_ (.A1(_0718_),
    .A2(_3055_),
    .B1(_1410_),
    .C1(_1411_),
    .D1(_1412_),
    .X(_1413_));
 sky130_fd_sc_hd__nand2_1 _4906_ (.A(_3092_),
    .B(_3109_),
    .Y(_1414_));
 sky130_fd_sc_hd__nand2_1 _4907_ (.A(_3098_),
    .B(\egd_top.BitStream_buffer.BS_buffer[108] ),
    .Y(_1415_));
 sky130_fd_sc_hd__or2_1 _4908_ (.A(_0804_),
    .B(_3105_),
    .X(_1416_));
 sky130_fd_sc_hd__o2111a_1 _4909_ (.A1(_0727_),
    .A2(_3089_),
    .B1(_1414_),
    .C1(_1415_),
    .D1(_1416_),
    .X(_1417_));
 sky130_fd_sc_hd__nand2_1 _4910_ (.A(_3126_),
    .B(_3075_),
    .Y(_1418_));
 sky130_fd_sc_hd__nand2_1 _4911_ (.A(_3112_),
    .B(_3169_),
    .Y(_1419_));
 sky130_fd_sc_hd__nand2_1 _4912_ (.A(_3116_),
    .B(_3164_),
    .Y(_1420_));
 sky130_fd_sc_hd__o2111a_1 _4913_ (.A1(_1035_),
    .A2(_3122_),
    .B1(_1418_),
    .C1(_1419_),
    .D1(_1420_),
    .X(_1421_));
 sky130_fd_sc_hd__nand2_1 _4914_ (.A(_3073_),
    .B(_3157_),
    .Y(_1422_));
 sky130_fd_sc_hd__o21ai_1 _4915_ (.A1(_2983_),
    .A2(_0728_),
    .B1(_1422_),
    .Y(_1423_));
 sky130_fd_sc_hd__a221oi_1 _4916_ (.A1(_3204_),
    .A2(_3078_),
    .B1(_0746_),
    .B2(_3080_),
    .C1(_1423_),
    .Y(_1424_));
 sky130_fd_sc_hd__and4_1 _4917_ (.A(_1413_),
    .B(_1417_),
    .C(_1421_),
    .D(_1424_),
    .X(_1425_));
 sky130_fd_sc_hd__inv_2 _4918_ (.A(\egd_top.BitStream_buffer.BS_buffer[77] ),
    .Y(_1426_));
 sky130_fd_sc_hd__nand2_1 _4919_ (.A(_3223_),
    .B(\egd_top.BitStream_buffer.BS_buffer[76] ),
    .Y(_1427_));
 sky130_fd_sc_hd__o21ai_1 _4920_ (.A1(_1426_),
    .A2(_1145_),
    .B1(_1427_),
    .Y(_1428_));
 sky130_fd_sc_hd__a221oi_1 _4921_ (.A1(_3248_),
    .A2(_3215_),
    .B1(_3252_),
    .B2(_3219_),
    .C1(_1428_),
    .Y(_1429_));
 sky130_fd_sc_hd__inv_2 _4922_ (.A(\egd_top.BitStream_buffer.BS_buffer[71] ),
    .Y(_1430_));
 sky130_fd_sc_hd__nand2_1 _4923_ (.A(_3242_),
    .B(\egd_top.BitStream_buffer.BS_buffer[70] ),
    .Y(_1431_));
 sky130_fd_sc_hd__nand2_1 _4924_ (.A(_3232_),
    .B(_3256_),
    .Y(_1432_));
 sky130_fd_sc_hd__nand2_1 _4925_ (.A(_3235_),
    .B(_3264_),
    .Y(_1433_));
 sky130_fd_sc_hd__o2111a_1 _4926_ (.A1(_1430_),
    .A2(_3239_),
    .B1(_1431_),
    .C1(_1432_),
    .D1(_1433_),
    .X(_1434_));
 sky130_fd_sc_hd__nand2_1 _4927_ (.A(_3262_),
    .B(\egd_top.BitStream_buffer.BS_buffer[79] ),
    .Y(_1435_));
 sky130_fd_sc_hd__nand2_1 _4928_ (.A(_3254_),
    .B(_3302_),
    .Y(_1436_));
 sky130_fd_sc_hd__nand2_1 _4929_ (.A(_3259_),
    .B(\egd_top.BitStream_buffer.BS_buffer[78] ),
    .Y(_1437_));
 sky130_fd_sc_hd__nand2_1 _4930_ (.A(_3250_),
    .B(\egd_top.BitStream_buffer.BS_buffer[80] ),
    .Y(_1438_));
 sky130_fd_sc_hd__and4_1 _4931_ (.A(_1435_),
    .B(_1436_),
    .C(_1437_),
    .D(_1438_),
    .X(_1439_));
 sky130_fd_sc_hd__nand2_1 _4932_ (.A(_3270_),
    .B(\egd_top.BitStream_buffer.BS_buffer[82] ),
    .Y(_1440_));
 sky130_fd_sc_hd__o21ai_1 _4933_ (.A1(_1007_),
    .A2(_3273_),
    .B1(_1440_),
    .Y(_1441_));
 sky130_fd_sc_hd__a221oi_1 _4934_ (.A1(_3315_),
    .A2(_3282_),
    .B1(_0774_),
    .B2(_1153_),
    .C1(_1441_),
    .Y(_1442_));
 sky130_fd_sc_hd__and4_1 _4935_ (.A(_1429_),
    .B(_1434_),
    .C(_1439_),
    .D(_1442_),
    .X(_1443_));
 sky130_fd_sc_hd__nand2_1 _4936_ (.A(_3193_),
    .B(\egd_top.BitStream_buffer.BS_buffer[124] ),
    .Y(_1444_));
 sky130_fd_sc_hd__nand2_1 _4937_ (.A(_3202_),
    .B(\egd_top.BitStream_buffer.BS_buffer[122] ),
    .Y(_1445_));
 sky130_fd_sc_hd__nand2_1 _4938_ (.A(_3196_),
    .B(_3177_),
    .Y(_1446_));
 sky130_fd_sc_hd__o2111a_1 _4939_ (.A1(_3012_),
    .A2(_3199_),
    .B1(_1444_),
    .C1(_1445_),
    .D1(_1446_),
    .X(_1447_));
 sky130_fd_sc_hd__nand2_1 _4940_ (.A(_3162_),
    .B(\egd_top.BitStream_buffer.BS_buffer[119] ),
    .Y(_1448_));
 sky130_fd_sc_hd__nand2_1 _4941_ (.A(_3159_),
    .B(\egd_top.BitStream_buffer.BS_buffer[121] ),
    .Y(_1449_));
 sky130_fd_sc_hd__nand2_1 _4942_ (.A(_3155_),
    .B(\egd_top.BitStream_buffer.BS_buffer[120] ),
    .Y(_1450_));
 sky130_fd_sc_hd__nand2_1 _4943_ (.A(_3167_),
    .B(\egd_top.BitStream_buffer.BS_buffer[118] ),
    .Y(_1451_));
 sky130_fd_sc_hd__and4_1 _4944_ (.A(_1448_),
    .B(_1449_),
    .C(_1450_),
    .D(_1451_),
    .X(_1452_));
 sky130_fd_sc_hd__nand2_1 _4945_ (.A(_3147_),
    .B(\egd_top.BitStream_buffer.BS_buffer[127] ),
    .Y(_1453_));
 sky130_fd_sc_hd__nand2_1 _4946_ (.A(_3140_),
    .B(\egd_top.BitStream_buffer.BS_buffer[1] ),
    .Y(_1454_));
 sky130_fd_sc_hd__nand2_1 _4947_ (.A(_3136_),
    .B(\egd_top.BitStream_buffer.BS_buffer[0] ),
    .Y(_1455_));
 sky130_fd_sc_hd__nand2_1 _4948_ (.A(_3144_),
    .B(\egd_top.BitStream_buffer.BS_buffer[126] ),
    .Y(_1456_));
 sky130_fd_sc_hd__and4_1 _4949_ (.A(_1453_),
    .B(_1454_),
    .C(_1455_),
    .D(_1456_),
    .X(_1457_));
 sky130_fd_sc_hd__nand2_1 _4950_ (.A(_3185_),
    .B(_0568_),
    .Y(_1458_));
 sky130_fd_sc_hd__o21ai_1 _4951_ (.A1(_0682_),
    .A2(_3183_),
    .B1(_1458_),
    .Y(_1459_));
 sky130_fd_sc_hd__a221oi_1 _4952_ (.A1(_0930_),
    .A2(_3175_),
    .B1(_1076_),
    .B2(_3179_),
    .C1(_1459_),
    .Y(_1460_));
 sky130_fd_sc_hd__and4_1 _4953_ (.A(_1447_),
    .B(_1452_),
    .C(_1457_),
    .D(_1460_),
    .X(_1461_));
 sky130_fd_sc_hd__and4_1 _4954_ (.A(_1409_),
    .B(_1425_),
    .C(_1443_),
    .D(_1461_),
    .X(_1462_));
 sky130_fd_sc_hd__nand2_1 _4955_ (.A(_0622_),
    .B(_0562_),
    .Y(_1463_));
 sky130_fd_sc_hd__nand3_1 _4956_ (.A(_1394_),
    .B(_1462_),
    .C(_1463_),
    .Y(_1464_));
 sky130_fd_sc_hd__nor2_1 _4957_ (.A(_3026_),
    .B(_1464_),
    .Y(_1465_));
 sky130_fd_sc_hd__nor2_1 _4958_ (.A(_1335_),
    .B(_1465_),
    .Y(_0291_));
 sky130_fd_sc_hd__inv_2 _4959_ (.A(\egd_top.BitStream_buffer.BS_buffer[46] ),
    .Y(_1466_));
 sky130_fd_sc_hd__nand2_1 _4960_ (.A(_0353_),
    .B(_0400_),
    .Y(_1467_));
 sky130_fd_sc_hd__o21ai_1 _4961_ (.A1(_1466_),
    .A2(_0350_),
    .B1(_1467_),
    .Y(_1468_));
 sky130_fd_sc_hd__a221oi_1 _4962_ (.A1(_0869_),
    .A2(_0342_),
    .B1(_0345_),
    .B2(_0393_),
    .C1(_1468_),
    .Y(_1469_));
 sky130_fd_sc_hd__nand2_1 _4963_ (.A(_0371_),
    .B(_0347_),
    .Y(_1470_));
 sky130_fd_sc_hd__o21ai_1 _4964_ (.A1(_0629_),
    .A2(_0368_),
    .B1(_1470_),
    .Y(_1471_));
 sky130_fd_sc_hd__a221oi_1 _4965_ (.A1(_0379_),
    .A2(_0360_),
    .B1(_0363_),
    .B2(_0389_),
    .C1(_1471_),
    .Y(_1472_));
 sky130_fd_sc_hd__nand2_1 _4966_ (.A(_0388_),
    .B(_0948_),
    .Y(_1473_));
 sky130_fd_sc_hd__o21ai_1 _4967_ (.A1(_0659_),
    .A2(_0385_),
    .B1(_1473_),
    .Y(_1474_));
 sky130_fd_sc_hd__a221oi_1 _4968_ (.A1(_0642_),
    .A2(_0378_),
    .B1(_0874_),
    .B2(_0382_),
    .C1(_1474_),
    .Y(_1475_));
 sky130_fd_sc_hd__nand2_1 _4969_ (.A(_0406_),
    .B(_0655_),
    .Y(_1476_));
 sky130_fd_sc_hd__o21ai_1 _4970_ (.A1(_0653_),
    .A2(_0403_),
    .B1(_1476_),
    .Y(_1477_));
 sky130_fd_sc_hd__a221oi_1 _4971_ (.A1(_0416_),
    .A2(_0396_),
    .B1(_0399_),
    .B2(_0443_),
    .C1(_1477_),
    .Y(_1478_));
 sky130_fd_sc_hd__and4_1 _4972_ (.A(_1469_),
    .B(_1472_),
    .C(_1475_),
    .D(_1478_),
    .X(_1479_));
 sky130_fd_sc_hd__or2_1 _4973_ (.A(_0883_),
    .B(_0425_),
    .X(_1480_));
 sky130_fd_sc_hd__o21ai_1 _4974_ (.A1(_0965_),
    .A2(_0422_),
    .B1(_1480_),
    .Y(_1481_));
 sky130_fd_sc_hd__a221oi_1 _4975_ (.A1(_0461_),
    .A2(_0415_),
    .B1(_0459_),
    .B2(_0419_),
    .C1(_1481_),
    .Y(_1482_));
 sky130_fd_sc_hd__nand2_1 _4976_ (.A(_0442_),
    .B(_0447_),
    .Y(_1483_));
 sky130_fd_sc_hd__o21ai_1 _4977_ (.A1(_0647_),
    .A2(_0439_),
    .B1(_1483_),
    .Y(_1484_));
 sky130_fd_sc_hd__a221oi_1 _4978_ (.A1(_0471_),
    .A2(_0432_),
    .B1(_0435_),
    .B2(_0478_),
    .C1(_1484_),
    .Y(_1485_));
 sky130_fd_sc_hd__nand2_1 _4979_ (.A(_0453_),
    .B(_0664_),
    .Y(_1486_));
 sky130_fd_sc_hd__nand2_1 _4980_ (.A(_0458_),
    .B(_0751_),
    .Y(_1487_));
 sky130_fd_sc_hd__or2_1 _4981_ (.A(_1297_),
    .B(_0450_),
    .X(_1488_));
 sky130_fd_sc_hd__o2111a_1 _4982_ (.A1(_0663_),
    .A2(_0464_),
    .B1(_1486_),
    .C1(_1487_),
    .D1(_1488_),
    .X(_1489_));
 sky130_fd_sc_hd__nand2_1 _4983_ (.A(_0470_),
    .B(_3237_),
    .Y(_1490_));
 sky130_fd_sc_hd__o21ai_1 _4984_ (.A1(_1043_),
    .A2(_0472_),
    .B1(_1490_),
    .Y(_1491_));
 sky130_fd_sc_hd__a221oi_1 _4985_ (.A1(_3217_),
    .A2(_0477_),
    .B1(_3221_),
    .B2(_2936_),
    .C1(_1491_),
    .Y(_1492_));
 sky130_fd_sc_hd__and4_1 _4986_ (.A(_1482_),
    .B(_1485_),
    .C(_1489_),
    .D(_1492_),
    .X(_1493_));
 sky130_fd_sc_hd__nand2_1 _4987_ (.A(_1479_),
    .B(_1493_),
    .Y(_1494_));
 sky130_fd_sc_hd__a22o_1 _4988_ (.A1(\egd_top.BitStream_buffer.BS_buffer[27] ),
    .A2(_0503_),
    .B1(_0508_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[28] ),
    .X(_1495_));
 sky130_fd_sc_hd__a221oi_1 _4989_ (.A1(\egd_top.BitStream_buffer.BS_buffer[29] ),
    .A2(_0514_),
    .B1(_0537_),
    .B2(_0901_),
    .C1(_1495_),
    .Y(_1496_));
 sky130_fd_sc_hd__o22a_1 _4990_ (.A1(_0995_),
    .A2(_0530_),
    .B1(_0366_),
    .B2(_0534_),
    .X(_1497_));
 sky130_fd_sc_hd__o221a_1 _4991_ (.A1(_0907_),
    .A2(_0523_),
    .B1(_0633_),
    .B2(_0526_),
    .C1(_1497_),
    .X(_1498_));
 sky130_fd_sc_hd__nand2_1 _4992_ (.A(_0497_),
    .B(_0531_),
    .Y(_1499_));
 sky130_fd_sc_hd__o21ai_1 _4993_ (.A1(_0528_),
    .A2(_0495_),
    .B1(_1499_),
    .Y(_1500_));
 sky130_fd_sc_hd__a221oi_1 _4994_ (.A1(_0509_),
    .A2(_0487_),
    .B1(_0519_),
    .B2(_0490_),
    .C1(_1500_),
    .Y(_1501_));
 sky130_fd_sc_hd__nand2_1 _4995_ (.A(_0548_),
    .B(_0364_),
    .Y(_1502_));
 sky130_fd_sc_hd__o21ai_1 _4996_ (.A1(_0940_),
    .A2(_0546_),
    .B1(_1502_),
    .Y(_1503_));
 sky130_fd_sc_hd__a221oi_1 _4997_ (.A1(_0346_),
    .A2(_0539_),
    .B1(_0354_),
    .B2(_0542_),
    .C1(_1503_),
    .Y(_1504_));
 sky130_fd_sc_hd__and4_1 _4998_ (.A(_1496_),
    .B(_1498_),
    .C(_1501_),
    .D(_1504_),
    .X(_1505_));
 sky130_fd_sc_hd__nand2_1 _4999_ (.A(_0561_),
    .B(\egd_top.BitStream_buffer.BS_buffer[13] ),
    .Y(_1506_));
 sky130_fd_sc_hd__nand2_1 _5000_ (.A(_0565_),
    .B(\egd_top.BitStream_buffer.BS_buffer[11] ),
    .Y(_1507_));
 sky130_fd_sc_hd__or2_1 _5001_ (.A(_0676_),
    .B(_0571_),
    .X(_1508_));
 sky130_fd_sc_hd__o2111a_1 _5002_ (.A1(_0688_),
    .A2(_0558_),
    .B1(_1506_),
    .C1(_1507_),
    .D1(_1508_),
    .X(_1509_));
 sky130_fd_sc_hd__nand2_1 _5003_ (.A(_0582_),
    .B(\egd_top.BitStream_buffer.BS_buffer[17] ),
    .Y(_1510_));
 sky130_fd_sc_hd__nand2_1 _5004_ (.A(_0578_),
    .B(\egd_top.BitStream_buffer.BS_buffer[15] ),
    .Y(_1511_));
 sky130_fd_sc_hd__or2_1 _5005_ (.A(_0685_),
    .B(_0588_),
    .X(_1512_));
 sky130_fd_sc_hd__o2111a_1 _5006_ (.A1(_0492_),
    .A2(_0576_),
    .B1(_1510_),
    .C1(_1511_),
    .D1(_1512_),
    .X(_1513_));
 sky130_fd_sc_hd__or2_1 _5007_ (.A(_0670_),
    .B(_0596_),
    .X(_1514_));
 sky130_fd_sc_hd__o221a_1 _5008_ (.A1(_0586_),
    .A2(_0593_),
    .B1(_0679_),
    .B2(_0599_),
    .C1(_1514_),
    .X(_1515_));
 sky130_fd_sc_hd__nand2_1 _5009_ (.A(_0606_),
    .B(_0498_),
    .Y(_1516_));
 sky130_fd_sc_hd__nand2_1 _5010_ (.A(_0609_),
    .B(_0505_),
    .Y(_1517_));
 sky130_fd_sc_hd__or2_1 _5011_ (.A(_0897_),
    .B(_0613_),
    .X(_1518_));
 sky130_fd_sc_hd__o2111a_1 _5012_ (.A1(_1128_),
    .A2(_0604_),
    .B1(_1516_),
    .C1(_1517_),
    .D1(_1518_),
    .X(_1519_));
 sky130_fd_sc_hd__and4_1 _5013_ (.A(_1509_),
    .B(_1513_),
    .C(_1515_),
    .D(_1519_),
    .X(_1520_));
 sky130_fd_sc_hd__nand2_1 _5014_ (.A(_1505_),
    .B(_1520_),
    .Y(_1521_));
 sky130_fd_sc_hd__nor2_1 _5015_ (.A(_1494_),
    .B(_1521_),
    .Y(_1522_));
 sky130_fd_sc_hd__nand2_1 _5016_ (.A(_3061_),
    .B(_3109_),
    .Y(_1523_));
 sky130_fd_sc_hd__o21ai_1 _5017_ (.A1(_3119_),
    .A2(_3056_),
    .B1(_1523_),
    .Y(_1524_));
 sky130_fd_sc_hd__a221oi_1 _5018_ (.A1(_0714_),
    .A2(_3039_),
    .B1(_3128_),
    .B2(_3048_),
    .C1(_1524_),
    .Y(_1525_));
 sky130_fd_sc_hd__nand2_1 _5019_ (.A(_3093_),
    .B(_3118_),
    .Y(_1526_));
 sky130_fd_sc_hd__nand2_1 _5020_ (.A(_3099_),
    .B(_3070_),
    .Y(_1527_));
 sky130_fd_sc_hd__or2_1 _5021_ (.A(_1025_),
    .B(_3106_),
    .X(_1528_));
 sky130_fd_sc_hd__o2111a_1 _5022_ (.A1(_0808_),
    .A2(_3089_),
    .B1(_1526_),
    .C1(_1527_),
    .D1(_1528_),
    .X(_1529_));
 sky130_fd_sc_hd__nand2_1 _5023_ (.A(_3127_),
    .B(_3082_),
    .Y(_1530_));
 sky130_fd_sc_hd__o21ai_1 _5024_ (.A1(_2977_),
    .A2(_3123_),
    .B1(_1530_),
    .Y(_1531_));
 sky130_fd_sc_hd__a221oi_1 _5025_ (.A1(_3164_),
    .A2(_3113_),
    .B1(_3117_),
    .B2(_3153_),
    .C1(_1531_),
    .Y(_1532_));
 sky130_fd_sc_hd__nand2_1 _5026_ (.A(_3074_),
    .B(_3204_),
    .Y(_1533_));
 sky130_fd_sc_hd__o21ai_1 _5027_ (.A1(_2986_),
    .A2(_0729_),
    .B1(_1533_),
    .Y(_1534_));
 sky130_fd_sc_hd__a221oi_1 _5028_ (.A1(_0746_),
    .A2(_0726_),
    .B1(_3191_),
    .B2(_3081_),
    .C1(_1534_),
    .Y(_1535_));
 sky130_fd_sc_hd__and4_1 _5029_ (.A(_1525_),
    .B(_1529_),
    .C(_1532_),
    .D(_1535_),
    .X(_1536_));
 sky130_fd_sc_hd__nand2_1 _5030_ (.A(_3148_),
    .B(_0623_),
    .Y(_1537_));
 sky130_fd_sc_hd__o21ai_1 _5031_ (.A1(_3024_),
    .A2(_3145_),
    .B1(_1537_),
    .Y(_1538_));
 sky130_fd_sc_hd__a221oi_1 _5032_ (.A1(_0792_),
    .A2(_3137_),
    .B1(_0930_),
    .B2(_3141_),
    .C1(_1538_),
    .Y(_1539_));
 sky130_fd_sc_hd__nand2_1 _5033_ (.A(_3163_),
    .B(_0744_),
    .Y(_1540_));
 sky130_fd_sc_hd__nand2_1 _5034_ (.A(_3168_),
    .B(_3198_),
    .Y(_1541_));
 sky130_fd_sc_hd__nand2_1 _5035_ (.A(_1540_),
    .B(_1541_),
    .Y(_1542_));
 sky130_fd_sc_hd__a221oi_1 _5036_ (.A1(_3149_),
    .A2(_3156_),
    .B1(_3133_),
    .B2(_3160_),
    .C1(_1542_),
    .Y(_1543_));
 sky130_fd_sc_hd__nand2_1 _5037_ (.A(_3203_),
    .B(_3138_),
    .Y(_1544_));
 sky130_fd_sc_hd__o21ai_1 _5038_ (.A1(_3015_),
    .A2(_3200_),
    .B1(_1544_),
    .Y(_1545_));
 sky130_fd_sc_hd__a221oi_1 _5039_ (.A1(_3177_),
    .A2(_3194_),
    .B1(_3197_),
    .B2(_0741_),
    .C1(_1545_),
    .Y(_1546_));
 sky130_fd_sc_hd__nand2_1 _5040_ (.A(_3186_),
    .B(_0562_),
    .Y(_1547_));
 sky130_fd_sc_hd__o21ai_1 _5041_ (.A1(_0569_),
    .A2(_3183_),
    .B1(_1547_),
    .Y(_1548_));
 sky130_fd_sc_hd__a221oi_1 _5042_ (.A1(_1076_),
    .A2(_3176_),
    .B1(_0566_),
    .B2(_3180_),
    .C1(_1548_),
    .Y(_1549_));
 sky130_fd_sc_hd__and4_1 _5043_ (.A(_1539_),
    .B(_1543_),
    .C(_1546_),
    .D(_1549_),
    .X(_1550_));
 sky130_fd_sc_hd__nand2_1 _5044_ (.A(_1536_),
    .B(_1550_),
    .Y(_1551_));
 sky130_fd_sc_hd__nand2_1 _5045_ (.A(_3301_),
    .B(_3334_),
    .Y(_1552_));
 sky130_fd_sc_hd__o21ai_1 _5046_ (.A1(_3306_),
    .A2(_3299_),
    .B1(_1552_),
    .Y(_1553_));
 sky130_fd_sc_hd__a221oi_1 _5047_ (.A1(_0780_),
    .A2(_3292_),
    .B1(_3322_),
    .B2(_3295_),
    .C1(_1553_),
    .Y(_1554_));
 sky130_fd_sc_hd__nand2_1 _5048_ (.A(_3314_),
    .B(_3327_),
    .Y(_1555_));
 sky130_fd_sc_hd__nand2_1 _5049_ (.A(_3310_),
    .B(_0785_),
    .Y(_1556_));
 sky130_fd_sc_hd__or2_1 _5050_ (.A(_1003_),
    .B(_3319_),
    .X(_1557_));
 sky130_fd_sc_hd__o2111a_1 _5051_ (.A1(_0784_),
    .A2(_3308_),
    .B1(_1555_),
    .C1(_1556_),
    .D1(_1557_),
    .X(_1558_));
 sky130_fd_sc_hd__nand2_1 _5052_ (.A(_1554_),
    .B(_1558_),
    .Y(_1559_));
 sky130_fd_sc_hd__nand2_1 _5053_ (.A(_0323_),
    .B(_3100_),
    .Y(_1560_));
 sky130_fd_sc_hd__nand2_1 _5054_ (.A(_0329_),
    .B(_3062_),
    .Y(_1561_));
 sky130_fd_sc_hd__nand2_1 _5055_ (.A(_3340_),
    .B(_0716_),
    .Y(_1562_));
 sky130_fd_sc_hd__o2111ai_1 _5056_ (.A1(_0796_),
    .A2(_0327_),
    .B1(_1560_),
    .C1(_1561_),
    .D1(_1562_),
    .Y(_1563_));
 sky130_fd_sc_hd__inv_2 _5057_ (.A(_3329_),
    .Y(_1564_));
 sky130_fd_sc_hd__a22o_1 _5058_ (.A1(_3040_),
    .A2(_3323_),
    .B1(_3325_),
    .B2(_0708_),
    .X(_1565_));
 sky130_fd_sc_hd__a221o_1 _5059_ (.A1(_3028_),
    .A2(_1564_),
    .B1(_3341_),
    .B2(_3333_),
    .C1(_1565_),
    .X(_1566_));
 sky130_fd_sc_hd__nor3_1 _5060_ (.A(_1559_),
    .B(_1563_),
    .C(_1566_),
    .Y(_1567_));
 sky130_fd_sc_hd__nand2_1 _5061_ (.A(_3263_),
    .B(_0837_),
    .Y(_1568_));
 sky130_fd_sc_hd__o21ai_1 _5062_ (.A1(_3277_),
    .A2(_3260_),
    .B1(_1568_),
    .Y(_1569_));
 sky130_fd_sc_hd__a221oi_1 _5063_ (.A1(_3302_),
    .A2(_3251_),
    .B1(_3288_),
    .B2(_3255_),
    .C1(_1569_),
    .Y(_1570_));
 sky130_fd_sc_hd__nand2_1 _5064_ (.A(_3243_),
    .B(_3227_),
    .Y(_1571_));
 sky130_fd_sc_hd__o21ai_1 _5065_ (.A1(_3257_),
    .A2(_3240_),
    .B1(_1571_),
    .Y(_1572_));
 sky130_fd_sc_hd__a221oi_1 _5066_ (.A1(_3264_),
    .A2(_3233_),
    .B1(_3236_),
    .B2(_3248_),
    .C1(_1572_),
    .Y(_1573_));
 sky130_fd_sc_hd__inv_2 _5067_ (.A(\egd_top.BitStream_buffer.BS_buffer[78] ),
    .Y(_1574_));
 sky130_fd_sc_hd__nand2_1 _5068_ (.A(_3224_),
    .B(_3272_),
    .Y(_1575_));
 sky130_fd_sc_hd__o21ai_1 _5069_ (.A1(_1574_),
    .A2(_1145_),
    .B1(_1575_),
    .Y(_1576_));
 sky130_fd_sc_hd__a221oi_1 _5070_ (.A1(_3252_),
    .A2(_3216_),
    .B1(_3268_),
    .B2(_3220_),
    .C1(_1576_),
    .Y(_1577_));
 sky130_fd_sc_hd__nand2_1 _5071_ (.A(_3282_),
    .B(_0774_),
    .Y(_1578_));
 sky130_fd_sc_hd__o21ai_1 _5072_ (.A1(_0771_),
    .A2(_3279_),
    .B1(_1578_),
    .Y(_1579_));
 sky130_fd_sc_hd__a221oi_1 _5073_ (.A1(_3293_),
    .A2(_3271_),
    .B1(_3315_),
    .B2(_3275_),
    .C1(_1579_),
    .Y(_1580_));
 sky130_fd_sc_hd__and4_1 _5074_ (.A(_1570_),
    .B(_1573_),
    .C(_1577_),
    .D(_1580_),
    .X(_1581_));
 sky130_fd_sc_hd__nand2_1 _5075_ (.A(_1567_),
    .B(_1581_),
    .Y(_1582_));
 sky130_fd_sc_hd__nor2_1 _5076_ (.A(_1551_),
    .B(_1582_),
    .Y(_1583_));
 sky130_fd_sc_hd__nand2_1 _5077_ (.A(_0622_),
    .B(_0553_),
    .Y(_1584_));
 sky130_fd_sc_hd__nand3_1 _5078_ (.A(_1522_),
    .B(_1583_),
    .C(_1584_),
    .Y(_1585_));
 sky130_fd_sc_hd__clkinv_2 _5079_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[8] ),
    .Y(_1586_));
 sky130_fd_sc_hd__a21oi_1 _5080_ (.A1(_1586_),
    .A2(_3027_),
    .B1(_2905_),
    .Y(_1587_));
 sky130_fd_sc_hd__o21a_1 _5081_ (.A1(_3027_),
    .A2(_1585_),
    .B1(_1587_),
    .X(_0290_));
 sky130_fd_sc_hd__nand2_1 _5082_ (.A(_3061_),
    .B(_3118_),
    .Y(_1588_));
 sky130_fd_sc_hd__o21ai_1 _5083_ (.A1(_0721_),
    .A2(_3056_),
    .B1(_1588_),
    .Y(_1589_));
 sky130_fd_sc_hd__a221oi_1 _5084_ (.A1(_3128_),
    .A2(_3039_),
    .B1(_0722_),
    .B2(_3048_),
    .C1(_1589_),
    .Y(_1590_));
 sky130_fd_sc_hd__nand2_1 _5085_ (.A(_3093_),
    .B(_3066_),
    .Y(_1591_));
 sky130_fd_sc_hd__nand2_1 _5086_ (.A(_3099_),
    .B(_3075_),
    .Y(_1592_));
 sky130_fd_sc_hd__or2_1 _5087_ (.A(_0727_),
    .B(_3106_),
    .X(_1593_));
 sky130_fd_sc_hd__o2111a_1 _5088_ (.A1(_1035_),
    .A2(_3089_),
    .B1(_1591_),
    .C1(_1592_),
    .D1(_1593_),
    .X(_1594_));
 sky130_fd_sc_hd__nand2_1 _5089_ (.A(_3127_),
    .B(_3169_),
    .Y(_1595_));
 sky130_fd_sc_hd__o21ai_1 _5090_ (.A1(_2980_),
    .A2(_3123_),
    .B1(_1595_),
    .Y(_1596_));
 sky130_fd_sc_hd__a221oi_1 _5091_ (.A1(_3153_),
    .A2(_3113_),
    .B1(_3117_),
    .B2(_3157_),
    .C1(_1596_),
    .Y(_1597_));
 sky130_fd_sc_hd__nand2_1 _5092_ (.A(_3074_),
    .B(_0746_),
    .Y(_1598_));
 sky130_fd_sc_hd__o21ai_1 _5093_ (.A1(_2990_),
    .A2(_0729_),
    .B1(_1598_),
    .Y(_1599_));
 sky130_fd_sc_hd__a221oi_1 _5094_ (.A1(_3191_),
    .A2(_0726_),
    .B1(_3198_),
    .B2(_3081_),
    .C1(_1599_),
    .Y(_1600_));
 sky130_fd_sc_hd__and4_1 _5095_ (.A(_1590_),
    .B(_1594_),
    .C(_1597_),
    .D(_1600_),
    .X(_1601_));
 sky130_fd_sc_hd__inv_2 _5096_ (.A(\egd_top.BitStream_buffer.BS_buffer[0] ),
    .Y(_1602_));
 sky130_fd_sc_hd__nand2_1 _5097_ (.A(_3148_),
    .B(_0792_),
    .Y(_1603_));
 sky130_fd_sc_hd__o21ai_1 _5098_ (.A1(_1602_),
    .A2(_3145_),
    .B1(_1603_),
    .Y(_1604_));
 sky130_fd_sc_hd__a221oi_1 _5099_ (.A1(_0930_),
    .A2(_3137_),
    .B1(_1076_),
    .B2(_3141_),
    .C1(_1604_),
    .Y(_1605_));
 sky130_fd_sc_hd__nand2_1 _5100_ (.A(_3163_),
    .B(_3149_),
    .Y(_1606_));
 sky130_fd_sc_hd__nand2_1 _5101_ (.A(_3168_),
    .B(_0744_),
    .Y(_1607_));
 sky130_fd_sc_hd__nand2_1 _5102_ (.A(_1606_),
    .B(_1607_),
    .Y(_1608_));
 sky130_fd_sc_hd__a221oi_1 _5103_ (.A1(_3133_),
    .A2(_3156_),
    .B1(_3138_),
    .B2(_3160_),
    .C1(_1608_),
    .Y(_1609_));
 sky130_fd_sc_hd__nand2_1 _5104_ (.A(_3203_),
    .B(_3173_),
    .Y(_1610_));
 sky130_fd_sc_hd__o21ai_1 _5105_ (.A1(_3018_),
    .A2(_3200_),
    .B1(_1610_),
    .Y(_1611_));
 sky130_fd_sc_hd__a221oi_1 _5106_ (.A1(_0741_),
    .A2(_3194_),
    .B1(_3197_),
    .B2(_3187_),
    .C1(_1611_),
    .Y(_1612_));
 sky130_fd_sc_hd__nand2_1 _5107_ (.A(_3186_),
    .B(_0553_),
    .Y(_1613_));
 sky130_fd_sc_hd__o21ai_1 _5108_ (.A1(_0673_),
    .A2(_3183_),
    .B1(_1613_),
    .Y(_1614_));
 sky130_fd_sc_hd__a221oi_1 _5109_ (.A1(_0566_),
    .A2(_3176_),
    .B1(_0568_),
    .B2(_3180_),
    .C1(_1614_),
    .Y(_1615_));
 sky130_fd_sc_hd__and4_1 _5110_ (.A(_1605_),
    .B(_1609_),
    .C(_1612_),
    .D(_1615_),
    .X(_1616_));
 sky130_fd_sc_hd__nand2_1 _5111_ (.A(_1601_),
    .B(_1616_),
    .Y(_1617_));
 sky130_fd_sc_hd__a22o_1 _5112_ (.A1(_3288_),
    .A2(_3251_),
    .B1(_3255_),
    .B2(_3293_),
    .X(_1618_));
 sky130_fd_sc_hd__a221oi_1 _5113_ (.A1(_0837_),
    .A2(_3259_),
    .B1(_3302_),
    .B2(_3263_),
    .C1(_1618_),
    .Y(_1619_));
 sky130_fd_sc_hd__nand2_1 _5114_ (.A(_3243_),
    .B(_3256_),
    .Y(_1620_));
 sky130_fd_sc_hd__o21ai_1 _5115_ (.A1(_0759_),
    .A2(_3240_),
    .B1(_1620_),
    .Y(_1621_));
 sky130_fd_sc_hd__a221oi_1 _5116_ (.A1(_3248_),
    .A2(_3233_),
    .B1(_3236_),
    .B2(_3252_),
    .C1(_1621_),
    .Y(_1622_));
 sky130_fd_sc_hd__nand2_1 _5117_ (.A(_3224_),
    .B(_3283_),
    .Y(_1623_));
 sky130_fd_sc_hd__o21ai_1 _5118_ (.A1(_3277_),
    .A2(_1145_),
    .B1(_1623_),
    .Y(_1624_));
 sky130_fd_sc_hd__a221oi_1 _5119_ (.A1(_3268_),
    .A2(_3216_),
    .B1(_3272_),
    .B2(_3220_),
    .C1(_1624_),
    .Y(_1625_));
 sky130_fd_sc_hd__nand2_1 _5120_ (.A(_3282_),
    .B(_3311_),
    .Y(_1626_));
 sky130_fd_sc_hd__o21ai_1 _5121_ (.A1(_3306_),
    .A2(_3279_),
    .B1(_1626_),
    .Y(_1627_));
 sky130_fd_sc_hd__a221oi_1 _5122_ (.A1(_3315_),
    .A2(_3271_),
    .B1(_0774_),
    .B2(_3275_),
    .C1(_1627_),
    .Y(_1628_));
 sky130_fd_sc_hd__and4_1 _5123_ (.A(_1619_),
    .B(_1622_),
    .C(_1625_),
    .D(_1628_),
    .X(_1629_));
 sky130_fd_sc_hd__nand2_1 _5124_ (.A(_3301_),
    .B(_0780_),
    .Y(_1630_));
 sky130_fd_sc_hd__o21ai_1 _5125_ (.A1(_0776_),
    .A2(_3299_),
    .B1(_1630_),
    .Y(_1631_));
 sky130_fd_sc_hd__a221oi_1 _5126_ (.A1(_3322_),
    .A2(_3292_),
    .B1(_3327_),
    .B2(_3295_),
    .C1(_1631_),
    .Y(_1632_));
 sky130_fd_sc_hd__nand2_1 _5127_ (.A(_3314_),
    .B(_0330_),
    .Y(_1633_));
 sky130_fd_sc_hd__nand2_1 _5128_ (.A(_3310_),
    .B(_3338_),
    .Y(_1634_));
 sky130_fd_sc_hd__or2_1 _5129_ (.A(_0324_),
    .B(_3319_),
    .X(_1635_));
 sky130_fd_sc_hd__o2111a_1 _5130_ (.A1(_0854_),
    .A2(_3308_),
    .B1(_1633_),
    .C1(_1634_),
    .D1(_1635_),
    .X(_1636_));
 sky130_fd_sc_hd__nand2_1 _5131_ (.A(_3333_),
    .B(_3028_),
    .Y(_1637_));
 sky130_fd_sc_hd__o21ai_1 _5132_ (.A1(_1169_),
    .A2(_3330_),
    .B1(_1637_),
    .Y(_1638_));
 sky130_fd_sc_hd__a221oi_1 _5133_ (.A1(_0708_),
    .A2(_3324_),
    .B1(_3326_),
    .B2(_3062_),
    .C1(_1638_),
    .Y(_1639_));
 sky130_fd_sc_hd__nand2_1 _5134_ (.A(_0329_),
    .B(_3094_),
    .Y(_1640_));
 sky130_fd_sc_hd__o21ai_1 _5135_ (.A1(_3102_),
    .A2(_0327_),
    .B1(_1640_),
    .Y(_1641_));
 sky130_fd_sc_hd__a221oi_1 _5136_ (.A1(_3100_),
    .A2(_3340_),
    .B1(_0714_),
    .B2(_0323_),
    .C1(_1641_),
    .Y(_1642_));
 sky130_fd_sc_hd__and4_1 _5137_ (.A(_1632_),
    .B(_1636_),
    .C(_1639_),
    .D(_1642_),
    .X(_1643_));
 sky130_fd_sc_hd__nand2_1 _5138_ (.A(_1629_),
    .B(_1643_),
    .Y(_1644_));
 sky130_fd_sc_hd__nor2_1 _5139_ (.A(_1617_),
    .B(_1644_),
    .Y(_1645_));
 sky130_fd_sc_hd__nand2_1 _5140_ (.A(_0353_),
    .B(_0407_),
    .Y(_1646_));
 sky130_fd_sc_hd__o21ai_1 _5141_ (.A1(_0401_),
    .A2(_0350_),
    .B1(_1646_),
    .Y(_1647_));
 sky130_fd_sc_hd__a221oi_1 _5142_ (.A1(_0393_),
    .A2(_0342_),
    .B1(_0345_),
    .B2(_0400_),
    .C1(_1647_),
    .Y(_1648_));
 sky130_fd_sc_hd__nand2_1 _5143_ (.A(_0388_),
    .B(_0412_),
    .Y(_1649_));
 sky130_fd_sc_hd__o21ai_1 _5144_ (.A1(_0879_),
    .A2(_0385_),
    .B1(_1649_),
    .Y(_1650_));
 sky130_fd_sc_hd__a221oi_1 _5145_ (.A1(_0874_),
    .A2(_0378_),
    .B1(_0948_),
    .B2(_0382_),
    .C1(_1650_),
    .Y(_1651_));
 sky130_fd_sc_hd__nand2_1 _5146_ (.A(_0371_),
    .B(_0375_),
    .Y(_1652_));
 sky130_fd_sc_hd__o21ai_1 _5147_ (.A1(_0861_),
    .A2(_0368_),
    .B1(_1652_),
    .Y(_1653_));
 sky130_fd_sc_hd__a221oi_1 _5148_ (.A1(_0389_),
    .A2(_0360_),
    .B1(_0363_),
    .B2(_0869_),
    .C1(_1653_),
    .Y(_1654_));
 sky130_fd_sc_hd__nand2_1 _5149_ (.A(_0406_),
    .B(_0429_),
    .Y(_1655_));
 sky130_fd_sc_hd__o21ai_1 _5150_ (.A1(_0883_),
    .A2(_0403_),
    .B1(_1655_),
    .Y(_1656_));
 sky130_fd_sc_hd__a221oi_1 _5151_ (.A1(_0443_),
    .A2(_0396_),
    .B1(_0399_),
    .B2(_0655_),
    .C1(_1656_),
    .Y(_1657_));
 sky130_fd_sc_hd__and4_1 _5152_ (.A(_1648_),
    .B(_1651_),
    .C(_1654_),
    .D(_1657_),
    .X(_1658_));
 sky130_fd_sc_hd__or2_1 _5153_ (.A(_0965_),
    .B(_0425_),
    .X(_1659_));
 sky130_fd_sc_hd__o21ai_1 _5154_ (.A1(_0462_),
    .A2(_0422_),
    .B1(_1659_),
    .Y(_1660_));
 sky130_fd_sc_hd__a221oi_1 _5155_ (.A1(_0459_),
    .A2(_0415_),
    .B1(_0447_),
    .B2(_0419_),
    .C1(_1660_),
    .Y(_1661_));
 sky130_fd_sc_hd__nand2_1 _5156_ (.A(_0442_),
    .B(_0467_),
    .Y(_1662_));
 sky130_fd_sc_hd__o21ai_1 _5157_ (.A1(_0887_),
    .A2(_0439_),
    .B1(_1662_),
    .Y(_1663_));
 sky130_fd_sc_hd__a221oi_1 _5158_ (.A1(_0478_),
    .A2(_0432_),
    .B1(_0435_),
    .B2(_0664_),
    .C1(_1663_),
    .Y(_1664_));
 sky130_fd_sc_hd__nand2_1 _5159_ (.A(_0458_),
    .B(_3230_),
    .Y(_1665_));
 sky130_fd_sc_hd__nand2_1 _5160_ (.A(_0453_),
    .B(_3244_),
    .Y(_1666_));
 sky130_fd_sc_hd__or2_1 _5161_ (.A(_3238_),
    .B(_0464_),
    .X(_1667_));
 sky130_fd_sc_hd__o2111a_1 _5162_ (.A1(_0829_),
    .A2(_0450_),
    .B1(_1665_),
    .C1(_1666_),
    .D1(_1667_),
    .X(_1668_));
 sky130_fd_sc_hd__nand2_1 _5163_ (.A(_0470_),
    .B(_3210_),
    .Y(_1669_));
 sky130_fd_sc_hd__o21ai_1 _5164_ (.A1(_1360_),
    .A2(_0472_),
    .B1(_1669_),
    .Y(_1670_));
 sky130_fd_sc_hd__a221oi_1 _5165_ (.A1(_3221_),
    .A2(_0477_),
    .B1(_3227_),
    .B2(_2936_),
    .C1(_1670_),
    .Y(_1671_));
 sky130_fd_sc_hd__and4_1 _5166_ (.A(_1661_),
    .B(_1664_),
    .C(_1668_),
    .D(_1671_),
    .X(_1672_));
 sky130_fd_sc_hd__nand2_1 _5167_ (.A(_1658_),
    .B(_1672_),
    .Y(_1673_));
 sky130_fd_sc_hd__nand2_1 _5168_ (.A(_0497_),
    .B(\egd_top.BitStream_buffer.BS_buffer[27] ),
    .Y(_1674_));
 sky130_fd_sc_hd__o21ai_1 _5169_ (.A1(_0532_),
    .A2(_0495_),
    .B1(_1674_),
    .Y(_1675_));
 sky130_fd_sc_hd__a221oi_1 _5170_ (.A1(_0519_),
    .A2(_0487_),
    .B1(_0527_),
    .B2(_0490_),
    .C1(_1675_),
    .Y(_1676_));
 sky130_fd_sc_hd__nand2_1 _5171_ (.A(_0514_),
    .B(_0537_),
    .Y(_1677_));
 sky130_fd_sc_hd__o21ai_1 _5172_ (.A1(_0907_),
    .A2(_0512_),
    .B1(_1677_),
    .Y(_1678_));
 sky130_fd_sc_hd__a221oi_1 _5173_ (.A1(\egd_top.BitStream_buffer.BS_buffer[28] ),
    .A2(_0504_),
    .B1(\egd_top.BitStream_buffer.BS_buffer[29] ),
    .B2(_0508_),
    .C1(_1678_),
    .Y(_1679_));
 sky130_fd_sc_hd__o22a_1 _5174_ (.A1(_0366_),
    .A2(_0530_),
    .B1(_0633_),
    .B2(_0534_),
    .X(_1680_));
 sky130_fd_sc_hd__o221a_1 _5175_ (.A1(_0995_),
    .A2(_0523_),
    .B1(_0865_),
    .B2(_0526_),
    .C1(_1680_),
    .X(_1681_));
 sky130_fd_sc_hd__nand2_1 _5176_ (.A(_0548_),
    .B(_0337_),
    .Y(_1682_));
 sky130_fd_sc_hd__o21ai_1 _5177_ (.A1(_1084_),
    .A2(_0546_),
    .B1(_1682_),
    .Y(_1683_));
 sky130_fd_sc_hd__a221oi_1 _5178_ (.A1(_0354_),
    .A2(_0539_),
    .B1(_0347_),
    .B2(_0542_),
    .C1(_1683_),
    .Y(_1684_));
 sky130_fd_sc_hd__and4_1 _5179_ (.A(_1676_),
    .B(_1679_),
    .C(_1681_),
    .D(_1684_),
    .X(_1685_));
 sky130_fd_sc_hd__nand2_1 _5180_ (.A(_0565_),
    .B(\egd_top.BitStream_buffer.BS_buffer[12] ),
    .Y(_1686_));
 sky130_fd_sc_hd__nand2_1 _5181_ (.A(_0561_),
    .B(\egd_top.BitStream_buffer.BS_buffer[14] ),
    .Y(_1687_));
 sky130_fd_sc_hd__or2_1 _5182_ (.A(_0611_),
    .B(_0571_),
    .X(_1688_));
 sky130_fd_sc_hd__o2111a_1 _5183_ (.A1(_0602_),
    .A2(_0558_),
    .B1(_1686_),
    .C1(_1687_),
    .D1(_1688_),
    .X(_1689_));
 sky130_fd_sc_hd__nand2_1 _5184_ (.A(_0582_),
    .B(_0491_),
    .Y(_1690_));
 sky130_fd_sc_hd__nand2_1 _5185_ (.A(_0578_),
    .B(\egd_top.BitStream_buffer.BS_buffer[16] ),
    .Y(_1691_));
 sky130_fd_sc_hd__or2_1 _5186_ (.A(_0922_),
    .B(_0588_),
    .X(_1692_));
 sky130_fd_sc_hd__o2111a_1 _5187_ (.A1(_0692_),
    .A2(_0576_),
    .B1(_1690_),
    .C1(_1691_),
    .D1(_1692_),
    .X(_1693_));
 sky130_fd_sc_hd__or2_1 _5188_ (.A(_0586_),
    .B(_0595_),
    .X(_1694_));
 sky130_fd_sc_hd__o221a_1 _5189_ (.A1(_0679_),
    .A2(_0593_),
    .B1(_0574_),
    .B2(_0599_),
    .C1(_1694_),
    .X(_1695_));
 sky130_fd_sc_hd__nand2_1 _5190_ (.A(_0606_),
    .B(_0502_),
    .Y(_1696_));
 sky130_fd_sc_hd__nand2_1 _5191_ (.A(_0609_),
    .B(_0515_),
    .Y(_1697_));
 sky130_fd_sc_hd__or2_1 _5192_ (.A(_0986_),
    .B(_0613_),
    .X(_1698_));
 sky130_fd_sc_hd__o2111a_1 _5193_ (.A1(_0510_),
    .A2(_0604_),
    .B1(_1696_),
    .C1(_1697_),
    .D1(_1698_),
    .X(_1699_));
 sky130_fd_sc_hd__and4_1 _5194_ (.A(_1689_),
    .B(_1693_),
    .C(_1695_),
    .D(_1699_),
    .X(_1700_));
 sky130_fd_sc_hd__nand2_1 _5195_ (.A(_1685_),
    .B(_1700_),
    .Y(_1701_));
 sky130_fd_sc_hd__nor2_1 _5196_ (.A(_1673_),
    .B(_1701_),
    .Y(_1702_));
 sky130_fd_sc_hd__nand2_1 _5197_ (.A(_0622_),
    .B(_0579_),
    .Y(_1703_));
 sky130_fd_sc_hd__nand3_1 _5198_ (.A(_1645_),
    .B(_1702_),
    .C(_1703_),
    .Y(_1704_));
 sky130_fd_sc_hd__clkinv_2 _5199_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[7] ),
    .Y(_1705_));
 sky130_fd_sc_hd__a21oi_1 _5200_ (.A1(_1705_),
    .A2(_3027_),
    .B1(_2905_),
    .Y(_1706_));
 sky130_fd_sc_hd__o21a_1 _5201_ (.A1(_3027_),
    .A2(_1704_),
    .B1(_1706_),
    .X(_0289_));
 sky130_fd_sc_hd__o21ai_1 _5202_ (.A1(\egd_top.BitStream_buffer.BitStream_buffer_output[6] ),
    .A2(_2965_),
    .B1(_0627_),
    .Y(_1707_));
 sky130_fd_sc_hd__a22o_1 _5203_ (.A1(\egd_top.BitStream_buffer.BS_buffer[119] ),
    .A2(_3078_),
    .B1(_3080_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[120] ),
    .X(_1708_));
 sky130_fd_sc_hd__a221oi_1 _5204_ (.A1(_0746_),
    .A2(_3069_),
    .B1(_3191_),
    .B2(_3074_),
    .C1(_1708_),
    .Y(_1709_));
 sky130_fd_sc_hd__nand2_1 _5205_ (.A(_3127_),
    .B(_3164_),
    .Y(_1710_));
 sky130_fd_sc_hd__o21ai_1 _5206_ (.A1(_2983_),
    .A2(_3123_),
    .B1(_1710_),
    .Y(_1711_));
 sky130_fd_sc_hd__a221oi_1 _5207_ (.A1(_3157_),
    .A2(_3113_),
    .B1(_3117_),
    .B2(_3204_),
    .C1(_1711_),
    .Y(_1712_));
 sky130_fd_sc_hd__nand2_1 _5208_ (.A(_3038_),
    .B(_0722_),
    .Y(_1713_));
 sky130_fd_sc_hd__nand2_1 _5209_ (.A(_3060_),
    .B(_3066_),
    .Y(_1714_));
 sky130_fd_sc_hd__nand2_1 _5210_ (.A(_3047_),
    .B(_3109_),
    .Y(_1715_));
 sky130_fd_sc_hd__o2111a_1 _5211_ (.A1(_0804_),
    .A2(_3055_),
    .B1(_1713_),
    .C1(_1714_),
    .D1(_1715_),
    .X(_1716_));
 sky130_fd_sc_hd__nand2_1 _5212_ (.A(_3098_),
    .B(_3082_),
    .Y(_1717_));
 sky130_fd_sc_hd__nand2_1 _5213_ (.A(_3092_),
    .B(_3070_),
    .Y(_1718_));
 sky130_fd_sc_hd__or2_1 _5214_ (.A(_0808_),
    .B(_3105_),
    .X(_1719_));
 sky130_fd_sc_hd__o2111a_1 _5215_ (.A1(_2977_),
    .A2(_3089_),
    .B1(_1717_),
    .C1(_1718_),
    .D1(_1719_),
    .X(_1720_));
 sky130_fd_sc_hd__and4_1 _5216_ (.A(_1709_),
    .B(_1712_),
    .C(_1716_),
    .D(_1720_),
    .X(_1721_));
 sky130_fd_sc_hd__nand2_1 _5217_ (.A(_3291_),
    .B(_3327_),
    .Y(_1722_));
 sky130_fd_sc_hd__nand2_1 _5218_ (.A(_3300_),
    .B(_3322_),
    .Y(_1723_));
 sky130_fd_sc_hd__nand2_1 _5219_ (.A(_3295_),
    .B(_0330_),
    .Y(_1724_));
 sky130_fd_sc_hd__o2111a_1 _5220_ (.A1(_3328_),
    .A2(_3298_),
    .B1(_1722_),
    .C1(_1723_),
    .D1(_1724_),
    .X(_1725_));
 sky130_fd_sc_hd__nand2_1 _5221_ (.A(_3309_),
    .B(_3341_),
    .Y(_1726_));
 sky130_fd_sc_hd__nand2_1 _5222_ (.A(_3313_),
    .B(_0785_),
    .Y(_1727_));
 sky130_fd_sc_hd__or2_1 _5223_ (.A(_1016_),
    .B(_3307_),
    .X(_1728_));
 sky130_fd_sc_hd__o2111a_1 _5224_ (.A1(_0784_),
    .A2(_3319_),
    .B1(_1726_),
    .C1(_1727_),
    .D1(_1728_),
    .X(_1729_));
 sky130_fd_sc_hd__nand2_1 _5225_ (.A(_3332_),
    .B(_3040_),
    .Y(_1730_));
 sky130_fd_sc_hd__nand2_1 _5226_ (.A(_3323_),
    .B(_3062_),
    .Y(_1731_));
 sky130_fd_sc_hd__nand2_1 _5227_ (.A(_3325_),
    .B(_3094_),
    .Y(_1732_));
 sky130_fd_sc_hd__o2111a_1 _5228_ (.A1(_3049_),
    .A2(_3329_),
    .B1(_1730_),
    .C1(_1731_),
    .D1(_1732_),
    .X(_1733_));
 sky130_fd_sc_hd__nand2_1 _5229_ (.A(_0328_),
    .B(_0716_),
    .Y(_1734_));
 sky130_fd_sc_hd__o21ai_1 _5230_ (.A1(_0713_),
    .A2(_0326_),
    .B1(_1734_),
    .Y(_1735_));
 sky130_fd_sc_hd__a221oi_1 _5231_ (.A1(_0714_),
    .A2(_3339_),
    .B1(_3128_),
    .B2(_0322_),
    .C1(_1735_),
    .Y(_1736_));
 sky130_fd_sc_hd__and4_1 _5232_ (.A(_1725_),
    .B(_1729_),
    .C(_1733_),
    .D(_1736_),
    .X(_1737_));
 sky130_fd_sc_hd__nand2_1 _5233_ (.A(_3251_),
    .B(_3293_),
    .Y(_1738_));
 sky130_fd_sc_hd__nand2_1 _5234_ (.A(_3254_),
    .B(\egd_top.BitStream_buffer.BS_buffer[84] ),
    .Y(_1739_));
 sky130_fd_sc_hd__nand2_1 _5235_ (.A(_3263_),
    .B(_3288_),
    .Y(_1740_));
 sky130_fd_sc_hd__o2111a_1 _5236_ (.A1(_0767_),
    .A2(_3260_),
    .B1(_1738_),
    .C1(_1739_),
    .D1(_1740_),
    .X(_1741_));
 sky130_fd_sc_hd__nand2_1 _5237_ (.A(_3232_),
    .B(_3252_),
    .Y(_1742_));
 sky130_fd_sc_hd__nand2_1 _5238_ (.A(_3243_),
    .B(_3264_),
    .Y(_1743_));
 sky130_fd_sc_hd__nand2_1 _5239_ (.A(_3235_),
    .B(_3268_),
    .Y(_1744_));
 sky130_fd_sc_hd__o2111a_1 _5240_ (.A1(_0833_),
    .A2(_3240_),
    .B1(_1742_),
    .C1(_1743_),
    .D1(_1744_),
    .X(_1745_));
 sky130_fd_sc_hd__nand2_1 _5241_ (.A(_3215_),
    .B(_3272_),
    .Y(_1746_));
 sky130_fd_sc_hd__nand2_1 _5242_ (.A(_3223_),
    .B(_3276_),
    .Y(_1747_));
 sky130_fd_sc_hd__nand2_1 _5243_ (.A(_3219_),
    .B(_3283_),
    .Y(_1748_));
 sky130_fd_sc_hd__o2111a_1 _5244_ (.A1(_3296_),
    .A2(_1145_),
    .B1(_1746_),
    .C1(_1747_),
    .D1(_1748_),
    .X(_1749_));
 sky130_fd_sc_hd__nand2_1 _5245_ (.A(_3270_),
    .B(_0774_),
    .Y(_1750_));
 sky130_fd_sc_hd__o21ai_1 _5246_ (.A1(_0771_),
    .A2(_3273_),
    .B1(_1750_),
    .Y(_1751_));
 sky130_fd_sc_hd__a221oi_1 _5247_ (.A1(_0772_),
    .A2(_3282_),
    .B1(_3334_),
    .B2(_1153_),
    .C1(_1751_),
    .Y(_1752_));
 sky130_fd_sc_hd__and4_1 _5248_ (.A(_1741_),
    .B(_1745_),
    .C(_1749_),
    .D(_1752_),
    .X(_1753_));
 sky130_fd_sc_hd__a22o_1 _5249_ (.A1(_0792_),
    .A2(_3144_),
    .B1(_3148_),
    .B2(_0930_),
    .X(_1754_));
 sky130_fd_sc_hd__a22o_1 _5250_ (.A1(_1076_),
    .A2(_3137_),
    .B1(_3141_),
    .B2(_0566_),
    .X(_1755_));
 sky130_fd_sc_hd__and3_1 _5251_ (.A(_3067_),
    .B(_0568_),
    .C(_3142_),
    .X(_1756_));
 sky130_fd_sc_hd__nand2_1 _5252_ (.A(_3185_),
    .B(_0579_),
    .Y(_1757_));
 sky130_fd_sc_hd__o21ai_1 _5253_ (.A1(_0554_),
    .A2(_3182_),
    .B1(_1757_),
    .Y(_1758_));
 sky130_fd_sc_hd__a211o_1 _5254_ (.A1(_0562_),
    .A2(_3179_),
    .B1(_1756_),
    .C1(_1758_),
    .X(_1759_));
 sky130_fd_sc_hd__nor3_1 _5255_ (.A(_1754_),
    .B(_1755_),
    .C(_1759_),
    .Y(_1760_));
 sky130_fd_sc_hd__nand2_1 _5256_ (.A(_3162_),
    .B(_3133_),
    .Y(_1761_));
 sky130_fd_sc_hd__nand2_1 _5257_ (.A(_3167_),
    .B(_3149_),
    .Y(_1762_));
 sky130_fd_sc_hd__nand2_1 _5258_ (.A(_1761_),
    .B(_1762_),
    .Y(_1763_));
 sky130_fd_sc_hd__a221oi_1 _5259_ (.A1(_3138_),
    .A2(_3155_),
    .B1(_3173_),
    .B2(_3159_),
    .C1(_1763_),
    .Y(_1764_));
 sky130_fd_sc_hd__nand2_1 _5260_ (.A(_3202_),
    .B(_3177_),
    .Y(_1765_));
 sky130_fd_sc_hd__o21ai_1 _5261_ (.A1(_3021_),
    .A2(_3199_),
    .B1(_1765_),
    .Y(_1766_));
 sky130_fd_sc_hd__a221oi_1 _5262_ (.A1(_3187_),
    .A2(_3193_),
    .B1(_3196_),
    .B2(_0623_),
    .C1(_1766_),
    .Y(_1767_));
 sky130_fd_sc_hd__and3_1 _5263_ (.A(_1760_),
    .B(_1764_),
    .C(_1767_),
    .X(_1768_));
 sky130_fd_sc_hd__and4_1 _5264_ (.A(_1721_),
    .B(_1737_),
    .C(_1753_),
    .D(_1768_),
    .X(_1769_));
 sky130_fd_sc_hd__or2_1 _5265_ (.A(_0462_),
    .B(_0425_),
    .X(_1770_));
 sky130_fd_sc_hd__o21ai_1 _5266_ (.A1(_0650_),
    .A2(_0422_),
    .B1(_1770_),
    .Y(_1771_));
 sky130_fd_sc_hd__a221oi_1 _5267_ (.A1(_0447_),
    .A2(_0415_),
    .B1(_0467_),
    .B2(_0419_),
    .C1(_1771_),
    .Y(_1772_));
 sky130_fd_sc_hd__nand2_1 _5268_ (.A(_0442_),
    .B(_0471_),
    .Y(_1773_));
 sky130_fd_sc_hd__o21ai_1 _5269_ (.A1(_0955_),
    .A2(_0439_),
    .B1(_1773_),
    .Y(_1774_));
 sky130_fd_sc_hd__a221oi_1 _5270_ (.A1(_0664_),
    .A2(_0432_),
    .B1(_0435_),
    .B2(_3244_),
    .C1(_1774_),
    .Y(_1775_));
 sky130_fd_sc_hd__nand2_1 _5271_ (.A(_0458_),
    .B(_3237_),
    .Y(_1776_));
 sky130_fd_sc_hd__nand2_1 _5272_ (.A(_0453_),
    .B(_0751_),
    .Y(_1777_));
 sky130_fd_sc_hd__or2_1 _5273_ (.A(_1043_),
    .B(_0449_),
    .X(_1778_));
 sky130_fd_sc_hd__o2111a_1 _5274_ (.A1(_1297_),
    .A2(_0464_),
    .B1(_1776_),
    .C1(_1777_),
    .D1(_1778_),
    .X(_1779_));
 sky130_fd_sc_hd__nand2_1 _5275_ (.A(_0477_),
    .B(_3227_),
    .Y(_1780_));
 sky130_fd_sc_hd__o21ai_1 _5276_ (.A1(_3257_),
    .A2(_2935_),
    .B1(_1780_),
    .Y(_1781_));
 sky130_fd_sc_hd__a221oi_1 _5277_ (.A1(_3217_),
    .A2(_0470_),
    .B1(_3221_),
    .B2(_0473_),
    .C1(_1781_),
    .Y(_1782_));
 sky130_fd_sc_hd__and4_1 _5278_ (.A(_1772_),
    .B(_1775_),
    .C(_1779_),
    .D(_1782_),
    .X(_1783_));
 sky130_fd_sc_hd__nand2_1 _5279_ (.A(_0371_),
    .B(_0379_),
    .Y(_1784_));
 sky130_fd_sc_hd__o21ai_1 _5280_ (.A1(_0936_),
    .A2(_0368_),
    .B1(_1784_),
    .Y(_1785_));
 sky130_fd_sc_hd__a221oi_1 _5281_ (.A1(_0869_),
    .A2(_0360_),
    .B1(_0363_),
    .B2(_0393_),
    .C1(_1785_),
    .Y(_1786_));
 sky130_fd_sc_hd__nand2_1 _5282_ (.A(_0388_),
    .B(_0416_),
    .Y(_1787_));
 sky130_fd_sc_hd__o21ai_1 _5283_ (.A1(_0960_),
    .A2(_0385_),
    .B1(_1787_),
    .Y(_1788_));
 sky130_fd_sc_hd__a221oi_1 _5284_ (.A1(_0948_),
    .A2(_0378_),
    .B1(_0412_),
    .B2(_0382_),
    .C1(_1788_),
    .Y(_1789_));
 sky130_fd_sc_hd__a22o_1 _5285_ (.A1(_0400_),
    .A2(_0341_),
    .B1(_0344_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[46] ),
    .X(_1790_));
 sky130_fd_sc_hd__a32o_1 _5286_ (.A1(_3087_),
    .A2(_0874_),
    .A3(_0339_),
    .B1(_0642_),
    .B2(_0352_),
    .X(_1791_));
 sky130_fd_sc_hd__nor2_1 _5287_ (.A(_1790_),
    .B(_1791_),
    .Y(_1792_));
 sky130_fd_sc_hd__nand2_1 _5288_ (.A(_0406_),
    .B(_0436_),
    .Y(_1793_));
 sky130_fd_sc_hd__o21ai_1 _5289_ (.A1(_0965_),
    .A2(_0403_),
    .B1(_1793_),
    .Y(_1794_));
 sky130_fd_sc_hd__a221oi_1 _5290_ (.A1(_0655_),
    .A2(_0396_),
    .B1(_0399_),
    .B2(_0429_),
    .C1(_1794_),
    .Y(_1795_));
 sky130_fd_sc_hd__and4_1 _5291_ (.A(_1786_),
    .B(_1789_),
    .C(_1792_),
    .D(_1795_),
    .X(_1796_));
 sky130_fd_sc_hd__nand2_1 _5292_ (.A(_1783_),
    .B(_1796_),
    .Y(_1797_));
 sky130_fd_sc_hd__nand2_1 _5293_ (.A(_0497_),
    .B(\egd_top.BitStream_buffer.BS_buffer[28] ),
    .Y(_1798_));
 sky130_fd_sc_hd__o21ai_1 _5294_ (.A1(_0524_),
    .A2(_0495_),
    .B1(_1798_),
    .Y(_1799_));
 sky130_fd_sc_hd__a221oi_1 _5295_ (.A1(_0527_),
    .A2(_0487_),
    .B1(_0531_),
    .B2(_0490_),
    .C1(_1799_),
    .Y(_1800_));
 sky130_fd_sc_hd__nand2_1 _5296_ (.A(_0514_),
    .B(_0540_),
    .Y(_1801_));
 sky130_fd_sc_hd__o21ai_1 _5297_ (.A1(_0995_),
    .A2(_0512_),
    .B1(_1801_),
    .Y(_1802_));
 sky130_fd_sc_hd__a221oi_1 _5298_ (.A1(\egd_top.BitStream_buffer.BS_buffer[29] ),
    .A2(_0504_),
    .B1(_0537_),
    .B2(_0508_),
    .C1(_1802_),
    .Y(_1803_));
 sky130_fd_sc_hd__o22a_1 _5299_ (.A1(_0633_),
    .A2(_0530_),
    .B1(_0865_),
    .B2(_0534_),
    .X(_1804_));
 sky130_fd_sc_hd__o221a_1 _5300_ (.A1(_0366_),
    .A2(_0523_),
    .B1(_0940_),
    .B2(_0526_),
    .C1(_1804_),
    .X(_1805_));
 sky130_fd_sc_hd__nand2_1 _5301_ (.A(_0548_),
    .B(_0346_),
    .Y(_1806_));
 sky130_fd_sc_hd__o21ai_1 _5302_ (.A1(_1276_),
    .A2(_0546_),
    .B1(_1806_),
    .Y(_1807_));
 sky130_fd_sc_hd__a221oi_1 _5303_ (.A1(_0347_),
    .A2(_0539_),
    .B1(_0375_),
    .B2(_0542_),
    .C1(_1807_),
    .Y(_1808_));
 sky130_fd_sc_hd__and4_1 _5304_ (.A(_1800_),
    .B(_1803_),
    .C(_1805_),
    .D(_1808_),
    .X(_1809_));
 sky130_fd_sc_hd__nand2_1 _5305_ (.A(_0561_),
    .B(\egd_top.BitStream_buffer.BS_buffer[15] ),
    .Y(_1810_));
 sky130_fd_sc_hd__nand2_1 _5306_ (.A(_0565_),
    .B(\egd_top.BitStream_buffer.BS_buffer[13] ),
    .Y(_1811_));
 sky130_fd_sc_hd__or2_1 _5307_ (.A(_0688_),
    .B(_0571_),
    .X(_1812_));
 sky130_fd_sc_hd__o2111a_1 _5308_ (.A1(_0685_),
    .A2(_0558_),
    .B1(_1810_),
    .C1(_1811_),
    .D1(_1812_),
    .X(_1813_));
 sky130_fd_sc_hd__nand2_1 _5309_ (.A(_0578_),
    .B(\egd_top.BitStream_buffer.BS_buffer[17] ),
    .Y(_1814_));
 sky130_fd_sc_hd__nand2_1 _5310_ (.A(_0582_),
    .B(_0498_),
    .Y(_1815_));
 sky130_fd_sc_hd__or2_1 _5311_ (.A(_0492_),
    .B(_0588_),
    .X(_1816_));
 sky130_fd_sc_hd__o2111a_1 _5312_ (.A1(_0897_),
    .A2(_0576_),
    .B1(_1814_),
    .C1(_1815_),
    .D1(_1816_),
    .X(_1817_));
 sky130_fd_sc_hd__or2_1 _5313_ (.A(_0676_),
    .B(_0599_),
    .X(_1818_));
 sky130_fd_sc_hd__o221a_1 _5314_ (.A1(_0574_),
    .A2(_0593_),
    .B1(_0679_),
    .B2(_0596_),
    .C1(_1818_),
    .X(_1819_));
 sky130_fd_sc_hd__nand2_1 _5315_ (.A(_0609_),
    .B(_0509_),
    .Y(_1820_));
 sky130_fd_sc_hd__nand2_1 _5316_ (.A(_0606_),
    .B(_0505_),
    .Y(_1821_));
 sky130_fd_sc_hd__or2_1 _5317_ (.A(_1128_),
    .B(_0613_),
    .X(_1822_));
 sky130_fd_sc_hd__o2111a_1 _5318_ (.A1(_0520_),
    .A2(_0604_),
    .B1(_1820_),
    .C1(_1821_),
    .D1(_1822_),
    .X(_1823_));
 sky130_fd_sc_hd__and4_1 _5319_ (.A(_1813_),
    .B(_1817_),
    .C(_1819_),
    .D(_1823_),
    .X(_1824_));
 sky130_fd_sc_hd__nand2_1 _5320_ (.A(_1809_),
    .B(_1824_),
    .Y(_1825_));
 sky130_fd_sc_hd__nor2_1 _5321_ (.A(_1797_),
    .B(_1825_),
    .Y(_1826_));
 sky130_fd_sc_hd__nand2_1 _5322_ (.A(_0621_),
    .B(_0585_),
    .Y(_1827_));
 sky130_fd_sc_hd__nand3_1 _5323_ (.A(_1769_),
    .B(_1826_),
    .C(_1827_),
    .Y(_1828_));
 sky130_fd_sc_hd__nor2_1 _5324_ (.A(_3026_),
    .B(_1828_),
    .Y(_1829_));
 sky130_fd_sc_hd__nor2_1 _5325_ (.A(_1707_),
    .B(_1829_),
    .Y(_0288_));
 sky130_fd_sc_hd__nand2_1 _5326_ (.A(_0371_),
    .B(_0389_),
    .Y(_1830_));
 sky130_fd_sc_hd__o21ai_1 _5327_ (.A1(_0383_),
    .A2(_0368_),
    .B1(_1830_),
    .Y(_1831_));
 sky130_fd_sc_hd__a221oi_1 _5328_ (.A1(_0393_),
    .A2(_0360_),
    .B1(_0363_),
    .B2(_0400_),
    .C1(_1831_),
    .Y(_1832_));
 sky130_fd_sc_hd__nand2_1 _5329_ (.A(_0353_),
    .B(_0874_),
    .Y(_1833_));
 sky130_fd_sc_hd__o21ai_1 _5330_ (.A1(_0420_),
    .A2(_0350_),
    .B1(_1833_),
    .Y(_1834_));
 sky130_fd_sc_hd__a221oi_1 _5331_ (.A1(_0407_),
    .A2(_0342_),
    .B1(_0345_),
    .B2(_0642_),
    .C1(_1834_),
    .Y(_1835_));
 sky130_fd_sc_hd__nand2_1 _5332_ (.A(_0378_),
    .B(_0412_),
    .Y(_1836_));
 sky130_fd_sc_hd__o21ai_1 _5333_ (.A1(_0879_),
    .A2(_0380_),
    .B1(_1836_),
    .Y(_1837_));
 sky130_fd_sc_hd__a221oi_1 _5334_ (.A1(_0443_),
    .A2(_0388_),
    .B1(_0655_),
    .B2(_0944_),
    .C1(_1837_),
    .Y(_1838_));
 sky130_fd_sc_hd__nor2_1 _5335_ (.A(_0462_),
    .B(_0403_),
    .Y(_1839_));
 sky130_fd_sc_hd__a22o_1 _5336_ (.A1(_0429_),
    .A2(_0395_),
    .B1(_0398_),
    .B2(_0436_),
    .X(_1840_));
 sky130_fd_sc_hd__a211oi_1 _5337_ (.A1(_0454_),
    .A2(_0406_),
    .B1(_1839_),
    .C1(_1840_),
    .Y(_1841_));
 sky130_fd_sc_hd__and4_1 _5338_ (.A(_1832_),
    .B(_1835_),
    .C(_1838_),
    .D(_1841_),
    .X(_1842_));
 sky130_fd_sc_hd__or2_1 _5339_ (.A(_0650_),
    .B(_0425_),
    .X(_1843_));
 sky130_fd_sc_hd__o21ai_1 _5340_ (.A1(_0448_),
    .A2(_0422_),
    .B1(_1843_),
    .Y(_1844_));
 sky130_fd_sc_hd__a221oi_1 _5341_ (.A1(_0467_),
    .A2(_0415_),
    .B1(_0471_),
    .B2(_0419_),
    .C1(_1844_),
    .Y(_1845_));
 sky130_fd_sc_hd__nand2_1 _5342_ (.A(_0442_),
    .B(_0478_),
    .Y(_1846_));
 sky130_fd_sc_hd__o21ai_1 _5343_ (.A1(_0474_),
    .A2(_0439_),
    .B1(_1846_),
    .Y(_1847_));
 sky130_fd_sc_hd__a221oi_1 _5344_ (.A1(_3244_),
    .A2(_0432_),
    .B1(_0435_),
    .B2(_0751_),
    .C1(_1847_),
    .Y(_1848_));
 sky130_fd_sc_hd__nand2_1 _5345_ (.A(_0453_),
    .B(_3230_),
    .Y(_1849_));
 sky130_fd_sc_hd__nand2_1 _5346_ (.A(_0458_),
    .B(_3210_),
    .Y(_1850_));
 sky130_fd_sc_hd__or2_1 _5347_ (.A(_0829_),
    .B(_0464_),
    .X(_1851_));
 sky130_fd_sc_hd__o2111a_1 _5348_ (.A1(_1360_),
    .A2(_0450_),
    .B1(_1849_),
    .C1(_1850_),
    .D1(_1851_),
    .X(_1852_));
 sky130_fd_sc_hd__nand2_1 _5349_ (.A(_0477_),
    .B(_3256_),
    .Y(_1853_));
 sky130_fd_sc_hd__o21ai_1 _5350_ (.A1(_0759_),
    .A2(_2935_),
    .B1(_1853_),
    .Y(_1854_));
 sky130_fd_sc_hd__a221oi_1 _5351_ (.A1(_3221_),
    .A2(_0470_),
    .B1(_3227_),
    .B2(_0473_),
    .C1(_1854_),
    .Y(_1855_));
 sky130_fd_sc_hd__and4_1 _5352_ (.A(_1845_),
    .B(_1848_),
    .C(_1852_),
    .D(_1855_),
    .X(_1856_));
 sky130_fd_sc_hd__nand2_1 _5353_ (.A(_1842_),
    .B(_1856_),
    .Y(_1857_));
 sky130_fd_sc_hd__a22o_1 _5354_ (.A1(\egd_top.BitStream_buffer.BS_buffer[32] ),
    .A2(_0514_),
    .B1(_0901_),
    .B2(_0365_),
    .X(_1858_));
 sky130_fd_sc_hd__a221oi_1 _5355_ (.A1(_0537_),
    .A2(_0504_),
    .B1(_0540_),
    .B2(_0508_),
    .C1(_1858_),
    .Y(_1859_));
 sky130_fd_sc_hd__o22a_1 _5356_ (.A1(_0865_),
    .A2(_0530_),
    .B1(_0940_),
    .B2(_0534_),
    .X(_1860_));
 sky130_fd_sc_hd__o221a_1 _5357_ (.A1(_0633_),
    .A2(_0523_),
    .B1(_1084_),
    .B2(_0526_),
    .C1(_1860_),
    .X(_1861_));
 sky130_fd_sc_hd__nand2_1 _5358_ (.A(_0497_),
    .B(\egd_top.BitStream_buffer.BS_buffer[29] ),
    .Y(_1862_));
 sky130_fd_sc_hd__o21ai_1 _5359_ (.A1(_0699_),
    .A2(_0495_),
    .B1(_1862_),
    .Y(_1863_));
 sky130_fd_sc_hd__a221oi_1 _5360_ (.A1(_0531_),
    .A2(_0487_),
    .B1(\egd_top.BitStream_buffer.BS_buffer[27] ),
    .B2(_0490_),
    .C1(_1863_),
    .Y(_1864_));
 sky130_fd_sc_hd__nand2_1 _5361_ (.A(_0548_),
    .B(_0354_),
    .Y(_1865_));
 sky130_fd_sc_hd__o21ai_1 _5362_ (.A1(_0348_),
    .A2(_0546_),
    .B1(_1865_),
    .Y(_1866_));
 sky130_fd_sc_hd__a221oi_1 _5363_ (.A1(_0375_),
    .A2(_0539_),
    .B1(_0379_),
    .B2(_0542_),
    .C1(_1866_),
    .Y(_1867_));
 sky130_fd_sc_hd__and4_1 _5364_ (.A(_1859_),
    .B(_1861_),
    .C(_1864_),
    .D(_1867_),
    .X(_1868_));
 sky130_fd_sc_hd__nand2_1 _5365_ (.A(_0565_),
    .B(\egd_top.BitStream_buffer.BS_buffer[14] ),
    .Y(_1869_));
 sky130_fd_sc_hd__nand2_1 _5366_ (.A(_0561_),
    .B(\egd_top.BitStream_buffer.BS_buffer[16] ),
    .Y(_1870_));
 sky130_fd_sc_hd__or2_1 _5367_ (.A(_0602_),
    .B(_0571_),
    .X(_1871_));
 sky130_fd_sc_hd__o2111a_1 _5368_ (.A1(_0922_),
    .A2(_0558_),
    .B1(_1869_),
    .C1(_1870_),
    .D1(_1871_),
    .X(_1872_));
 sky130_fd_sc_hd__nand2_1 _5369_ (.A(_0578_),
    .B(_0491_),
    .Y(_1873_));
 sky130_fd_sc_hd__nand2_1 _5370_ (.A(_0582_),
    .B(_0502_),
    .Y(_1874_));
 sky130_fd_sc_hd__or2_1 _5371_ (.A(_0692_),
    .B(_0588_),
    .X(_1875_));
 sky130_fd_sc_hd__o2111a_1 _5372_ (.A1(_0986_),
    .A2(_0576_),
    .B1(_1873_),
    .C1(_1874_),
    .D1(_1875_),
    .X(_1876_));
 sky130_fd_sc_hd__or2_1 _5373_ (.A(_0574_),
    .B(_0596_),
    .X(_1877_));
 sky130_fd_sc_hd__o221a_1 _5374_ (.A1(_0676_),
    .A2(_0593_),
    .B1(_0611_),
    .B2(_0599_),
    .C1(_1877_),
    .X(_1878_));
 sky130_fd_sc_hd__nand2_1 _5375_ (.A(_0609_),
    .B(_0519_),
    .Y(_1879_));
 sky130_fd_sc_hd__nand2_1 _5376_ (.A(_0606_),
    .B(_0515_),
    .Y(_1880_));
 sky130_fd_sc_hd__or2_1 _5377_ (.A(_0510_),
    .B(_0613_),
    .X(_1881_));
 sky130_fd_sc_hd__o2111a_1 _5378_ (.A1(_0528_),
    .A2(_0604_),
    .B1(_1879_),
    .C1(_1880_),
    .D1(_1881_),
    .X(_1882_));
 sky130_fd_sc_hd__and4_1 _5379_ (.A(_1872_),
    .B(_1876_),
    .C(_1878_),
    .D(_1882_),
    .X(_1883_));
 sky130_fd_sc_hd__nand2_1 _5380_ (.A(_1868_),
    .B(_1883_),
    .Y(_1884_));
 sky130_fd_sc_hd__nor2_1 _5381_ (.A(_1857_),
    .B(_1884_),
    .Y(_1885_));
 sky130_fd_sc_hd__nor2_1 _5382_ (.A(_0709_),
    .B(_3330_),
    .Y(_1886_));
 sky130_fd_sc_hd__a22o_1 _5383_ (.A1(_3094_),
    .A2(_3323_),
    .B1(_3325_),
    .B2(_0716_),
    .X(_1887_));
 sky130_fd_sc_hd__a211oi_1 _5384_ (.A1(_0708_),
    .A2(_3333_),
    .B1(_1886_),
    .C1(_1887_),
    .Y(_1888_));
 sky130_fd_sc_hd__nand2_1 _5385_ (.A(_3301_),
    .B(_3327_),
    .Y(_1889_));
 sky130_fd_sc_hd__o21ai_1 _5386_ (.A1(_0779_),
    .A2(_3299_),
    .B1(_1889_),
    .Y(_1890_));
 sky130_fd_sc_hd__a221oi_1 _5387_ (.A1(_0330_),
    .A2(_3292_),
    .B1(_0785_),
    .B2(_3295_),
    .C1(_1890_),
    .Y(_1891_));
 sky130_fd_sc_hd__nand2_1 _5388_ (.A(_3314_),
    .B(_3338_),
    .Y(_1892_));
 sky130_fd_sc_hd__nand2_1 _5389_ (.A(_3310_),
    .B(_3028_),
    .Y(_1893_));
 sky130_fd_sc_hd__or2_1 _5390_ (.A(_0854_),
    .B(_3319_),
    .X(_1894_));
 sky130_fd_sc_hd__o2111a_1 _5391_ (.A1(_1169_),
    .A2(_3308_),
    .B1(_1892_),
    .C1(_1893_),
    .D1(_1894_),
    .X(_1895_));
 sky130_fd_sc_hd__nand2_1 _5392_ (.A(_0329_),
    .B(_3100_),
    .Y(_1896_));
 sky130_fd_sc_hd__o21ai_1 _5393_ (.A1(_3085_),
    .A2(_0327_),
    .B1(_1896_),
    .Y(_1897_));
 sky130_fd_sc_hd__a221oi_1 _5394_ (.A1(_3128_),
    .A2(_3340_),
    .B1(_0722_),
    .B2(_0323_),
    .C1(_1897_),
    .Y(_1898_));
 sky130_fd_sc_hd__and4_1 _5395_ (.A(_1888_),
    .B(_1891_),
    .C(_1895_),
    .D(_1898_),
    .X(_1899_));
 sky130_fd_sc_hd__nand2_1 _5396_ (.A(_3263_),
    .B(_3293_),
    .Y(_1900_));
 sky130_fd_sc_hd__o21ai_1 _5397_ (.A1(_0842_),
    .A2(_3260_),
    .B1(_1900_),
    .Y(_1901_));
 sky130_fd_sc_hd__a221oi_1 _5398_ (.A1(_3315_),
    .A2(_3251_),
    .B1(_0774_),
    .B2(_3255_),
    .C1(_1901_),
    .Y(_1902_));
 sky130_fd_sc_hd__nand2_1 _5399_ (.A(_3243_),
    .B(_3248_),
    .Y(_1903_));
 sky130_fd_sc_hd__o21ai_1 _5400_ (.A1(_1144_),
    .A2(_3240_),
    .B1(_1903_),
    .Y(_1904_));
 sky130_fd_sc_hd__a221oi_1 _5401_ (.A1(_3268_),
    .A2(_3233_),
    .B1(_3236_),
    .B2(_3272_),
    .C1(_1904_),
    .Y(_1905_));
 sky130_fd_sc_hd__nand2_1 _5402_ (.A(_3224_),
    .B(_0837_),
    .Y(_1906_));
 sky130_fd_sc_hd__o21ai_1 _5403_ (.A1(_0767_),
    .A2(_1145_),
    .B1(_1906_),
    .Y(_1907_));
 sky130_fd_sc_hd__a221oi_1 _5404_ (.A1(_3283_),
    .A2(_3216_),
    .B1(_3276_),
    .B2(_3220_),
    .C1(_1907_),
    .Y(_1908_));
 sky130_fd_sc_hd__nand2_1 _5405_ (.A(_3282_),
    .B(_3334_),
    .Y(_1909_));
 sky130_fd_sc_hd__o21ai_1 _5406_ (.A1(_3328_),
    .A2(_3279_),
    .B1(_1909_),
    .Y(_1910_));
 sky130_fd_sc_hd__a221oi_1 _5407_ (.A1(_3311_),
    .A2(_3271_),
    .B1(_0772_),
    .B2(_3275_),
    .C1(_1910_),
    .Y(_1911_));
 sky130_fd_sc_hd__and4_1 _5408_ (.A(_1902_),
    .B(_1905_),
    .C(_1908_),
    .D(_1911_),
    .X(_1912_));
 sky130_fd_sc_hd__nand2_1 _5409_ (.A(_1899_),
    .B(_1912_),
    .Y(_1913_));
 sky130_fd_sc_hd__nor2_1 _5410_ (.A(_2986_),
    .B(_3123_),
    .Y(_1914_));
 sky130_fd_sc_hd__a22o_1 _5411_ (.A1(_3204_),
    .A2(_3112_),
    .B1(_3116_),
    .B2(_0746_),
    .X(_1915_));
 sky130_fd_sc_hd__a211oi_1 _5412_ (.A1(_3153_),
    .A2(_3127_),
    .B1(_1914_),
    .C1(_1915_),
    .Y(_1916_));
 sky130_fd_sc_hd__nand2_1 _5413_ (.A(_3061_),
    .B(_3070_),
    .Y(_1917_));
 sky130_fd_sc_hd__o21ai_1 _5414_ (.A1(_1025_),
    .A2(_3056_),
    .B1(_1917_),
    .Y(_1918_));
 sky130_fd_sc_hd__a221oi_1 _5415_ (.A1(_3109_),
    .A2(_3039_),
    .B1(_3118_),
    .B2(_3048_),
    .C1(_1918_),
    .Y(_1919_));
 sky130_fd_sc_hd__nand2_1 _5416_ (.A(_3099_),
    .B(_3169_),
    .Y(_1920_));
 sky130_fd_sc_hd__nand2_1 _5417_ (.A(_3093_),
    .B(_3075_),
    .Y(_1921_));
 sky130_fd_sc_hd__or2_1 _5418_ (.A(_1035_),
    .B(_3106_),
    .X(_1922_));
 sky130_fd_sc_hd__o2111a_1 _5419_ (.A1(_2980_),
    .A2(_3089_),
    .B1(_1920_),
    .C1(_1921_),
    .D1(_1922_),
    .X(_1923_));
 sky130_fd_sc_hd__nand2_1 _5420_ (.A(_3074_),
    .B(_3198_),
    .Y(_1924_));
 sky130_fd_sc_hd__o21ai_1 _5421_ (.A1(_2996_),
    .A2(_0729_),
    .B1(_1924_),
    .Y(_1925_));
 sky130_fd_sc_hd__a221oi_1 _5422_ (.A1(_0744_),
    .A2(_0726_),
    .B1(_3149_),
    .B2(_3081_),
    .C1(_1925_),
    .Y(_1926_));
 sky130_fd_sc_hd__and4_1 _5423_ (.A(_1916_),
    .B(_1919_),
    .C(_1923_),
    .D(_1926_),
    .X(_1927_));
 sky130_fd_sc_hd__nand2_1 _5424_ (.A(_3148_),
    .B(_1076_),
    .Y(_1928_));
 sky130_fd_sc_hd__o21ai_1 _5425_ (.A1(_0591_),
    .A2(_3145_),
    .B1(_1928_),
    .Y(_1929_));
 sky130_fd_sc_hd__a221oi_1 _5426_ (.A1(_0566_),
    .A2(_3137_),
    .B1(_0568_),
    .B2(_3141_),
    .C1(_1929_),
    .Y(_1930_));
 sky130_fd_sc_hd__nand2_1 _5427_ (.A(_3163_),
    .B(_3138_),
    .Y(_1931_));
 sky130_fd_sc_hd__nand2_1 _5428_ (.A(_3168_),
    .B(_3133_),
    .Y(_1932_));
 sky130_fd_sc_hd__nand2_1 _5429_ (.A(_1931_),
    .B(_1932_),
    .Y(_1933_));
 sky130_fd_sc_hd__a221oi_1 _5430_ (.A1(_3173_),
    .A2(_3156_),
    .B1(_3177_),
    .B2(_3160_),
    .C1(_1933_),
    .Y(_1934_));
 sky130_fd_sc_hd__a22o_1 _5431_ (.A1(_3181_),
    .A2(_0579_),
    .B1(_0562_),
    .B2(_3176_),
    .X(_1935_));
 sky130_fd_sc_hd__a221oi_1 _5432_ (.A1(_0553_),
    .A2(_3180_),
    .B1(_0585_),
    .B2(_3186_),
    .C1(_1935_),
    .Y(_1936_));
 sky130_fd_sc_hd__nand2_1 _5433_ (.A(_3203_),
    .B(_0741_),
    .Y(_1937_));
 sky130_fd_sc_hd__o21ai_1 _5434_ (.A1(_3024_),
    .A2(_3200_),
    .B1(_1937_),
    .Y(_1938_));
 sky130_fd_sc_hd__a221oi_1 _5435_ (.A1(_0623_),
    .A2(_3194_),
    .B1(_3197_),
    .B2(_0792_),
    .C1(_1938_),
    .Y(_1939_));
 sky130_fd_sc_hd__and4_1 _5436_ (.A(_1930_),
    .B(_1934_),
    .C(_1936_),
    .D(_1939_),
    .X(_1940_));
 sky130_fd_sc_hd__nand2_1 _5437_ (.A(_1927_),
    .B(_1940_),
    .Y(_1941_));
 sky130_fd_sc_hd__nor2_1 _5438_ (.A(_1913_),
    .B(_1941_),
    .Y(_1942_));
 sky130_fd_sc_hd__nand2_1 _5439_ (.A(_0622_),
    .B(_0583_),
    .Y(_1943_));
 sky130_fd_sc_hd__nand3_1 _5440_ (.A(_1885_),
    .B(_1942_),
    .C(_1943_),
    .Y(_1944_));
 sky130_fd_sc_hd__inv_2 _5441_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[5] ),
    .Y(_1945_));
 sky130_fd_sc_hd__a21oi_1 _5442_ (.A1(_1945_),
    .A2(_3027_),
    .B1(_2905_),
    .Y(_1946_));
 sky130_fd_sc_hd__o21a_1 _5443_ (.A1(_3027_),
    .A2(_1944_),
    .B1(_1946_),
    .X(_0287_));
 sky130_fd_sc_hd__o21ai_1 _5444_ (.A1(\egd_top.BitStream_buffer.BitStream_buffer_output[4] ),
    .A2(_2965_),
    .B1(_0627_),
    .Y(_1947_));
 sky130_fd_sc_hd__nand2_1 _5445_ (.A(_3333_),
    .B(_3062_),
    .Y(_1948_));
 sky130_fd_sc_hd__o21ai_1 _5446_ (.A1(_0796_),
    .A2(_3330_),
    .B1(_1948_),
    .Y(_1949_));
 sky130_fd_sc_hd__a221oi_1 _5447_ (.A1(_0716_),
    .A2(_3324_),
    .B1(_3326_),
    .B2(_3100_),
    .C1(_1949_),
    .Y(_1950_));
 sky130_fd_sc_hd__nand2_1 _5448_ (.A(_3291_),
    .B(_0785_),
    .Y(_1951_));
 sky130_fd_sc_hd__nand2_1 _5449_ (.A(_3294_),
    .B(_3338_),
    .Y(_1952_));
 sky130_fd_sc_hd__nand2_1 _5450_ (.A(_3300_),
    .B(_0330_),
    .Y(_1953_));
 sky130_fd_sc_hd__o2111a_1 _5451_ (.A1(_0850_),
    .A2(_3298_),
    .B1(_1951_),
    .C1(_1952_),
    .D1(_1953_),
    .X(_1954_));
 sky130_fd_sc_hd__nand2_1 _5452_ (.A(_3313_),
    .B(_3341_),
    .Y(_1955_));
 sky130_fd_sc_hd__nand2_1 _5453_ (.A(_3309_),
    .B(_3040_),
    .Y(_1956_));
 sky130_fd_sc_hd__or2_1 _5454_ (.A(_1016_),
    .B(_3318_),
    .X(_1957_));
 sky130_fd_sc_hd__o2111a_1 _5455_ (.A1(_3049_),
    .A2(_3308_),
    .B1(_1955_),
    .C1(_1956_),
    .D1(_1957_),
    .X(_1958_));
 sky130_fd_sc_hd__nand2_1 _5456_ (.A(_0328_),
    .B(_0714_),
    .Y(_1959_));
 sky130_fd_sc_hd__o21ai_1 _5457_ (.A1(_0718_),
    .A2(_0326_),
    .B1(_1959_),
    .Y(_1960_));
 sky130_fd_sc_hd__a221oi_1 _5458_ (.A1(_0722_),
    .A2(_3339_),
    .B1(_3109_),
    .B2(_0322_),
    .C1(_1960_),
    .Y(_1961_));
 sky130_fd_sc_hd__and4_1 _5459_ (.A(_1950_),
    .B(_1954_),
    .C(_1958_),
    .D(_1961_),
    .X(_1962_));
 sky130_fd_sc_hd__nand2_1 _5460_ (.A(_3126_),
    .B(_3157_),
    .Y(_1963_));
 sky130_fd_sc_hd__o21ai_1 _5461_ (.A1(_2990_),
    .A2(_3122_),
    .B1(_1963_),
    .Y(_1964_));
 sky130_fd_sc_hd__a221oi_1 _5462_ (.A1(_0746_),
    .A2(_3113_),
    .B1(_3117_),
    .B2(_3191_),
    .C1(_1964_),
    .Y(_1965_));
 sky130_fd_sc_hd__nand2_1 _5463_ (.A(_3038_),
    .B(_3118_),
    .Y(_1966_));
 sky130_fd_sc_hd__nand2_1 _5464_ (.A(_3047_),
    .B(_3066_),
    .Y(_1967_));
 sky130_fd_sc_hd__nand2_1 _5465_ (.A(_3060_),
    .B(_3075_),
    .Y(_1968_));
 sky130_fd_sc_hd__o2111a_1 _5466_ (.A1(_0727_),
    .A2(_3055_),
    .B1(_1966_),
    .C1(_1967_),
    .D1(_1968_),
    .X(_1969_));
 sky130_fd_sc_hd__nand2_1 _5467_ (.A(_3092_),
    .B(_3082_),
    .Y(_1970_));
 sky130_fd_sc_hd__nand2_1 _5468_ (.A(_3098_),
    .B(\egd_top.BitStream_buffer.BS_buffer[113] ),
    .Y(_1971_));
 sky130_fd_sc_hd__or2_1 _5469_ (.A(_2977_),
    .B(_3105_),
    .X(_1972_));
 sky130_fd_sc_hd__o2111a_1 _5470_ (.A1(_2983_),
    .A2(_3089_),
    .B1(_1970_),
    .C1(_1971_),
    .D1(_1972_),
    .X(_1973_));
 sky130_fd_sc_hd__nand2_1 _5471_ (.A(_3073_),
    .B(_0744_),
    .Y(_1974_));
 sky130_fd_sc_hd__o21ai_1 _5472_ (.A1(_2999_),
    .A2(_0729_),
    .B1(_1974_),
    .Y(_1975_));
 sky130_fd_sc_hd__a221oi_1 _5473_ (.A1(_3149_),
    .A2(_0726_),
    .B1(_3133_),
    .B2(_3080_),
    .C1(_1975_),
    .Y(_1976_));
 sky130_fd_sc_hd__and4_1 _5474_ (.A(_1965_),
    .B(_1969_),
    .C(_1973_),
    .D(_1976_),
    .X(_1977_));
 sky130_fd_sc_hd__nand2_1 _5475_ (.A(_3223_),
    .B(_3302_),
    .Y(_1978_));
 sky130_fd_sc_hd__o21ai_1 _5476_ (.A1(_0842_),
    .A2(_1145_),
    .B1(_1978_),
    .Y(_1979_));
 sky130_fd_sc_hd__a221oi_1 _5477_ (.A1(_3276_),
    .A2(_3216_),
    .B1(_0837_),
    .B2(_3220_),
    .C1(_1979_),
    .Y(_1980_));
 sky130_fd_sc_hd__nand2_1 _5478_ (.A(_3242_),
    .B(\egd_top.BitStream_buffer.BS_buffer[75] ),
    .Y(_1981_));
 sky130_fd_sc_hd__nand2_1 _5479_ (.A(_3232_),
    .B(_3272_),
    .Y(_1982_));
 sky130_fd_sc_hd__nand2_1 _5480_ (.A(_3235_),
    .B(_3283_),
    .Y(_1983_));
 sky130_fd_sc_hd__o2111a_1 _5481_ (.A1(_1149_),
    .A2(_3240_),
    .B1(_1981_),
    .C1(_1982_),
    .D1(_1983_),
    .X(_1984_));
 sky130_fd_sc_hd__nand2_1 _5482_ (.A(_3254_),
    .B(_3311_),
    .Y(_1985_));
 sky130_fd_sc_hd__nand2_1 _5483_ (.A(_3262_),
    .B(\egd_top.BitStream_buffer.BS_buffer[84] ),
    .Y(_1986_));
 sky130_fd_sc_hd__nand2_1 _5484_ (.A(_3259_),
    .B(\egd_top.BitStream_buffer.BS_buffer[83] ),
    .Y(_1987_));
 sky130_fd_sc_hd__nand2_1 _5485_ (.A(_3250_),
    .B(\egd_top.BitStream_buffer.BS_buffer[85] ),
    .Y(_1988_));
 sky130_fd_sc_hd__and4_1 _5486_ (.A(_1985_),
    .B(_1986_),
    .C(_1987_),
    .D(_1988_),
    .X(_1989_));
 sky130_fd_sc_hd__nand2_1 _5487_ (.A(_3281_),
    .B(_0780_),
    .Y(_1990_));
 sky130_fd_sc_hd__o21ai_1 _5488_ (.A1(_0779_),
    .A2(_3279_),
    .B1(_1990_),
    .Y(_1991_));
 sky130_fd_sc_hd__a221oi_1 _5489_ (.A1(_0772_),
    .A2(_3270_),
    .B1(_3334_),
    .B2(_3275_),
    .C1(_1991_),
    .Y(_1992_));
 sky130_fd_sc_hd__and4_1 _5490_ (.A(_1980_),
    .B(_1984_),
    .C(_1989_),
    .D(_1992_),
    .X(_1993_));
 sky130_fd_sc_hd__nand2_1 _5491_ (.A(_3203_),
    .B(_3187_),
    .Y(_1994_));
 sky130_fd_sc_hd__o21ai_1 _5492_ (.A1(_1602_),
    .A2(_3200_),
    .B1(_1994_),
    .Y(_1995_));
 sky130_fd_sc_hd__a221oi_1 _5493_ (.A1(_0792_),
    .A2(_3194_),
    .B1(_3197_),
    .B2(_0930_),
    .C1(_1995_),
    .Y(_1996_));
 sky130_fd_sc_hd__nand2_1 _5494_ (.A(_3162_),
    .B(\egd_top.BitStream_buffer.BS_buffer[124] ),
    .Y(_1997_));
 sky130_fd_sc_hd__nand2_1 _5495_ (.A(_3159_),
    .B(_0741_),
    .Y(_1998_));
 sky130_fd_sc_hd__nand2_1 _5496_ (.A(_3167_),
    .B(\egd_top.BitStream_buffer.BS_buffer[123] ),
    .Y(_1999_));
 sky130_fd_sc_hd__nand2_1 _5497_ (.A(_3155_),
    .B(\egd_top.BitStream_buffer.BS_buffer[125] ),
    .Y(_2000_));
 sky130_fd_sc_hd__and4_1 _5498_ (.A(_1997_),
    .B(_1998_),
    .C(_1999_),
    .D(_2000_),
    .X(_2001_));
 sky130_fd_sc_hd__nand2_1 _5499_ (.A(_3147_),
    .B(_0566_),
    .Y(_2002_));
 sky130_fd_sc_hd__nand2_1 _5500_ (.A(_3140_),
    .B(_0562_),
    .Y(_2003_));
 sky130_fd_sc_hd__nand2_1 _5501_ (.A(_3144_),
    .B(_1076_),
    .Y(_2004_));
 sky130_fd_sc_hd__nand2_1 _5502_ (.A(_3136_),
    .B(_0568_),
    .Y(_2005_));
 sky130_fd_sc_hd__and4_1 _5503_ (.A(_2002_),
    .B(_2003_),
    .C(_2004_),
    .D(_2005_),
    .X(_2006_));
 sky130_fd_sc_hd__nand2_1 _5504_ (.A(_3175_),
    .B(_0553_),
    .Y(_2007_));
 sky130_fd_sc_hd__o21ai_1 _5505_ (.A1(_0586_),
    .A2(_3183_),
    .B1(_2007_),
    .Y(_2008_));
 sky130_fd_sc_hd__a221oi_1 _5506_ (.A1(_3186_),
    .A2(_0583_),
    .B1(_0579_),
    .B2(_3180_),
    .C1(_2008_),
    .Y(_2009_));
 sky130_fd_sc_hd__and4_1 _5507_ (.A(_1996_),
    .B(_2001_),
    .C(_2006_),
    .D(_2009_),
    .X(_2010_));
 sky130_fd_sc_hd__and4_1 _5508_ (.A(_1962_),
    .B(_1977_),
    .C(_1993_),
    .D(_2010_),
    .X(_2011_));
 sky130_fd_sc_hd__nand2_1 _5509_ (.A(_0353_),
    .B(_0948_),
    .Y(_2012_));
 sky130_fd_sc_hd__o21ai_1 _5510_ (.A1(_0659_),
    .A2(_0350_),
    .B1(_2012_),
    .Y(_2013_));
 sky130_fd_sc_hd__a221oi_1 _5511_ (.A1(_0642_),
    .A2(_0342_),
    .B1(_0345_),
    .B2(_0874_),
    .C1(_2013_),
    .Y(_2014_));
 sky130_fd_sc_hd__nand2_1 _5512_ (.A(_0371_),
    .B(_0869_),
    .Y(_2015_));
 sky130_fd_sc_hd__o21ai_1 _5513_ (.A1(_0637_),
    .A2(_0368_),
    .B1(_2015_),
    .Y(_2016_));
 sky130_fd_sc_hd__a221oi_1 _5514_ (.A1(_0400_),
    .A2(_0360_),
    .B1(_0363_),
    .B2(_0407_),
    .C1(_2016_),
    .Y(_2017_));
 sky130_fd_sc_hd__nand2_1 _5515_ (.A(_0377_),
    .B(_0416_),
    .Y(_2018_));
 sky130_fd_sc_hd__o21ai_1 _5516_ (.A1(_0960_),
    .A2(_0380_),
    .B1(_2018_),
    .Y(_2019_));
 sky130_fd_sc_hd__a221oi_1 _5517_ (.A1(_0655_),
    .A2(_0388_),
    .B1(_0429_),
    .B2(_0944_),
    .C1(_2019_),
    .Y(_2020_));
 sky130_fd_sc_hd__nand2_1 _5518_ (.A(_0406_),
    .B(_0461_),
    .Y(_2021_));
 sky130_fd_sc_hd__o21ai_1 _5519_ (.A1(_0650_),
    .A2(_0403_),
    .B1(_2021_),
    .Y(_2022_));
 sky130_fd_sc_hd__a221oi_1 _5520_ (.A1(_0436_),
    .A2(_0396_),
    .B1(_0399_),
    .B2(_0454_),
    .C1(_2022_),
    .Y(_2023_));
 sky130_fd_sc_hd__and4_1 _5521_ (.A(_2014_),
    .B(_2017_),
    .C(_2020_),
    .D(_2023_),
    .X(_2024_));
 sky130_fd_sc_hd__or2_1 _5522_ (.A(_0448_),
    .B(_0425_),
    .X(_2025_));
 sky130_fd_sc_hd__o21ai_1 _5523_ (.A1(_0647_),
    .A2(_0422_),
    .B1(_2025_),
    .Y(_2026_));
 sky130_fd_sc_hd__a221oi_1 _5524_ (.A1(_0471_),
    .A2(_0415_),
    .B1(_0478_),
    .B2(_0419_),
    .C1(_2026_),
    .Y(_2027_));
 sky130_fd_sc_hd__nand2_1 _5525_ (.A(_0442_),
    .B(_0664_),
    .Y(_2028_));
 sky130_fd_sc_hd__o21ai_1 _5526_ (.A1(_0663_),
    .A2(_0439_),
    .B1(_2028_),
    .Y(_2029_));
 sky130_fd_sc_hd__a221oi_1 _5527_ (.A1(_0751_),
    .A2(_0432_),
    .B1(_0435_),
    .B2(_3230_),
    .C1(_2029_),
    .Y(_2030_));
 sky130_fd_sc_hd__nand2_1 _5528_ (.A(_0453_),
    .B(_3237_),
    .Y(_2031_));
 sky130_fd_sc_hd__nand2_1 _5529_ (.A(_0458_),
    .B(_3217_),
    .Y(_2032_));
 sky130_fd_sc_hd__or2_1 _5530_ (.A(_0755_),
    .B(_0449_),
    .X(_2033_));
 sky130_fd_sc_hd__o2111a_1 _5531_ (.A1(_1043_),
    .A2(_0464_),
    .B1(_2031_),
    .C1(_2032_),
    .D1(_2033_),
    .X(_2034_));
 sky130_fd_sc_hd__nand2_1 _5532_ (.A(_0469_),
    .B(_3227_),
    .Y(_2035_));
 sky130_fd_sc_hd__o21ai_1 _5533_ (.A1(_3257_),
    .A2(_0472_),
    .B1(_2035_),
    .Y(_2036_));
 sky130_fd_sc_hd__a221oi_1 _5534_ (.A1(_3264_),
    .A2(_0477_),
    .B1(_3248_),
    .B2(_2936_),
    .C1(_2036_),
    .Y(_2037_));
 sky130_fd_sc_hd__and4_1 _5535_ (.A(_2027_),
    .B(_2030_),
    .C(_2034_),
    .D(_2037_),
    .X(_2038_));
 sky130_fd_sc_hd__nand2_1 _5536_ (.A(_2024_),
    .B(_2038_),
    .Y(_2039_));
 sky130_fd_sc_hd__nand2_1 _5537_ (.A(_0497_),
    .B(_0537_),
    .Y(_2040_));
 sky130_fd_sc_hd__o21ai_1 _5538_ (.A1(_0543_),
    .A2(_0495_),
    .B1(_2040_),
    .Y(_2041_));
 sky130_fd_sc_hd__a221oi_1 _5539_ (.A1(\egd_top.BitStream_buffer.BS_buffer[27] ),
    .A2(_0487_),
    .B1(\egd_top.BitStream_buffer.BS_buffer[28] ),
    .B2(_0490_),
    .C1(_2041_),
    .Y(_2042_));
 sky130_fd_sc_hd__nand2_1 _5540_ (.A(_0514_),
    .B(_0365_),
    .Y(_2043_));
 sky130_fd_sc_hd__o21ai_1 _5541_ (.A1(_0633_),
    .A2(_0512_),
    .B1(_2043_),
    .Y(_2044_));
 sky130_fd_sc_hd__a221oi_1 _5542_ (.A1(_0540_),
    .A2(_0504_),
    .B1(\egd_top.BitStream_buffer.BS_buffer[32] ),
    .B2(_0508_),
    .C1(_2044_),
    .Y(_2045_));
 sky130_fd_sc_hd__o22a_1 _5543_ (.A1(_0940_),
    .A2(_0530_),
    .B1(_1084_),
    .B2(_0534_),
    .X(_2046_));
 sky130_fd_sc_hd__o221a_1 _5544_ (.A1(_0865_),
    .A2(_0523_),
    .B1(_1276_),
    .B2(_0526_),
    .C1(_2046_),
    .X(_2047_));
 sky130_fd_sc_hd__nand2_1 _5545_ (.A(_0548_),
    .B(_0347_),
    .Y(_2048_));
 sky130_fd_sc_hd__o21ai_1 _5546_ (.A1(_0629_),
    .A2(_0546_),
    .B1(_2048_),
    .Y(_2049_));
 sky130_fd_sc_hd__a221oi_1 _5547_ (.A1(_0379_),
    .A2(_0539_),
    .B1(_0389_),
    .B2(_0542_),
    .C1(_2049_),
    .Y(_2050_));
 sky130_fd_sc_hd__and4_1 _5548_ (.A(_2042_),
    .B(_2045_),
    .C(_2047_),
    .D(_2050_),
    .X(_2051_));
 sky130_fd_sc_hd__nand2_1 _5549_ (.A(_0561_),
    .B(\egd_top.BitStream_buffer.BS_buffer[17] ),
    .Y(_2052_));
 sky130_fd_sc_hd__nand2_1 _5550_ (.A(_0565_),
    .B(\egd_top.BitStream_buffer.BS_buffer[15] ),
    .Y(_2053_));
 sky130_fd_sc_hd__or2_1 _5551_ (.A(_0685_),
    .B(_0571_),
    .X(_2054_));
 sky130_fd_sc_hd__o2111a_1 _5552_ (.A1(_0492_),
    .A2(_0558_),
    .B1(_2052_),
    .C1(_2053_),
    .D1(_2054_),
    .X(_2055_));
 sky130_fd_sc_hd__nand2_1 _5553_ (.A(_0578_),
    .B(_0498_),
    .Y(_2056_));
 sky130_fd_sc_hd__nand2_1 _5554_ (.A(_0582_),
    .B(_0505_),
    .Y(_2057_));
 sky130_fd_sc_hd__or2_1 _5555_ (.A(_0897_),
    .B(_0588_),
    .X(_2058_));
 sky130_fd_sc_hd__o2111a_1 _5556_ (.A1(_1128_),
    .A2(_0576_),
    .B1(_2056_),
    .C1(_2057_),
    .D1(_2058_),
    .X(_2059_));
 sky130_fd_sc_hd__or2_1 _5557_ (.A(_0688_),
    .B(_0599_),
    .X(_2060_));
 sky130_fd_sc_hd__o221a_1 _5558_ (.A1(_0611_),
    .A2(_0593_),
    .B1(_0676_),
    .B2(_0596_),
    .C1(_2060_),
    .X(_2061_));
 sky130_fd_sc_hd__nand2_1 _5559_ (.A(_0606_),
    .B(_0509_),
    .Y(_2062_));
 sky130_fd_sc_hd__nand2_1 _5560_ (.A(_0609_),
    .B(_0527_),
    .Y(_2063_));
 sky130_fd_sc_hd__or2_1 _5561_ (.A(_0520_),
    .B(_0613_),
    .X(_2064_));
 sky130_fd_sc_hd__o2111a_1 _5562_ (.A1(_0532_),
    .A2(_0604_),
    .B1(_2062_),
    .C1(_2063_),
    .D1(_2064_),
    .X(_2065_));
 sky130_fd_sc_hd__and4_1 _5563_ (.A(_2055_),
    .B(_2059_),
    .C(_2061_),
    .D(_2065_),
    .X(_2066_));
 sky130_fd_sc_hd__nand2_1 _5564_ (.A(_2051_),
    .B(_2066_),
    .Y(_2067_));
 sky130_fd_sc_hd__nor2_1 _5565_ (.A(_2039_),
    .B(_2067_),
    .Y(_2068_));
 sky130_fd_sc_hd__nand2_1 _5566_ (.A(_0621_),
    .B(\egd_top.BitStream_buffer.BS_buffer[11] ),
    .Y(_2069_));
 sky130_fd_sc_hd__nand3_1 _5567_ (.A(_2011_),
    .B(_2068_),
    .C(_2069_),
    .Y(_2070_));
 sky130_fd_sc_hd__nor2_1 _5568_ (.A(_3026_),
    .B(_2070_),
    .Y(_2071_));
 sky130_fd_sc_hd__nor2_1 _5569_ (.A(_1947_),
    .B(_2071_),
    .Y(_0286_));
 sky130_fd_sc_hd__o21ai_1 _5570_ (.A1(\egd_top.BitStream_buffer.BitStream_buffer_output[3] ),
    .A2(_2965_),
    .B1(_0627_),
    .Y(_2072_));
 sky130_fd_sc_hd__nand2_1 _5571_ (.A(_0371_),
    .B(_0393_),
    .Y(_2073_));
 sky130_fd_sc_hd__o21ai_1 _5572_ (.A1(_0870_),
    .A2(_0368_),
    .B1(_2073_),
    .Y(_2074_));
 sky130_fd_sc_hd__a221oi_1 _5573_ (.A1(_0407_),
    .A2(_0360_),
    .B1(_0363_),
    .B2(_0642_),
    .C1(_2074_),
    .Y(_2075_));
 sky130_fd_sc_hd__nand2_1 _5574_ (.A(_0387_),
    .B(_0429_),
    .Y(_2076_));
 sky130_fd_sc_hd__o21ai_1 _5575_ (.A1(_0883_),
    .A2(_0385_),
    .B1(_2076_),
    .Y(_2077_));
 sky130_fd_sc_hd__a221oi_1 _5576_ (.A1(_0443_),
    .A2(_0378_),
    .B1(_0655_),
    .B2(_0382_),
    .C1(_2077_),
    .Y(_2078_));
 sky130_fd_sc_hd__a22o_1 _5577_ (.A1(\egd_top.BitStream_buffer.BS_buffer[48] ),
    .A2(_0341_),
    .B1(_0344_),
    .B2(_0948_),
    .X(_2079_));
 sky130_fd_sc_hd__a32o_1 _5578_ (.A1(_3087_),
    .A2(_0416_),
    .A3(_0339_),
    .B1(_0412_),
    .B2(_0352_),
    .X(_2080_));
 sky130_fd_sc_hd__nor2_1 _5579_ (.A(_2079_),
    .B(_2080_),
    .Y(_2081_));
 sky130_fd_sc_hd__nand2_1 _5580_ (.A(_0405_),
    .B(_0459_),
    .Y(_2082_));
 sky130_fd_sc_hd__o21ai_1 _5581_ (.A1(_0448_),
    .A2(_0402_),
    .B1(_2082_),
    .Y(_2083_));
 sky130_fd_sc_hd__a221oi_1 _5582_ (.A1(_0454_),
    .A2(_0395_),
    .B1(_0398_),
    .B2(_0461_),
    .C1(_2083_),
    .Y(_2084_));
 sky130_fd_sc_hd__and4_1 _5583_ (.A(_2075_),
    .B(_2078_),
    .C(_2081_),
    .D(_2084_),
    .X(_2085_));
 sky130_fd_sc_hd__or2_1 _5584_ (.A(_0647_),
    .B(_0424_),
    .X(_2086_));
 sky130_fd_sc_hd__o21ai_1 _5585_ (.A1(_0887_),
    .A2(_0421_),
    .B1(_2086_),
    .Y(_2087_));
 sky130_fd_sc_hd__a221oi_1 _5586_ (.A1(_0478_),
    .A2(_0414_),
    .B1(_0664_),
    .B2(_0418_),
    .C1(_2087_),
    .Y(_2088_));
 sky130_fd_sc_hd__nand2_1 _5587_ (.A(_0452_),
    .B(_3210_),
    .Y(_2089_));
 sky130_fd_sc_hd__nand2_1 _5588_ (.A(_0457_),
    .B(_3221_),
    .Y(_2090_));
 sky130_fd_sc_hd__or2_1 _5589_ (.A(_1360_),
    .B(_0463_),
    .X(_2091_));
 sky130_fd_sc_hd__o2111a_1 _5590_ (.A1(_1430_),
    .A2(_0450_),
    .B1(_2089_),
    .C1(_2090_),
    .D1(_2091_),
    .X(_2092_));
 sky130_fd_sc_hd__nand2_1 _5591_ (.A(_0441_),
    .B(_3244_),
    .Y(_2093_));
 sky130_fd_sc_hd__nand2_1 _5592_ (.A(_0432_),
    .B(_3230_),
    .Y(_2094_));
 sky130_fd_sc_hd__nand2_1 _5593_ (.A(_0434_),
    .B(_3237_),
    .Y(_2095_));
 sky130_fd_sc_hd__o2111a_1 _5594_ (.A1(_3238_),
    .A2(_0439_),
    .B1(_2093_),
    .C1(_2094_),
    .D1(_2095_),
    .X(_2096_));
 sky130_fd_sc_hd__nand2_1 _5595_ (.A(_0476_),
    .B(\egd_top.BitStream_buffer.BS_buffer[74] ),
    .Y(_2097_));
 sky130_fd_sc_hd__o21ai_1 _5596_ (.A1(_1144_),
    .A2(_2935_),
    .B1(_2097_),
    .Y(_2098_));
 sky130_fd_sc_hd__a221oi_1 _5597_ (.A1(_3256_),
    .A2(_0470_),
    .B1(_3264_),
    .B2(_0473_),
    .C1(_2098_),
    .Y(_2099_));
 sky130_fd_sc_hd__and4_1 _5598_ (.A(_2088_),
    .B(_2092_),
    .C(_2096_),
    .D(_2099_),
    .X(_2100_));
 sky130_fd_sc_hd__nand2_1 _5599_ (.A(_0560_),
    .B(_0491_),
    .Y(_2101_));
 sky130_fd_sc_hd__nand2_1 _5600_ (.A(_0564_),
    .B(\egd_top.BitStream_buffer.BS_buffer[16] ),
    .Y(_2102_));
 sky130_fd_sc_hd__or2_1 _5601_ (.A(_0922_),
    .B(_0570_),
    .X(_2103_));
 sky130_fd_sc_hd__o2111a_1 _5602_ (.A1(_0692_),
    .A2(_0557_),
    .B1(_2101_),
    .C1(_2102_),
    .D1(_2103_),
    .X(_2104_));
 sky130_fd_sc_hd__nand2_1 _5603_ (.A(_0577_),
    .B(_0502_),
    .Y(_2105_));
 sky130_fd_sc_hd__nand2_1 _5604_ (.A(_0581_),
    .B(_0515_),
    .Y(_2106_));
 sky130_fd_sc_hd__or2_1 _5605_ (.A(_0510_),
    .B(_0575_),
    .X(_2107_));
 sky130_fd_sc_hd__o2111a_1 _5606_ (.A1(_0986_),
    .A2(_0588_),
    .B1(_2105_),
    .C1(_2106_),
    .D1(_2107_),
    .X(_2108_));
 sky130_fd_sc_hd__or2_1 _5607_ (.A(_0602_),
    .B(_0598_),
    .X(_2109_));
 sky130_fd_sc_hd__o221a_1 _5608_ (.A1(_0688_),
    .A2(_0592_),
    .B1(_0611_),
    .B2(_0596_),
    .C1(_2109_),
    .X(_2110_));
 sky130_fd_sc_hd__nand2_1 _5609_ (.A(_0608_),
    .B(_0531_),
    .Y(_2111_));
 sky130_fd_sc_hd__nand2_1 _5610_ (.A(_0605_),
    .B(_0519_),
    .Y(_2112_));
 sky130_fd_sc_hd__or2_1 _5611_ (.A(_0528_),
    .B(_0612_),
    .X(_2113_));
 sky130_fd_sc_hd__o2111a_1 _5612_ (.A1(_0524_),
    .A2(_0603_),
    .B1(_2111_),
    .C1(_2112_),
    .D1(_2113_),
    .X(_2114_));
 sky130_fd_sc_hd__and4_1 _5613_ (.A(_2104_),
    .B(_2108_),
    .C(_2110_),
    .D(_2114_),
    .X(_2115_));
 sky130_fd_sc_hd__nand2_1 _5614_ (.A(_0486_),
    .B(\egd_top.BitStream_buffer.BS_buffer[28] ),
    .Y(_2116_));
 sky130_fd_sc_hd__nand2_1 _5615_ (.A(_0496_),
    .B(_0540_),
    .Y(_2117_));
 sky130_fd_sc_hd__nand2_1 _5616_ (.A(_0489_),
    .B(\egd_top.BitStream_buffer.BS_buffer[29] ),
    .Y(_2118_));
 sky130_fd_sc_hd__o2111a_1 _5617_ (.A1(_0702_),
    .A2(_0494_),
    .B1(_2116_),
    .C1(_2117_),
    .D1(_2118_),
    .X(_2119_));
 sky130_fd_sc_hd__nand2_1 _5618_ (.A(_0503_),
    .B(\egd_top.BitStream_buffer.BS_buffer[32] ),
    .Y(_2120_));
 sky130_fd_sc_hd__nand2_1 _5619_ (.A(_0513_),
    .B(\egd_top.BitStream_buffer.BS_buffer[34] ),
    .Y(_2121_));
 sky130_fd_sc_hd__nand2_1 _5620_ (.A(_0507_),
    .B(_0365_),
    .Y(_2122_));
 sky130_fd_sc_hd__o2111a_1 _5621_ (.A1(_0865_),
    .A2(_0511_),
    .B1(_2120_),
    .C1(_2121_),
    .D1(_2122_),
    .X(_2123_));
 sky130_fd_sc_hd__nand2_1 _5622_ (.A(_0547_),
    .B(_0375_),
    .Y(_2124_));
 sky130_fd_sc_hd__o21ai_1 _5623_ (.A1(_0861_),
    .A2(_0545_),
    .B1(_2124_),
    .Y(_2125_));
 sky130_fd_sc_hd__a221oi_1 _5624_ (.A1(_0389_),
    .A2(_0538_),
    .B1(_0869_),
    .B2(_0541_),
    .C1(_2125_),
    .Y(_2126_));
 sky130_fd_sc_hd__o22a_1 _5625_ (.A1(_1084_),
    .A2(_0529_),
    .B1(_0348_),
    .B2(_0525_),
    .X(_2127_));
 sky130_fd_sc_hd__o221a_1 _5626_ (.A1(_0940_),
    .A2(_0522_),
    .B1(_1276_),
    .B2(_0533_),
    .C1(_2127_),
    .X(_2128_));
 sky130_fd_sc_hd__and4_1 _5627_ (.A(_2119_),
    .B(_2123_),
    .C(_2126_),
    .D(_2128_),
    .X(_2129_));
 sky130_fd_sc_hd__and4_1 _5628_ (.A(_2085_),
    .B(_2100_),
    .C(_2115_),
    .D(_2129_),
    .X(_2130_));
 sky130_fd_sc_hd__nand2_1 _5629_ (.A(_3301_),
    .B(_0785_),
    .Y(_2131_));
 sky130_fd_sc_hd__o21ai_1 _5630_ (.A1(_1003_),
    .A2(_3299_),
    .B1(_2131_),
    .Y(_2132_));
 sky130_fd_sc_hd__a221oi_2 _5631_ (.A1(_3338_),
    .A2(_3292_),
    .B1(_3341_),
    .B2(_3295_),
    .C1(_2132_),
    .Y(_2133_));
 sky130_fd_sc_hd__nand2_1 _5632_ (.A(_3310_),
    .B(_0708_),
    .Y(_2134_));
 sky130_fd_sc_hd__nand2_1 _5633_ (.A(_3314_),
    .B(_3028_),
    .Y(_2135_));
 sky130_fd_sc_hd__or2_1 _5634_ (.A(_1169_),
    .B(_3319_),
    .X(_2136_));
 sky130_fd_sc_hd__o2111a_1 _5635_ (.A1(_0709_),
    .A2(_3308_),
    .B1(_2134_),
    .C1(_2135_),
    .D1(_2136_),
    .X(_2137_));
 sky130_fd_sc_hd__nand2_1 _5636_ (.A(_3333_),
    .B(_3094_),
    .Y(_2138_));
 sky130_fd_sc_hd__o21ai_1 _5637_ (.A1(_3102_),
    .A2(_3330_),
    .B1(_2138_),
    .Y(_2139_));
 sky130_fd_sc_hd__a221oi_1 _5638_ (.A1(_3100_),
    .A2(_3324_),
    .B1(_3326_),
    .B2(_0714_),
    .C1(_2139_),
    .Y(_2140_));
 sky130_fd_sc_hd__nand2_1 _5639_ (.A(_0329_),
    .B(_3128_),
    .Y(_2141_));
 sky130_fd_sc_hd__o21ai_1 _5640_ (.A1(_3119_),
    .A2(_0327_),
    .B1(_2141_),
    .Y(_2142_));
 sky130_fd_sc_hd__a221oi_1 _5641_ (.A1(_3109_),
    .A2(_3340_),
    .B1(_3118_),
    .B2(_0323_),
    .C1(_2142_),
    .Y(_2143_));
 sky130_fd_sc_hd__and4_1 _5642_ (.A(_2133_),
    .B(_2137_),
    .C(_2140_),
    .D(_2143_),
    .X(_2144_));
 sky130_fd_sc_hd__nand2_1 _5643_ (.A(_3263_),
    .B(_0774_),
    .Y(_2145_));
 sky130_fd_sc_hd__o21ai_1 _5644_ (.A1(_1158_),
    .A2(_3260_),
    .B1(_2145_),
    .Y(_2146_));
 sky130_fd_sc_hd__a221oi_1 _5645_ (.A1(_3311_),
    .A2(_3251_),
    .B1(_0772_),
    .B2(_3255_),
    .C1(_2146_),
    .Y(_2147_));
 sky130_fd_sc_hd__nand2_1 _5646_ (.A(_3243_),
    .B(_3268_),
    .Y(_2148_));
 sky130_fd_sc_hd__o21ai_1 _5647_ (.A1(_1426_),
    .A2(_3240_),
    .B1(_2148_),
    .Y(_2149_));
 sky130_fd_sc_hd__a221oi_1 _5648_ (.A1(_3283_),
    .A2(_3233_),
    .B1(_3236_),
    .B2(_3276_),
    .C1(_2149_),
    .Y(_2150_));
 sky130_fd_sc_hd__nand2_1 _5649_ (.A(_3224_),
    .B(_3288_),
    .Y(_2151_));
 sky130_fd_sc_hd__o21ai_1 _5650_ (.A1(_1007_),
    .A2(_1145_),
    .B1(_2151_),
    .Y(_2152_));
 sky130_fd_sc_hd__a221oi_1 _5651_ (.A1(_0837_),
    .A2(_3216_),
    .B1(_3302_),
    .B2(_3220_),
    .C1(_2152_),
    .Y(_2153_));
 sky130_fd_sc_hd__a22o_1 _5652_ (.A1(_3322_),
    .A2(_3281_),
    .B1(_1153_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[91] ),
    .X(_2154_));
 sky130_fd_sc_hd__a221oi_1 _5653_ (.A1(_3334_),
    .A2(_3271_),
    .B1(_0780_),
    .B2(_3275_),
    .C1(_2154_),
    .Y(_2155_));
 sky130_fd_sc_hd__and4_1 _5654_ (.A(_2147_),
    .B(_2150_),
    .C(_2153_),
    .D(_2155_),
    .X(_2156_));
 sky130_fd_sc_hd__nand2_1 _5655_ (.A(_2144_),
    .B(_2156_),
    .Y(_2157_));
 sky130_fd_sc_hd__a22o_1 _5656_ (.A1(_0562_),
    .A2(_3137_),
    .B1(_3141_),
    .B2(_0553_),
    .X(_2158_));
 sky130_fd_sc_hd__a221oi_1 _5657_ (.A1(_0566_),
    .A2(_3144_),
    .B1(_0568_),
    .B2(_3148_),
    .C1(_2158_),
    .Y(_2159_));
 sky130_fd_sc_hd__nand2_1 _5658_ (.A(_3163_),
    .B(_3177_),
    .Y(_2160_));
 sky130_fd_sc_hd__nand2_1 _5659_ (.A(_3168_),
    .B(_3173_),
    .Y(_2161_));
 sky130_fd_sc_hd__nand2_1 _5660_ (.A(_2160_),
    .B(_2161_),
    .Y(_2162_));
 sky130_fd_sc_hd__a221oi_1 _5661_ (.A1(_0741_),
    .A2(_3156_),
    .B1(_3187_),
    .B2(_3160_),
    .C1(_2162_),
    .Y(_2163_));
 sky130_fd_sc_hd__nand2_1 _5662_ (.A(_3203_),
    .B(_0623_),
    .Y(_2164_));
 sky130_fd_sc_hd__o21ai_1 _5663_ (.A1(_0594_),
    .A2(_3200_),
    .B1(_2164_),
    .Y(_2165_));
 sky130_fd_sc_hd__a221oi_1 _5664_ (.A1(_0930_),
    .A2(_3194_),
    .B1(_3197_),
    .B2(_1076_),
    .C1(_2165_),
    .Y(_2166_));
 sky130_fd_sc_hd__nand2_1 _5665_ (.A(_3186_),
    .B(\egd_top.BitStream_buffer.BS_buffer[11] ),
    .Y(_2167_));
 sky130_fd_sc_hd__o21ai_1 _5666_ (.A1(_0679_),
    .A2(_3183_),
    .B1(_2167_),
    .Y(_2168_));
 sky130_fd_sc_hd__a221oi_1 _5667_ (.A1(_0579_),
    .A2(_3176_),
    .B1(_0585_),
    .B2(_3180_),
    .C1(_2168_),
    .Y(_2169_));
 sky130_fd_sc_hd__and4_1 _5668_ (.A(_2159_),
    .B(_2163_),
    .C(_2166_),
    .D(_2169_),
    .X(_2170_));
 sky130_fd_sc_hd__nand2_1 _5669_ (.A(_3061_),
    .B(_3082_),
    .Y(_2171_));
 sky130_fd_sc_hd__o21ai_1 _5670_ (.A1(_0808_),
    .A2(_3056_),
    .B1(_2171_),
    .Y(_2172_));
 sky130_fd_sc_hd__a221oi_1 _5671_ (.A1(_3066_),
    .A2(_3039_),
    .B1(_3070_),
    .B2(_3048_),
    .C1(_2172_),
    .Y(_2173_));
 sky130_fd_sc_hd__nand2_1 _5672_ (.A(_3099_),
    .B(_3153_),
    .Y(_2174_));
 sky130_fd_sc_hd__nand2_1 _5673_ (.A(_3093_),
    .B(_3169_),
    .Y(_2175_));
 sky130_fd_sc_hd__or2_1 _5674_ (.A(_2986_),
    .B(_3088_),
    .X(_2176_));
 sky130_fd_sc_hd__o2111a_1 _5675_ (.A1(_2980_),
    .A2(_3106_),
    .B1(_2174_),
    .C1(_2175_),
    .D1(_2176_),
    .X(_2177_));
 sky130_fd_sc_hd__nand2_1 _5676_ (.A(_3127_),
    .B(_3204_),
    .Y(_2178_));
 sky130_fd_sc_hd__o21ai_1 _5677_ (.A1(_2993_),
    .A2(_3123_),
    .B1(_2178_),
    .Y(_2179_));
 sky130_fd_sc_hd__a221oi_1 _5678_ (.A1(_3191_),
    .A2(_3113_),
    .B1(_3117_),
    .B2(_3198_),
    .C1(_2179_),
    .Y(_2180_));
 sky130_fd_sc_hd__nand2_1 _5679_ (.A(_3074_),
    .B(_3149_),
    .Y(_2181_));
 sky130_fd_sc_hd__o21ai_1 _5680_ (.A1(_3003_),
    .A2(_0729_),
    .B1(_2181_),
    .Y(_2182_));
 sky130_fd_sc_hd__a221oi_1 _5681_ (.A1(_3133_),
    .A2(_0726_),
    .B1(_3138_),
    .B2(_3081_),
    .C1(_2182_),
    .Y(_2183_));
 sky130_fd_sc_hd__and4_1 _5682_ (.A(_2173_),
    .B(_2177_),
    .C(_2180_),
    .D(_2183_),
    .X(_2184_));
 sky130_fd_sc_hd__nand2_1 _5683_ (.A(_2170_),
    .B(_2184_),
    .Y(_2185_));
 sky130_fd_sc_hd__nor2_1 _5684_ (.A(_2157_),
    .B(_2185_),
    .Y(_2186_));
 sky130_fd_sc_hd__nand2_1 _5685_ (.A(_0621_),
    .B(\egd_top.BitStream_buffer.BS_buffer[12] ),
    .Y(_2187_));
 sky130_fd_sc_hd__nand3_1 _5686_ (.A(_2130_),
    .B(_2186_),
    .C(_2187_),
    .Y(_2188_));
 sky130_fd_sc_hd__nor2_1 _5687_ (.A(_3026_),
    .B(_2188_),
    .Y(_2189_));
 sky130_fd_sc_hd__nor2_1 _5688_ (.A(_2072_),
    .B(_2189_),
    .Y(_0285_));
 sky130_fd_sc_hd__o21ai_1 _5689_ (.A1(\egd_top.BitStream_buffer.BitStream_buffer_output[2] ),
    .A2(_2965_),
    .B1(_0627_),
    .Y(_2190_));
 sky130_fd_sc_hd__nand2_1 _5690_ (.A(_0352_),
    .B(_0416_),
    .Y(_2191_));
 sky130_fd_sc_hd__o21ai_1 _5691_ (.A1(_0960_),
    .A2(_0349_),
    .B1(_2191_),
    .Y(_2192_));
 sky130_fd_sc_hd__a221oi_1 _5692_ (.A1(_0948_),
    .A2(_0341_),
    .B1(_0344_),
    .B2(_0412_),
    .C1(_2192_),
    .Y(_2193_));
 sky130_fd_sc_hd__nand2_1 _5693_ (.A(_0370_),
    .B(_0400_),
    .Y(_2194_));
 sky130_fd_sc_hd__o21ai_1 _5694_ (.A1(_1466_),
    .A2(_0367_),
    .B1(_2194_),
    .Y(_2195_));
 sky130_fd_sc_hd__a221oi_1 _5695_ (.A1(_0642_),
    .A2(_0359_),
    .B1(_0362_),
    .B2(_0874_),
    .C1(_2195_),
    .Y(_2196_));
 sky130_fd_sc_hd__nand2_1 _5696_ (.A(_0387_),
    .B(_0436_),
    .Y(_2197_));
 sky130_fd_sc_hd__o21ai_1 _5697_ (.A1(_0965_),
    .A2(_0385_),
    .B1(_2197_),
    .Y(_2198_));
 sky130_fd_sc_hd__a221oi_1 _5698_ (.A1(_0655_),
    .A2(_0378_),
    .B1(_0429_),
    .B2(_0382_),
    .C1(_2198_),
    .Y(_2199_));
 sky130_fd_sc_hd__nand2_1 _5699_ (.A(_0405_),
    .B(_0447_),
    .Y(_2200_));
 sky130_fd_sc_hd__o21ai_1 _5700_ (.A1(_0647_),
    .A2(_0402_),
    .B1(_2200_),
    .Y(_2201_));
 sky130_fd_sc_hd__a221oi_1 _5701_ (.A1(_0461_),
    .A2(_0395_),
    .B1(_0398_),
    .B2(_0459_),
    .C1(_2201_),
    .Y(_2202_));
 sky130_fd_sc_hd__and4_1 _5702_ (.A(_2193_),
    .B(_2196_),
    .C(_2199_),
    .D(_2202_),
    .X(_2203_));
 sky130_fd_sc_hd__or2_1 _5703_ (.A(_0887_),
    .B(_0424_),
    .X(_2204_));
 sky130_fd_sc_hd__o21ai_1 _5704_ (.A1(_0955_),
    .A2(_0421_),
    .B1(_2204_),
    .Y(_2205_));
 sky130_fd_sc_hd__a221oi_1 _5705_ (.A1(_0664_),
    .A2(_0414_),
    .B1(_3244_),
    .B2(_0418_),
    .C1(_2205_),
    .Y(_2206_));
 sky130_fd_sc_hd__nand2_1 _5706_ (.A(_0457_),
    .B(\egd_top.BitStream_buffer.BS_buffer[71] ),
    .Y(_2207_));
 sky130_fd_sc_hd__nand2_1 _5707_ (.A(_0453_),
    .B(_3217_),
    .Y(_2208_));
 sky130_fd_sc_hd__or2_1 _5708_ (.A(_3257_),
    .B(_0449_),
    .X(_2209_));
 sky130_fd_sc_hd__o2111a_1 _5709_ (.A1(_0755_),
    .A2(_0464_),
    .B1(_2207_),
    .C1(_2208_),
    .D1(_2209_),
    .X(_2210_));
 sky130_fd_sc_hd__nand2_1 _5710_ (.A(_0431_),
    .B(_3237_),
    .Y(_2211_));
 sky130_fd_sc_hd__nand2_1 _5711_ (.A(_0442_),
    .B(_0751_),
    .Y(_2212_));
 sky130_fd_sc_hd__nand2_1 _5712_ (.A(_0434_),
    .B(_3210_),
    .Y(_2213_));
 sky130_fd_sc_hd__o2111a_1 _5713_ (.A1(_1297_),
    .A2(_0438_),
    .B1(_2211_),
    .C1(_2212_),
    .D1(_2213_),
    .X(_2214_));
 sky130_fd_sc_hd__nand2_1 _5714_ (.A(_0469_),
    .B(\egd_top.BitStream_buffer.BS_buffer[73] ),
    .Y(_2215_));
 sky130_fd_sc_hd__o21ai_1 _5715_ (.A1(_0833_),
    .A2(_0472_),
    .B1(_2215_),
    .Y(_2216_));
 sky130_fd_sc_hd__a221oi_1 _5716_ (.A1(_3252_),
    .A2(_0477_),
    .B1(_3268_),
    .B2(_2936_),
    .C1(_2216_),
    .Y(_2217_));
 sky130_fd_sc_hd__and4_1 _5717_ (.A(_2206_),
    .B(_2210_),
    .C(_2214_),
    .D(_2217_),
    .X(_2218_));
 sky130_fd_sc_hd__nand2_1 _5718_ (.A(_0560_),
    .B(_0498_),
    .Y(_2219_));
 sky130_fd_sc_hd__nand2_1 _5719_ (.A(_0564_),
    .B(\egd_top.BitStream_buffer.BS_buffer[17] ),
    .Y(_2220_));
 sky130_fd_sc_hd__or2_1 _5720_ (.A(_0492_),
    .B(_0570_),
    .X(_2221_));
 sky130_fd_sc_hd__o2111a_1 _5721_ (.A1(_0897_),
    .A2(_0557_),
    .B1(_2219_),
    .C1(_2220_),
    .D1(_2221_),
    .X(_2222_));
 sky130_fd_sc_hd__nand2_1 _5722_ (.A(_0577_),
    .B(_0505_),
    .Y(_2223_));
 sky130_fd_sc_hd__nand2_1 _5723_ (.A(_0581_),
    .B(_0509_),
    .Y(_2224_));
 sky130_fd_sc_hd__or2_1 _5724_ (.A(_1128_),
    .B(_0587_),
    .X(_2225_));
 sky130_fd_sc_hd__o2111a_1 _5725_ (.A1(_0520_),
    .A2(_0575_),
    .B1(_2223_),
    .C1(_2224_),
    .D1(_2225_),
    .X(_2226_));
 sky130_fd_sc_hd__or2_1 _5726_ (.A(_0685_),
    .B(_0598_),
    .X(_2227_));
 sky130_fd_sc_hd__o221a_1 _5727_ (.A1(_0602_),
    .A2(_0592_),
    .B1(_0688_),
    .B2(_0595_),
    .C1(_2227_),
    .X(_2228_));
 sky130_fd_sc_hd__nand2_1 _5728_ (.A(_0608_),
    .B(\egd_top.BitStream_buffer.BS_buffer[27] ),
    .Y(_2229_));
 sky130_fd_sc_hd__nand2_1 _5729_ (.A(_0605_),
    .B(_0527_),
    .Y(_2230_));
 sky130_fd_sc_hd__or2_1 _5730_ (.A(_0532_),
    .B(_0612_),
    .X(_2231_));
 sky130_fd_sc_hd__o2111a_1 _5731_ (.A1(_0699_),
    .A2(_0603_),
    .B1(_2229_),
    .C1(_2230_),
    .D1(_2231_),
    .X(_2232_));
 sky130_fd_sc_hd__and4_1 _5732_ (.A(_2222_),
    .B(_2226_),
    .C(_2228_),
    .D(_2232_),
    .X(_2233_));
 sky130_fd_sc_hd__nand2_1 _5733_ (.A(_0486_),
    .B(\egd_top.BitStream_buffer.BS_buffer[29] ),
    .Y(_2234_));
 sky130_fd_sc_hd__nand2_1 _5734_ (.A(_0489_),
    .B(_0537_),
    .Y(_2235_));
 sky130_fd_sc_hd__nand2_1 _5735_ (.A(_0496_),
    .B(\egd_top.BitStream_buffer.BS_buffer[32] ),
    .Y(_2236_));
 sky130_fd_sc_hd__o2111a_1 _5736_ (.A1(_0907_),
    .A2(_0494_),
    .B1(_2234_),
    .C1(_2235_),
    .D1(_2236_),
    .X(_2237_));
 sky130_fd_sc_hd__nand2_1 _5737_ (.A(_0513_),
    .B(_0364_),
    .Y(_2238_));
 sky130_fd_sc_hd__nand2_1 _5738_ (.A(_0503_),
    .B(_0365_),
    .Y(_2239_));
 sky130_fd_sc_hd__nand2_1 _5739_ (.A(_0901_),
    .B(_0337_),
    .Y(_2240_));
 sky130_fd_sc_hd__o2111a_1 _5740_ (.A1(_0633_),
    .A2(_0506_),
    .B1(_2238_),
    .C1(_2239_),
    .D1(_2240_),
    .X(_2241_));
 sky130_fd_sc_hd__nand2_1 _5741_ (.A(_0547_),
    .B(_0379_),
    .Y(_2242_));
 sky130_fd_sc_hd__o21ai_1 _5742_ (.A1(_0936_),
    .A2(_0545_),
    .B1(_2242_),
    .Y(_2243_));
 sky130_fd_sc_hd__a221oi_1 _5743_ (.A1(_0869_),
    .A2(_0538_),
    .B1(_0393_),
    .B2(_0541_),
    .C1(_2243_),
    .Y(_2244_));
 sky130_fd_sc_hd__o22a_1 _5744_ (.A1(_1276_),
    .A2(_0529_),
    .B1(_0348_),
    .B2(_0533_),
    .X(_2245_));
 sky130_fd_sc_hd__o221a_1 _5745_ (.A1(_1084_),
    .A2(_0522_),
    .B1(_0629_),
    .B2(_0525_),
    .C1(_2245_),
    .X(_2246_));
 sky130_fd_sc_hd__and4_1 _5746_ (.A(_2237_),
    .B(_2241_),
    .C(_2244_),
    .D(_2246_),
    .X(_2247_));
 sky130_fd_sc_hd__and4_1 _5747_ (.A(_2203_),
    .B(_2218_),
    .C(_2233_),
    .D(_2247_),
    .X(_2248_));
 sky130_fd_sc_hd__nand2_1 _5748_ (.A(_3061_),
    .B(_3169_),
    .Y(_2249_));
 sky130_fd_sc_hd__o21ai_1 _5749_ (.A1(_1035_),
    .A2(_3056_),
    .B1(_2249_),
    .Y(_2250_));
 sky130_fd_sc_hd__a221oi_2 _5750_ (.A1(_3070_),
    .A2(_3039_),
    .B1(_3075_),
    .B2(_3048_),
    .C1(_2250_),
    .Y(_2251_));
 sky130_fd_sc_hd__nand2_1 _5751_ (.A(_3099_),
    .B(_3157_),
    .Y(_2252_));
 sky130_fd_sc_hd__nand2_1 _5752_ (.A(_3093_),
    .B(_3164_),
    .Y(_2253_));
 sky130_fd_sc_hd__or2_1 _5753_ (.A(_2990_),
    .B(_3088_),
    .X(_2254_));
 sky130_fd_sc_hd__o2111a_1 _5754_ (.A1(_2983_),
    .A2(_3106_),
    .B1(_2252_),
    .C1(_2253_),
    .D1(_2254_),
    .X(_2255_));
 sky130_fd_sc_hd__nand2_1 _5755_ (.A(_3127_),
    .B(_0746_),
    .Y(_2256_));
 sky130_fd_sc_hd__o21ai_1 _5756_ (.A1(_2996_),
    .A2(_3123_),
    .B1(_2256_),
    .Y(_2257_));
 sky130_fd_sc_hd__a221oi_1 _5757_ (.A1(_3198_),
    .A2(_3113_),
    .B1(_3117_),
    .B2(_0744_),
    .C1(_2257_),
    .Y(_2258_));
 sky130_fd_sc_hd__nand2_1 _5758_ (.A(_3074_),
    .B(_3133_),
    .Y(_2259_));
 sky130_fd_sc_hd__o21ai_1 _5759_ (.A1(_3006_),
    .A2(_0729_),
    .B1(_2259_),
    .Y(_2260_));
 sky130_fd_sc_hd__a221oi_1 _5760_ (.A1(_3138_),
    .A2(_0726_),
    .B1(_3173_),
    .B2(_3081_),
    .C1(_2260_),
    .Y(_2261_));
 sky130_fd_sc_hd__and4_1 _5761_ (.A(_2251_),
    .B(_2255_),
    .C(_2258_),
    .D(_2261_),
    .X(_2262_));
 sky130_fd_sc_hd__nand2_1 _5762_ (.A(_3148_),
    .B(_0562_),
    .Y(_2263_));
 sky130_fd_sc_hd__o21ai_1 _5763_ (.A1(_0569_),
    .A2(_3145_),
    .B1(_2263_),
    .Y(_2264_));
 sky130_fd_sc_hd__a221oi_1 _5764_ (.A1(_0553_),
    .A2(_3137_),
    .B1(_0579_),
    .B2(_3141_),
    .C1(_2264_),
    .Y(_2265_));
 sky130_fd_sc_hd__nand2_1 _5765_ (.A(_3163_),
    .B(_0741_),
    .Y(_2266_));
 sky130_fd_sc_hd__nand2_1 _5766_ (.A(_3168_),
    .B(_3177_),
    .Y(_2267_));
 sky130_fd_sc_hd__nand2_1 _5767_ (.A(_2266_),
    .B(_2267_),
    .Y(_2268_));
 sky130_fd_sc_hd__a221oi_1 _5768_ (.A1(_3187_),
    .A2(_3156_),
    .B1(_0623_),
    .B2(_3160_),
    .C1(_2268_),
    .Y(_2269_));
 sky130_fd_sc_hd__nand2_1 _5769_ (.A(_3203_),
    .B(_0792_),
    .Y(_2270_));
 sky130_fd_sc_hd__o21ai_1 _5770_ (.A1(_0591_),
    .A2(_3200_),
    .B1(_2270_),
    .Y(_2271_));
 sky130_fd_sc_hd__a221oi_1 _5771_ (.A1(_1076_),
    .A2(_3194_),
    .B1(_3197_),
    .B2(_0566_),
    .C1(_2271_),
    .Y(_2272_));
 sky130_fd_sc_hd__nand2_1 _5772_ (.A(_3186_),
    .B(\egd_top.BitStream_buffer.BS_buffer[12] ),
    .Y(_2273_));
 sky130_fd_sc_hd__o21ai_1 _5773_ (.A1(_0574_),
    .A2(_3183_),
    .B1(_2273_),
    .Y(_2274_));
 sky130_fd_sc_hd__a221oi_1 _5774_ (.A1(_0585_),
    .A2(_3176_),
    .B1(_0583_),
    .B2(_3180_),
    .C1(_2274_),
    .Y(_2275_));
 sky130_fd_sc_hd__and4_1 _5775_ (.A(_2265_),
    .B(_2269_),
    .C(_2272_),
    .D(_2275_),
    .X(_2276_));
 sky130_fd_sc_hd__nand2_1 _5776_ (.A(_2262_),
    .B(_2276_),
    .Y(_2277_));
 sky130_fd_sc_hd__a22o_1 _5777_ (.A1(_3302_),
    .A2(_3215_),
    .B1(_3219_),
    .B2(_3288_),
    .X(_2278_));
 sky130_fd_sc_hd__a221oi_1 _5778_ (.A1(_3293_),
    .A2(_3224_),
    .B1(_3315_),
    .B2(_3226_),
    .C1(_2278_),
    .Y(_2279_));
 sky130_fd_sc_hd__nand2_1 _5779_ (.A(_3243_),
    .B(_3272_),
    .Y(_2280_));
 sky130_fd_sc_hd__o21ai_1 _5780_ (.A1(_1574_),
    .A2(_3240_),
    .B1(_2280_),
    .Y(_2281_));
 sky130_fd_sc_hd__a221oi_1 _5781_ (.A1(_3276_),
    .A2(_3233_),
    .B1(_3236_),
    .B2(_0837_),
    .C1(_2281_),
    .Y(_2282_));
 sky130_fd_sc_hd__nand2_1 _5782_ (.A(_3263_),
    .B(_3311_),
    .Y(_2283_));
 sky130_fd_sc_hd__o21ai_1 _5783_ (.A1(_3317_),
    .A2(_3260_),
    .B1(_2283_),
    .Y(_2284_));
 sky130_fd_sc_hd__a221oi_1 _5784_ (.A1(_0772_),
    .A2(_3251_),
    .B1(_3334_),
    .B2(_3255_),
    .C1(_2284_),
    .Y(_2285_));
 sky130_fd_sc_hd__nand2_1 _5785_ (.A(_3282_),
    .B(_3327_),
    .Y(_2286_));
 sky130_fd_sc_hd__o21ai_1 _5786_ (.A1(_1003_),
    .A2(_3279_),
    .B1(_2286_),
    .Y(_2287_));
 sky130_fd_sc_hd__a221oi_1 _5787_ (.A1(_0780_),
    .A2(_3271_),
    .B1(_3322_),
    .B2(_3275_),
    .C1(_2287_),
    .Y(_2288_));
 sky130_fd_sc_hd__and4_1 _5788_ (.A(_2279_),
    .B(_2282_),
    .C(_2285_),
    .D(_2288_),
    .X(_2289_));
 sky130_fd_sc_hd__nand2_1 _5789_ (.A(_3301_),
    .B(_3338_),
    .Y(_2290_));
 sky130_fd_sc_hd__o21ai_1 _5790_ (.A1(_0324_),
    .A2(_3299_),
    .B1(_2290_),
    .Y(_2291_));
 sky130_fd_sc_hd__a221oi_1 _5791_ (.A1(_3028_),
    .A2(_3295_),
    .B1(_3341_),
    .B2(_3292_),
    .C1(_2291_),
    .Y(_2292_));
 sky130_fd_sc_hd__nand2_1 _5792_ (.A(_3314_),
    .B(_3040_),
    .Y(_2293_));
 sky130_fd_sc_hd__nand2_1 _5793_ (.A(_3310_),
    .B(_3062_),
    .Y(_2294_));
 sky130_fd_sc_hd__or2_1 _5794_ (.A(_3049_),
    .B(_3319_),
    .X(_2295_));
 sky130_fd_sc_hd__o2111a_1 _5795_ (.A1(_0796_),
    .A2(_3308_),
    .B1(_2293_),
    .C1(_2294_),
    .D1(_2295_),
    .X(_2296_));
 sky130_fd_sc_hd__nand2_1 _5796_ (.A(_3333_),
    .B(_0716_),
    .Y(_2297_));
 sky130_fd_sc_hd__o21ai_1 _5797_ (.A1(_0713_),
    .A2(_3330_),
    .B1(_2297_),
    .Y(_2298_));
 sky130_fd_sc_hd__a221oi_1 _5798_ (.A1(_0714_),
    .A2(_3324_),
    .B1(_3326_),
    .B2(_3128_),
    .C1(_2298_),
    .Y(_2299_));
 sky130_fd_sc_hd__nand2_1 _5799_ (.A(_0329_),
    .B(_0722_),
    .Y(_2300_));
 sky130_fd_sc_hd__o21ai_1 _5800_ (.A1(_0721_),
    .A2(_0327_),
    .B1(_2300_),
    .Y(_2301_));
 sky130_fd_sc_hd__a221oi_1 _5801_ (.A1(_3118_),
    .A2(_3340_),
    .B1(_3066_),
    .B2(_0323_),
    .C1(_2301_),
    .Y(_2302_));
 sky130_fd_sc_hd__and4_1 _5802_ (.A(_2292_),
    .B(_2296_),
    .C(_2299_),
    .D(_2302_),
    .X(_2303_));
 sky130_fd_sc_hd__nand2_1 _5803_ (.A(_2289_),
    .B(_2303_),
    .Y(_2304_));
 sky130_fd_sc_hd__nor2_1 _5804_ (.A(_2277_),
    .B(_2304_),
    .Y(_2305_));
 sky130_fd_sc_hd__nand2_1 _5805_ (.A(_0621_),
    .B(\egd_top.BitStream_buffer.BS_buffer[13] ),
    .Y(_2306_));
 sky130_fd_sc_hd__nand3_1 _5806_ (.A(_2248_),
    .B(_2305_),
    .C(_2306_),
    .Y(_2307_));
 sky130_fd_sc_hd__nor2_1 _5807_ (.A(_3026_),
    .B(_2307_),
    .Y(_2308_));
 sky130_fd_sc_hd__nor2_1 _5808_ (.A(_2190_),
    .B(_2308_),
    .Y(_0284_));
 sky130_fd_sc_hd__o21ai_1 _5809_ (.A1(\egd_top.BitStream_buffer.BitStream_buffer_output[1] ),
    .A2(_2964_),
    .B1(_0627_),
    .Y(_2309_));
 sky130_fd_sc_hd__nand2_1 _5810_ (.A(_3243_),
    .B(_3283_),
    .Y(_2310_));
 sky130_fd_sc_hd__o21ai_1 _5811_ (.A1(_3277_),
    .A2(_3240_),
    .B1(_2310_),
    .Y(_2311_));
 sky130_fd_sc_hd__a221oi_1 _5812_ (.A1(_0837_),
    .A2(_3233_),
    .B1(_3236_),
    .B2(_3302_),
    .C1(_2311_),
    .Y(_2312_));
 sky130_fd_sc_hd__nand2_1 _5813_ (.A(_3223_),
    .B(_3315_),
    .Y(_2313_));
 sky130_fd_sc_hd__o21ai_1 _5814_ (.A1(_3317_),
    .A2(_1145_),
    .B1(_2313_),
    .Y(_2314_));
 sky130_fd_sc_hd__a221oi_1 _5815_ (.A1(_3288_),
    .A2(_3216_),
    .B1(_3293_),
    .B2(_3220_),
    .C1(_2314_),
    .Y(_2315_));
 sky130_fd_sc_hd__a22o_1 _5816_ (.A1(_0330_),
    .A2(_3281_),
    .B1(_1153_),
    .B2(_0785_),
    .X(_2316_));
 sky130_fd_sc_hd__a221oi_1 _5817_ (.A1(_3322_),
    .A2(_3271_),
    .B1(_3327_),
    .B2(_3275_),
    .C1(_2316_),
    .Y(_2317_));
 sky130_fd_sc_hd__nand2_1 _5818_ (.A(_3250_),
    .B(\egd_top.BitStream_buffer.BS_buffer[88] ),
    .Y(_2318_));
 sky130_fd_sc_hd__nand2_1 _5819_ (.A(_3262_),
    .B(_0772_),
    .Y(_2319_));
 sky130_fd_sc_hd__nand2_1 _5820_ (.A(_3255_),
    .B(_0780_),
    .Y(_2320_));
 sky130_fd_sc_hd__o2111a_1 _5821_ (.A1(_0771_),
    .A2(_3260_),
    .B1(_2318_),
    .C1(_2319_),
    .D1(_2320_),
    .X(_2321_));
 sky130_fd_sc_hd__and4_1 _5822_ (.A(_2312_),
    .B(_2315_),
    .C(_2317_),
    .D(_2321_),
    .X(_2322_));
 sky130_fd_sc_hd__nand2_1 _5823_ (.A(_3038_),
    .B(_3075_),
    .Y(_2323_));
 sky130_fd_sc_hd__nand2_1 _5824_ (.A(_3047_),
    .B(_3082_),
    .Y(_2324_));
 sky130_fd_sc_hd__nand2_1 _5825_ (.A(_3061_),
    .B(_3164_),
    .Y(_2325_));
 sky130_fd_sc_hd__o2111a_1 _5826_ (.A1(_2977_),
    .A2(_3056_),
    .B1(_2323_),
    .C1(_2324_),
    .D1(_2325_),
    .X(_2326_));
 sky130_fd_sc_hd__nand2_1 _5827_ (.A(_3092_),
    .B(_3153_),
    .Y(_2327_));
 sky130_fd_sc_hd__nand2_1 _5828_ (.A(_3099_),
    .B(\egd_top.BitStream_buffer.BS_buffer[116] ),
    .Y(_2328_));
 sky130_fd_sc_hd__or2_1 _5829_ (.A(_2986_),
    .B(_3105_),
    .X(_2329_));
 sky130_fd_sc_hd__o2111a_1 _5830_ (.A1(_2993_),
    .A2(_3089_),
    .B1(_2327_),
    .C1(_2328_),
    .D1(_2329_),
    .X(_2330_));
 sky130_fd_sc_hd__nand2_1 _5831_ (.A(_3126_),
    .B(_3191_),
    .Y(_2331_));
 sky130_fd_sc_hd__nand2_1 _5832_ (.A(_3112_),
    .B(_0744_),
    .Y(_2332_));
 sky130_fd_sc_hd__nand2_1 _5833_ (.A(_3116_),
    .B(_3149_),
    .Y(_2333_));
 sky130_fd_sc_hd__o2111a_1 _5834_ (.A1(_2999_),
    .A2(_3122_),
    .B1(_2331_),
    .C1(_2332_),
    .D1(_2333_),
    .X(_2334_));
 sky130_fd_sc_hd__nand2_1 _5835_ (.A(_3073_),
    .B(\egd_top.BitStream_buffer.BS_buffer[123] ),
    .Y(_2335_));
 sky130_fd_sc_hd__o21ai_1 _5836_ (.A1(_3009_),
    .A2(_0728_),
    .B1(_2335_),
    .Y(_2336_));
 sky130_fd_sc_hd__a221oi_1 _5837_ (.A1(_3173_),
    .A2(_3078_),
    .B1(_3177_),
    .B2(_3080_),
    .C1(_2336_),
    .Y(_2337_));
 sky130_fd_sc_hd__and4_1 _5838_ (.A(_2326_),
    .B(_2330_),
    .C(_2334_),
    .D(_2337_),
    .X(_2338_));
 sky130_fd_sc_hd__nand2_1 _5839_ (.A(_3332_),
    .B(_3100_),
    .Y(_2339_));
 sky130_fd_sc_hd__o21ai_1 _5840_ (.A1(_3085_),
    .A2(_3329_),
    .B1(_2339_),
    .Y(_2340_));
 sky130_fd_sc_hd__a221oi_1 _5841_ (.A1(_3128_),
    .A2(_3323_),
    .B1(_3325_),
    .B2(_0722_),
    .C1(_2340_),
    .Y(_2341_));
 sky130_fd_sc_hd__nand2_1 _5842_ (.A(_3313_),
    .B(_0708_),
    .Y(_2342_));
 sky130_fd_sc_hd__nand2_1 _5843_ (.A(_3309_),
    .B(_3094_),
    .Y(_2343_));
 sky130_fd_sc_hd__or2_1 _5844_ (.A(_0709_),
    .B(_3318_),
    .X(_2344_));
 sky130_fd_sc_hd__o2111a_1 _5845_ (.A1(_3102_),
    .A2(_3307_),
    .B1(_2342_),
    .C1(_2343_),
    .D1(_2344_),
    .X(_2345_));
 sky130_fd_sc_hd__nand2_1 _5846_ (.A(_3294_),
    .B(\egd_top.BitStream_buffer.BS_buffer[97] ),
    .Y(_2346_));
 sky130_fd_sc_hd__nand2_1 _5847_ (.A(_3300_),
    .B(\egd_top.BitStream_buffer.BS_buffer[95] ),
    .Y(_2347_));
 sky130_fd_sc_hd__or2_1 _5848_ (.A(_0784_),
    .B(_3298_),
    .X(_2348_));
 sky130_fd_sc_hd__nand2_1 _5849_ (.A(_3291_),
    .B(\egd_top.BitStream_buffer.BS_buffer[96] ),
    .Y(_2349_));
 sky130_fd_sc_hd__and4_1 _5850_ (.A(_2346_),
    .B(_2347_),
    .C(_2348_),
    .D(_2349_),
    .X(_2350_));
 sky130_fd_sc_hd__nand2_1 _5851_ (.A(_0328_),
    .B(_3109_),
    .Y(_2351_));
 sky130_fd_sc_hd__o21ai_1 _5852_ (.A1(_0804_),
    .A2(_0326_),
    .B1(_2351_),
    .Y(_2352_));
 sky130_fd_sc_hd__a221oi_1 _5853_ (.A1(_3066_),
    .A2(_3339_),
    .B1(_3070_),
    .B2(_0322_),
    .C1(_2352_),
    .Y(_2353_));
 sky130_fd_sc_hd__and4_1 _5854_ (.A(_2341_),
    .B(_2345_),
    .C(_2350_),
    .D(_2353_),
    .X(_2354_));
 sky130_fd_sc_hd__nand2_1 _5855_ (.A(_3202_),
    .B(_0930_),
    .Y(_2355_));
 sky130_fd_sc_hd__o21ai_1 _5856_ (.A1(_0597_),
    .A2(_3199_),
    .B1(_2355_),
    .Y(_2356_));
 sky130_fd_sc_hd__a221oi_1 _5857_ (.A1(_0566_),
    .A2(_3193_),
    .B1(_3196_),
    .B2(_0568_),
    .C1(_2356_),
    .Y(_2357_));
 sky130_fd_sc_hd__nand2_1 _5858_ (.A(_3162_),
    .B(_3187_),
    .Y(_2358_));
 sky130_fd_sc_hd__nand2_1 _5859_ (.A(_3159_),
    .B(_0792_),
    .Y(_2359_));
 sky130_fd_sc_hd__nand2_1 _5860_ (.A(_3167_),
    .B(\egd_top.BitStream_buffer.BS_buffer[126] ),
    .Y(_2360_));
 sky130_fd_sc_hd__nand2_1 _5861_ (.A(_3155_),
    .B(\egd_top.BitStream_buffer.BS_buffer[0] ),
    .Y(_2361_));
 sky130_fd_sc_hd__and4_1 _5862_ (.A(_2358_),
    .B(_2359_),
    .C(_2360_),
    .D(_2361_),
    .X(_2362_));
 sky130_fd_sc_hd__nand2_1 _5863_ (.A(_3147_),
    .B(_0553_),
    .Y(_2363_));
 sky130_fd_sc_hd__nand2_1 _5864_ (.A(_3140_),
    .B(_0585_),
    .Y(_2364_));
 sky130_fd_sc_hd__nand2_1 _5865_ (.A(_3136_),
    .B(_0579_),
    .Y(_2365_));
 sky130_fd_sc_hd__nand2_1 _5866_ (.A(_3144_),
    .B(_0562_),
    .Y(_2366_));
 sky130_fd_sc_hd__and4_1 _5867_ (.A(_2363_),
    .B(_2364_),
    .C(_2365_),
    .D(_2366_),
    .X(_2367_));
 sky130_fd_sc_hd__nand2_1 _5868_ (.A(_3185_),
    .B(\egd_top.BitStream_buffer.BS_buffer[13] ),
    .Y(_2368_));
 sky130_fd_sc_hd__o21ai_1 _5869_ (.A1(_0676_),
    .A2(_3183_),
    .B1(_2368_),
    .Y(_2369_));
 sky130_fd_sc_hd__a221oi_1 _5870_ (.A1(_0583_),
    .A2(_3176_),
    .B1(\egd_top.BitStream_buffer.BS_buffer[11] ),
    .B2(_3179_),
    .C1(_2369_),
    .Y(_2370_));
 sky130_fd_sc_hd__and4_1 _5871_ (.A(_2357_),
    .B(_2362_),
    .C(_2367_),
    .D(_2370_),
    .X(_2371_));
 sky130_fd_sc_hd__and4_1 _5872_ (.A(_2322_),
    .B(_2338_),
    .C(_2354_),
    .D(_2371_),
    .X(_2372_));
 sky130_fd_sc_hd__nand2_1 _5873_ (.A(_0353_),
    .B(_0443_),
    .Y(_2373_));
 sky130_fd_sc_hd__o21ai_1 _5874_ (.A1(_0437_),
    .A2(_0350_),
    .B1(_2373_),
    .Y(_2374_));
 sky130_fd_sc_hd__a221oi_1 _5875_ (.A1(_0412_),
    .A2(_0342_),
    .B1(_0345_),
    .B2(_0416_),
    .C1(_2374_),
    .Y(_2375_));
 sky130_fd_sc_hd__nand2_1 _5876_ (.A(_0388_),
    .B(_0454_),
    .Y(_2376_));
 sky130_fd_sc_hd__o21ai_1 _5877_ (.A1(_0462_),
    .A2(_0385_),
    .B1(_2376_),
    .Y(_2377_));
 sky130_fd_sc_hd__a221oi_1 _5878_ (.A1(_0429_),
    .A2(_0378_),
    .B1(_0436_),
    .B2(_0382_),
    .C1(_2377_),
    .Y(_2378_));
 sky130_fd_sc_hd__nand2_1 _5879_ (.A(_0371_),
    .B(_0407_),
    .Y(_2379_));
 sky130_fd_sc_hd__o21ai_1 _5880_ (.A1(_0401_),
    .A2(_0368_),
    .B1(_2379_),
    .Y(_2380_));
 sky130_fd_sc_hd__a221oi_1 _5881_ (.A1(_0874_),
    .A2(_0360_),
    .B1(_0363_),
    .B2(_0948_),
    .C1(_2380_),
    .Y(_2381_));
 sky130_fd_sc_hd__nand2_1 _5882_ (.A(_0406_),
    .B(_0467_),
    .Y(_2382_));
 sky130_fd_sc_hd__o21ai_1 _5883_ (.A1(_0887_),
    .A2(_0403_),
    .B1(_2382_),
    .Y(_2383_));
 sky130_fd_sc_hd__a221oi_1 _5884_ (.A1(_0459_),
    .A2(_0396_),
    .B1(_0399_),
    .B2(_0447_),
    .C1(_2383_),
    .Y(_2384_));
 sky130_fd_sc_hd__and4_1 _5885_ (.A(_2375_),
    .B(_2378_),
    .C(_2381_),
    .D(_2384_),
    .X(_2385_));
 sky130_fd_sc_hd__or2_1 _5886_ (.A(_0955_),
    .B(_0425_),
    .X(_2386_));
 sky130_fd_sc_hd__o21ai_1 _5887_ (.A1(_0474_),
    .A2(_0422_),
    .B1(_2386_),
    .Y(_2387_));
 sky130_fd_sc_hd__a221oi_1 _5888_ (.A1(_3244_),
    .A2(_0415_),
    .B1(_0751_),
    .B2(_0419_),
    .C1(_2387_),
    .Y(_2388_));
 sky130_fd_sc_hd__nand2_1 _5889_ (.A(_0442_),
    .B(_3230_),
    .Y(_2389_));
 sky130_fd_sc_hd__o21ai_1 _5890_ (.A1(_0829_),
    .A2(_0439_),
    .B1(_2389_),
    .Y(_2390_));
 sky130_fd_sc_hd__a221oi_1 _5891_ (.A1(_3210_),
    .A2(_0432_),
    .B1(_0435_),
    .B2(_3217_),
    .C1(_2390_),
    .Y(_2391_));
 sky130_fd_sc_hd__nand2_1 _5892_ (.A(_0453_),
    .B(_3221_),
    .Y(_2392_));
 sky130_fd_sc_hd__nand2_1 _5893_ (.A(_0458_),
    .B(_3256_),
    .Y(_2393_));
 sky130_fd_sc_hd__or2_1 _5894_ (.A(_1430_),
    .B(_0464_),
    .X(_2394_));
 sky130_fd_sc_hd__o2111a_1 _5895_ (.A1(_0759_),
    .A2(_0450_),
    .B1(_2392_),
    .C1(_2393_),
    .D1(_2394_),
    .X(_2395_));
 sky130_fd_sc_hd__nand2_1 _5896_ (.A(_0477_),
    .B(_3268_),
    .Y(_2396_));
 sky130_fd_sc_hd__o21ai_1 _5897_ (.A1(_1426_),
    .A2(_2935_),
    .B1(_2396_),
    .Y(_2397_));
 sky130_fd_sc_hd__a221oi_1 _5898_ (.A1(_3248_),
    .A2(_0470_),
    .B1(_3252_),
    .B2(_0473_),
    .C1(_2397_),
    .Y(_2398_));
 sky130_fd_sc_hd__and4_1 _5899_ (.A(_2388_),
    .B(_2391_),
    .C(_2395_),
    .D(_2398_),
    .X(_2399_));
 sky130_fd_sc_hd__nand2_1 _5900_ (.A(_2385_),
    .B(_2399_),
    .Y(_2400_));
 sky130_fd_sc_hd__nand2_1 _5901_ (.A(_0497_),
    .B(_0365_),
    .Y(_2401_));
 sky130_fd_sc_hd__o21ai_1 _5902_ (.A1(_0995_),
    .A2(_0495_),
    .B1(_2401_),
    .Y(_2402_));
 sky130_fd_sc_hd__a221oi_1 _5903_ (.A1(_0537_),
    .A2(_0487_),
    .B1(_0540_),
    .B2(_0490_),
    .C1(_2402_),
    .Y(_2403_));
 sky130_fd_sc_hd__nand2_1 _5904_ (.A(_0514_),
    .B(_0337_),
    .Y(_2404_));
 sky130_fd_sc_hd__o21ai_1 _5905_ (.A1(_1084_),
    .A2(_0512_),
    .B1(_2404_),
    .Y(_2405_));
 sky130_fd_sc_hd__a221oi_1 _5906_ (.A1(\egd_top.BitStream_buffer.BS_buffer[34] ),
    .A2(_0504_),
    .B1(_0364_),
    .B2(_0508_),
    .C1(_2405_),
    .Y(_2406_));
 sky130_fd_sc_hd__o22a_1 _5907_ (.A1(_0348_),
    .A2(_0530_),
    .B1(_0629_),
    .B2(_0534_),
    .X(_2407_));
 sky130_fd_sc_hd__o221a_1 _5908_ (.A1(_1276_),
    .A2(_0523_),
    .B1(_0861_),
    .B2(_0526_),
    .C1(_2407_),
    .X(_2408_));
 sky130_fd_sc_hd__nand2_1 _5909_ (.A(_0548_),
    .B(_0389_),
    .Y(_2409_));
 sky130_fd_sc_hd__o21ai_1 _5910_ (.A1(_0383_),
    .A2(_0546_),
    .B1(_2409_),
    .Y(_2410_));
 sky130_fd_sc_hd__a221oi_1 _5911_ (.A1(_0393_),
    .A2(_0539_),
    .B1(_0400_),
    .B2(_0542_),
    .C1(_2410_),
    .Y(_2411_));
 sky130_fd_sc_hd__and4_1 _5912_ (.A(_2403_),
    .B(_2406_),
    .C(_2408_),
    .D(_2411_),
    .X(_2412_));
 sky130_fd_sc_hd__nand2_1 _5913_ (.A(_0561_),
    .B(_0502_),
    .Y(_2413_));
 sky130_fd_sc_hd__nand2_1 _5914_ (.A(_0565_),
    .B(_0491_),
    .Y(_2414_));
 sky130_fd_sc_hd__or2_1 _5915_ (.A(_0986_),
    .B(_0557_),
    .X(_2415_));
 sky130_fd_sc_hd__o2111a_1 _5916_ (.A1(_0692_),
    .A2(_0571_),
    .B1(_2413_),
    .C1(_2414_),
    .D1(_2415_),
    .X(_2416_));
 sky130_fd_sc_hd__nand2_1 _5917_ (.A(_0578_),
    .B(_0515_),
    .Y(_2417_));
 sky130_fd_sc_hd__nand2_1 _5918_ (.A(_0582_),
    .B(_0519_),
    .Y(_2418_));
 sky130_fd_sc_hd__or2_1 _5919_ (.A(_0510_),
    .B(_0588_),
    .X(_2419_));
 sky130_fd_sc_hd__o2111a_1 _5920_ (.A1(_0528_),
    .A2(_0576_),
    .B1(_2417_),
    .C1(_2418_),
    .D1(_2419_),
    .X(_2420_));
 sky130_fd_sc_hd__or2_1 _5921_ (.A(_0602_),
    .B(_0595_),
    .X(_2421_));
 sky130_fd_sc_hd__o221a_1 _5922_ (.A1(_0685_),
    .A2(_0593_),
    .B1(_0922_),
    .B2(_0599_),
    .C1(_2421_),
    .X(_2422_));
 sky130_fd_sc_hd__nand2_1 _5923_ (.A(_0609_),
    .B(\egd_top.BitStream_buffer.BS_buffer[28] ),
    .Y(_2423_));
 sky130_fd_sc_hd__nand2_1 _5924_ (.A(_0606_),
    .B(_0531_),
    .Y(_2424_));
 sky130_fd_sc_hd__or2_1 _5925_ (.A(_0524_),
    .B(_0613_),
    .X(_2425_));
 sky130_fd_sc_hd__o2111a_1 _5926_ (.A1(_0543_),
    .A2(_0604_),
    .B1(_2423_),
    .C1(_2424_),
    .D1(_2425_),
    .X(_2426_));
 sky130_fd_sc_hd__and4_1 _5927_ (.A(_2416_),
    .B(_2420_),
    .C(_2422_),
    .D(_2426_),
    .X(_2427_));
 sky130_fd_sc_hd__nand2_1 _5928_ (.A(_2412_),
    .B(_2427_),
    .Y(_2428_));
 sky130_fd_sc_hd__nor2_1 _5929_ (.A(_2400_),
    .B(_2428_),
    .Y(_2429_));
 sky130_fd_sc_hd__nand2_1 _5930_ (.A(_0621_),
    .B(\egd_top.BitStream_buffer.BS_buffer[14] ),
    .Y(_2430_));
 sky130_fd_sc_hd__nand3_1 _5931_ (.A(_2372_),
    .B(_2429_),
    .C(_2430_),
    .Y(_2431_));
 sky130_fd_sc_hd__nor2_1 _5932_ (.A(_3026_),
    .B(_2431_),
    .Y(_2432_));
 sky130_fd_sc_hd__nor2_1 _5933_ (.A(_2309_),
    .B(_2432_),
    .Y(_0283_));
 sky130_fd_sc_hd__nand2_1 _5934_ (.A(_2972_),
    .B(_2967_),
    .Y(_2433_));
 sky130_fd_sc_hd__and3_1 _5935_ (.A(_2974_),
    .B(_2901_),
    .C(_2433_),
    .X(_2434_));
 sky130_fd_sc_hd__clkbuf_1 _5936_ (.A(_2434_),
    .X(_0282_));
 sky130_fd_sc_hd__nand2_1 _5937_ (.A(_2971_),
    .B(_2938_),
    .Y(_2435_));
 sky130_fd_sc_hd__and3_1 _5938_ (.A(_2972_),
    .B(_2901_),
    .C(_2435_),
    .X(_2436_));
 sky130_fd_sc_hd__clkbuf_1 _5939_ (.A(_2436_),
    .X(_0281_));
 sky130_fd_sc_hd__inv_2 _5940_ (.A(_2970_),
    .Y(_2437_));
 sky130_fd_sc_hd__nand2_1 _5941_ (.A(_2437_),
    .B(_2939_),
    .Y(_2438_));
 sky130_fd_sc_hd__and3_1 _5942_ (.A(_2438_),
    .B(_2901_),
    .C(_2971_),
    .X(_2439_));
 sky130_fd_sc_hd__clkbuf_1 _5943_ (.A(_2439_),
    .X(_0280_));
 sky130_fd_sc_hd__or2_1 _5944_ (.A(_2944_),
    .B(_2437_),
    .X(_2440_));
 sky130_fd_sc_hd__clkbuf_2 _5945_ (.A(_2440_),
    .X(_2441_));
 sky130_fd_sc_hd__buf_2 _5946_ (.A(_2441_),
    .X(_2442_));
 sky130_fd_sc_hd__clkbuf_4 _5947_ (.A(_2441_),
    .X(_2443_));
 sky130_fd_sc_hd__nand2_1 _5948_ (.A(_2443_),
    .B(_1602_),
    .Y(_2444_));
 sky130_fd_sc_hd__o211a_1 _5949_ (.A1(_2966_),
    .A2(_2442_),
    .B1(_3002_),
    .C1(_2444_),
    .X(_0279_));
 sky130_fd_sc_hd__nand2_1 _5950_ (.A(_2443_),
    .B(_0594_),
    .Y(_2445_));
 sky130_fd_sc_hd__o211a_1 _5951_ (.A1(_2979_),
    .A2(_2442_),
    .B1(_3002_),
    .C1(_2445_),
    .X(_0278_));
 sky130_fd_sc_hd__buf_2 _5952_ (.A(_2901_),
    .X(_2446_));
 sky130_fd_sc_hd__nand2_1 _5953_ (.A(_2443_),
    .B(_0591_),
    .Y(_2447_));
 sky130_fd_sc_hd__o211a_1 _5954_ (.A1(_2982_),
    .A2(_2442_),
    .B1(_2446_),
    .C1(_2447_),
    .X(_0277_));
 sky130_fd_sc_hd__nand2_1 _5955_ (.A(_2443_),
    .B(_0597_),
    .Y(_2448_));
 sky130_fd_sc_hd__o211a_1 _5956_ (.A1(_2985_),
    .A2(_2442_),
    .B1(_2446_),
    .C1(_2448_),
    .X(_0276_));
 sky130_fd_sc_hd__clkbuf_4 _5957_ (.A(_2441_),
    .X(_2449_));
 sky130_fd_sc_hd__nand2_1 _5958_ (.A(_2449_),
    .B(_0682_),
    .Y(_2450_));
 sky130_fd_sc_hd__o211a_1 _5959_ (.A1(_2988_),
    .A2(_2442_),
    .B1(_2446_),
    .C1(_2450_),
    .X(_0275_));
 sky130_fd_sc_hd__nand2_1 _5960_ (.A(_2449_),
    .B(_0569_),
    .Y(_2451_));
 sky130_fd_sc_hd__o211a_1 _5961_ (.A1(_2992_),
    .A2(_2442_),
    .B1(_2446_),
    .C1(_2451_),
    .X(_0274_));
 sky130_fd_sc_hd__nand2_1 _5962_ (.A(_2449_),
    .B(_0673_),
    .Y(_2452_));
 sky130_fd_sc_hd__o211a_1 _5963_ (.A1(_2995_),
    .A2(_2442_),
    .B1(_2446_),
    .C1(_2452_),
    .X(_0273_));
 sky130_fd_sc_hd__nand2_1 _5964_ (.A(_2449_),
    .B(_0554_),
    .Y(_2453_));
 sky130_fd_sc_hd__o211a_1 _5965_ (.A1(_2998_),
    .A2(_2442_),
    .B1(_2446_),
    .C1(_2453_),
    .X(_0272_));
 sky130_fd_sc_hd__nand2_1 _5966_ (.A(_2449_),
    .B(_0670_),
    .Y(_2454_));
 sky130_fd_sc_hd__o211a_1 _5967_ (.A1(_3001_),
    .A2(_2442_),
    .B1(_2446_),
    .C1(_2454_),
    .X(_0271_));
 sky130_fd_sc_hd__nand2_1 _5968_ (.A(_2449_),
    .B(_0586_),
    .Y(_2455_));
 sky130_fd_sc_hd__o211a_1 _5969_ (.A1(_3005_),
    .A2(_2442_),
    .B1(_2446_),
    .C1(_2455_),
    .X(_0270_));
 sky130_fd_sc_hd__nand2_1 _5970_ (.A(_2449_),
    .B(_0679_),
    .Y(_2456_));
 sky130_fd_sc_hd__o211a_1 _5971_ (.A1(_3008_),
    .A2(_2443_),
    .B1(_2446_),
    .C1(_2456_),
    .X(_0269_));
 sky130_fd_sc_hd__nand2_1 _5972_ (.A(_2449_),
    .B(_0574_),
    .Y(_2457_));
 sky130_fd_sc_hd__o211a_1 _5973_ (.A1(_3011_),
    .A2(_2443_),
    .B1(_2446_),
    .C1(_2457_),
    .X(_0268_));
 sky130_fd_sc_hd__buf_2 _5974_ (.A(_2901_),
    .X(_2458_));
 sky130_fd_sc_hd__nand2_1 _5975_ (.A(_2449_),
    .B(_0676_),
    .Y(_2459_));
 sky130_fd_sc_hd__o211a_1 _5976_ (.A1(_3014_),
    .A2(_2443_),
    .B1(_2458_),
    .C1(_2459_),
    .X(_0267_));
 sky130_fd_sc_hd__nand2_1 _5977_ (.A(_2449_),
    .B(_0611_),
    .Y(_2460_));
 sky130_fd_sc_hd__o211a_1 _5978_ (.A1(_3017_),
    .A2(_2443_),
    .B1(_2458_),
    .C1(_2460_),
    .X(_0266_));
 sky130_fd_sc_hd__nand2_1 _5979_ (.A(_2441_),
    .B(_0688_),
    .Y(_2461_));
 sky130_fd_sc_hd__o211a_1 _5980_ (.A1(_3020_),
    .A2(_2443_),
    .B1(_2458_),
    .C1(_2461_),
    .X(_0265_));
 sky130_fd_sc_hd__nand2_1 _5981_ (.A(_2441_),
    .B(_0602_),
    .Y(_2462_));
 sky130_fd_sc_hd__o211a_1 _5982_ (.A1(_3023_),
    .A2(_2443_),
    .B1(_2458_),
    .C1(_2462_),
    .X(_0264_));
 sky130_fd_sc_hd__or3_1 _5983_ (.A(\egd_top.BitStream_buffer.buffer_index[6] ),
    .B(\egd_top.BitStream_buffer.buffer_index[5] ),
    .C(_2971_),
    .X(_2463_));
 sky130_fd_sc_hd__clkbuf_2 _5984_ (.A(_2463_),
    .X(_2464_));
 sky130_fd_sc_hd__buf_2 _5985_ (.A(_2464_),
    .X(_2465_));
 sky130_fd_sc_hd__buf_2 _5986_ (.A(_2464_),
    .X(_2466_));
 sky130_fd_sc_hd__nand2_1 _5987_ (.A(_2466_),
    .B(_0685_),
    .Y(_2467_));
 sky130_fd_sc_hd__o211a_1 _5988_ (.A1(_2966_),
    .A2(_2465_),
    .B1(_2458_),
    .C1(_2467_),
    .X(_0263_));
 sky130_fd_sc_hd__nand2_1 _5989_ (.A(_2466_),
    .B(_0922_),
    .Y(_2468_));
 sky130_fd_sc_hd__o211a_1 _5990_ (.A1(_2979_),
    .A2(_2465_),
    .B1(_2458_),
    .C1(_2468_),
    .X(_0262_));
 sky130_fd_sc_hd__nand2_1 _5991_ (.A(_2466_),
    .B(_0492_),
    .Y(_2469_));
 sky130_fd_sc_hd__o211a_1 _5992_ (.A1(_2982_),
    .A2(_2465_),
    .B1(_2458_),
    .C1(_2469_),
    .X(_0261_));
 sky130_fd_sc_hd__nand2_1 _5993_ (.A(_2466_),
    .B(_0692_),
    .Y(_2470_));
 sky130_fd_sc_hd__o211a_1 _5994_ (.A1(_2985_),
    .A2(_2465_),
    .B1(_2458_),
    .C1(_2470_),
    .X(_0260_));
 sky130_fd_sc_hd__buf_2 _5995_ (.A(_2464_),
    .X(_2471_));
 sky130_fd_sc_hd__nand2_1 _5996_ (.A(_2471_),
    .B(_0897_),
    .Y(_2472_));
 sky130_fd_sc_hd__o211a_1 _5997_ (.A1(_2988_),
    .A2(_2465_),
    .B1(_2458_),
    .C1(_2472_),
    .X(_0259_));
 sky130_fd_sc_hd__nand2_1 _5998_ (.A(_2471_),
    .B(_0986_),
    .Y(_2473_));
 sky130_fd_sc_hd__o211a_1 _5999_ (.A1(_2992_),
    .A2(_2465_),
    .B1(_2458_),
    .C1(_2473_),
    .X(_0258_));
 sky130_fd_sc_hd__buf_2 _6000_ (.A(_2901_),
    .X(_2474_));
 sky130_fd_sc_hd__nand2_1 _6001_ (.A(_2471_),
    .B(_1128_),
    .Y(_2475_));
 sky130_fd_sc_hd__o211a_1 _6002_ (.A1(_2995_),
    .A2(_2465_),
    .B1(_2474_),
    .C1(_2475_),
    .X(_0257_));
 sky130_fd_sc_hd__nand2_1 _6003_ (.A(_2471_),
    .B(_0510_),
    .Y(_2476_));
 sky130_fd_sc_hd__o211a_1 _6004_ (.A1(_2998_),
    .A2(_2465_),
    .B1(_2474_),
    .C1(_2476_),
    .X(_0256_));
 sky130_fd_sc_hd__nand2_1 _6005_ (.A(_2471_),
    .B(_0520_),
    .Y(_2477_));
 sky130_fd_sc_hd__o211a_1 _6006_ (.A1(_3001_),
    .A2(_2465_),
    .B1(_2474_),
    .C1(_2477_),
    .X(_0255_));
 sky130_fd_sc_hd__nand2_1 _6007_ (.A(_2471_),
    .B(_0528_),
    .Y(_2478_));
 sky130_fd_sc_hd__o211a_1 _6008_ (.A1(_3005_),
    .A2(_2465_),
    .B1(_2474_),
    .C1(_2478_),
    .X(_0254_));
 sky130_fd_sc_hd__nand2_1 _6009_ (.A(_2471_),
    .B(_0532_),
    .Y(_2479_));
 sky130_fd_sc_hd__o211a_1 _6010_ (.A1(_3008_),
    .A2(_2466_),
    .B1(_2474_),
    .C1(_2479_),
    .X(_0253_));
 sky130_fd_sc_hd__nand2_1 _6011_ (.A(_2471_),
    .B(_0524_),
    .Y(_2480_));
 sky130_fd_sc_hd__o211a_1 _6012_ (.A1(_3011_),
    .A2(_2466_),
    .B1(_2474_),
    .C1(_2480_),
    .X(_0252_));
 sky130_fd_sc_hd__nand2_1 _6013_ (.A(_2471_),
    .B(_0699_),
    .Y(_2481_));
 sky130_fd_sc_hd__o211a_1 _6014_ (.A1(_3014_),
    .A2(_2466_),
    .B1(_2474_),
    .C1(_2481_),
    .X(_0251_));
 sky130_fd_sc_hd__nand2_1 _6015_ (.A(_2471_),
    .B(_0543_),
    .Y(_2482_));
 sky130_fd_sc_hd__o211a_1 _6016_ (.A1(_3017_),
    .A2(_2466_),
    .B1(_2474_),
    .C1(_2482_),
    .X(_0250_));
 sky130_fd_sc_hd__nand2_1 _6017_ (.A(_2464_),
    .B(_0702_),
    .Y(_2483_));
 sky130_fd_sc_hd__o211a_1 _6018_ (.A1(_3020_),
    .A2(_2466_),
    .B1(_2474_),
    .C1(_2483_),
    .X(_0249_));
 sky130_fd_sc_hd__nand2_1 _6019_ (.A(_2464_),
    .B(_0907_),
    .Y(_2484_));
 sky130_fd_sc_hd__o211a_1 _6020_ (.A1(_3023_),
    .A2(_2466_),
    .B1(_2474_),
    .C1(_2484_),
    .X(_0248_));
 sky130_fd_sc_hd__or4_1 _6021_ (.A(\egd_top.BitStream_buffer.buffer_index[6] ),
    .B(_2938_),
    .C(\egd_top.BitStream_buffer.buffer_index[4] ),
    .D(_2437_),
    .X(_2485_));
 sky130_fd_sc_hd__clkbuf_2 _6022_ (.A(_2485_),
    .X(_2486_));
 sky130_fd_sc_hd__buf_2 _6023_ (.A(_2486_),
    .X(_2487_));
 sky130_fd_sc_hd__buf_2 _6024_ (.A(_2904_),
    .X(_2488_));
 sky130_fd_sc_hd__buf_2 _6025_ (.A(_2486_),
    .X(_2489_));
 sky130_fd_sc_hd__nand2_1 _6026_ (.A(_2489_),
    .B(_0995_),
    .Y(_2490_));
 sky130_fd_sc_hd__o211a_1 _6027_ (.A1(_2966_),
    .A2(_2487_),
    .B1(_2488_),
    .C1(_2490_),
    .X(_0247_));
 sky130_fd_sc_hd__nand2_1 _6028_ (.A(_2489_),
    .B(_0366_),
    .Y(_2491_));
 sky130_fd_sc_hd__o211a_1 _6029_ (.A1(_2979_),
    .A2(_2487_),
    .B1(_2488_),
    .C1(_2491_),
    .X(_0246_));
 sky130_fd_sc_hd__nand2_1 _6030_ (.A(_2489_),
    .B(_0633_),
    .Y(_2492_));
 sky130_fd_sc_hd__o211a_1 _6031_ (.A1(_2982_),
    .A2(_2487_),
    .B1(_2488_),
    .C1(_2492_),
    .X(_0245_));
 sky130_fd_sc_hd__nand2_1 _6032_ (.A(_2489_),
    .B(_0865_),
    .Y(_2493_));
 sky130_fd_sc_hd__o211a_1 _6033_ (.A1(_2985_),
    .A2(_2487_),
    .B1(_2488_),
    .C1(_2493_),
    .X(_0244_));
 sky130_fd_sc_hd__buf_2 _6034_ (.A(_2486_),
    .X(_2494_));
 sky130_fd_sc_hd__nand2_1 _6035_ (.A(_2494_),
    .B(_0940_),
    .Y(_2495_));
 sky130_fd_sc_hd__o211a_1 _6036_ (.A1(_2988_),
    .A2(_2487_),
    .B1(_2488_),
    .C1(_2495_),
    .X(_0243_));
 sky130_fd_sc_hd__nand2_1 _6037_ (.A(_2494_),
    .B(_1084_),
    .Y(_2496_));
 sky130_fd_sc_hd__o211a_1 _6038_ (.A1(_2992_),
    .A2(_2487_),
    .B1(_2488_),
    .C1(_2496_),
    .X(_0242_));
 sky130_fd_sc_hd__nand2_1 _6039_ (.A(_2494_),
    .B(_1276_),
    .Y(_2497_));
 sky130_fd_sc_hd__o211a_1 _6040_ (.A1(_2995_),
    .A2(_2487_),
    .B1(_2488_),
    .C1(_2497_),
    .X(_0241_));
 sky130_fd_sc_hd__nand2_1 _6041_ (.A(_2494_),
    .B(_0348_),
    .Y(_2498_));
 sky130_fd_sc_hd__o211a_1 _6042_ (.A1(_2998_),
    .A2(_2487_),
    .B1(_2488_),
    .C1(_2498_),
    .X(_0240_));
 sky130_fd_sc_hd__nand2_1 _6043_ (.A(_2494_),
    .B(_0629_),
    .Y(_2499_));
 sky130_fd_sc_hd__o211a_1 _6044_ (.A1(_3001_),
    .A2(_2487_),
    .B1(_2488_),
    .C1(_2499_),
    .X(_0239_));
 sky130_fd_sc_hd__nand2_1 _6045_ (.A(_2494_),
    .B(_0861_),
    .Y(_2500_));
 sky130_fd_sc_hd__o211a_1 _6046_ (.A1(_3005_),
    .A2(_2487_),
    .B1(_2488_),
    .C1(_2500_),
    .X(_0238_));
 sky130_fd_sc_hd__buf_2 _6047_ (.A(_2904_),
    .X(_2501_));
 sky130_fd_sc_hd__nand2_1 _6048_ (.A(_2494_),
    .B(_0936_),
    .Y(_2502_));
 sky130_fd_sc_hd__o211a_1 _6049_ (.A1(_3008_),
    .A2(_2489_),
    .B1(_2501_),
    .C1(_2502_),
    .X(_0237_));
 sky130_fd_sc_hd__nand2_1 _6050_ (.A(_2494_),
    .B(_0383_),
    .Y(_2503_));
 sky130_fd_sc_hd__o211a_1 _6051_ (.A1(_3011_),
    .A2(_2489_),
    .B1(_2501_),
    .C1(_2503_),
    .X(_0236_));
 sky130_fd_sc_hd__nand2_1 _6052_ (.A(_2494_),
    .B(_0637_),
    .Y(_2504_));
 sky130_fd_sc_hd__o211a_1 _6053_ (.A1(_3014_),
    .A2(_2489_),
    .B1(_2501_),
    .C1(_2504_),
    .X(_0235_));
 sky130_fd_sc_hd__nand2_1 _6054_ (.A(_2494_),
    .B(_0870_),
    .Y(_2505_));
 sky130_fd_sc_hd__o211a_1 _6055_ (.A1(_3017_),
    .A2(_2489_),
    .B1(_2501_),
    .C1(_2505_),
    .X(_0234_));
 sky130_fd_sc_hd__nand2_1 _6056_ (.A(_2486_),
    .B(_1466_),
    .Y(_2506_));
 sky130_fd_sc_hd__o211a_1 _6057_ (.A1(_3020_),
    .A2(_2489_),
    .B1(_2501_),
    .C1(_2506_),
    .X(_0233_));
 sky130_fd_sc_hd__nand2_1 _6058_ (.A(_2486_),
    .B(_0401_),
    .Y(_2507_));
 sky130_fd_sc_hd__o211a_1 _6059_ (.A1(_3023_),
    .A2(_2489_),
    .B1(_2501_),
    .C1(_2507_),
    .X(_0232_));
 sky130_fd_sc_hd__nor2_1 _6060_ (.A(\egd_top.BitStream_buffer.buffer_index[6] ),
    .B(_2972_),
    .Y(_2508_));
 sky130_fd_sc_hd__clkinv_2 _6061_ (.A(_2508_),
    .Y(_2509_));
 sky130_fd_sc_hd__buf_2 _6062_ (.A(_2509_),
    .X(_2510_));
 sky130_fd_sc_hd__buf_2 _6063_ (.A(_2509_),
    .X(_2511_));
 sky130_fd_sc_hd__nand2_1 _6064_ (.A(_2511_),
    .B(_0423_),
    .Y(_2512_));
 sky130_fd_sc_hd__o211a_1 _6065_ (.A1(_2966_),
    .A2(_2510_),
    .B1(_2501_),
    .C1(_2512_),
    .X(_0231_));
 sky130_fd_sc_hd__nand2_1 _6066_ (.A(_2511_),
    .B(_0420_),
    .Y(_2513_));
 sky130_fd_sc_hd__o211a_1 _6067_ (.A1(_2979_),
    .A2(_2510_),
    .B1(_2501_),
    .C1(_2513_),
    .X(_0230_));
 sky130_fd_sc_hd__nand2_1 _6068_ (.A(_2511_),
    .B(_0659_),
    .Y(_2514_));
 sky130_fd_sc_hd__o211a_1 _6069_ (.A1(_2982_),
    .A2(_2510_),
    .B1(_2501_),
    .C1(_2514_),
    .X(_0229_));
 sky130_fd_sc_hd__nand2_1 _6070_ (.A(_2511_),
    .B(_0879_),
    .Y(_2515_));
 sky130_fd_sc_hd__o211a_1 _6071_ (.A1(_2985_),
    .A2(_2510_),
    .B1(_2501_),
    .C1(_2515_),
    .X(_0228_));
 sky130_fd_sc_hd__buf_2 _6072_ (.A(_2904_),
    .X(_2516_));
 sky130_fd_sc_hd__buf_2 _6073_ (.A(_2509_),
    .X(_2517_));
 sky130_fd_sc_hd__nand2_1 _6074_ (.A(_2517_),
    .B(_0960_),
    .Y(_2518_));
 sky130_fd_sc_hd__o211a_1 _6075_ (.A1(_2988_),
    .A2(_2510_),
    .B1(_2516_),
    .C1(_2518_),
    .X(_0227_));
 sky130_fd_sc_hd__nand2_1 _6076_ (.A(_2517_),
    .B(_0437_),
    .Y(_2519_));
 sky130_fd_sc_hd__o211a_1 _6077_ (.A1(_2992_),
    .A2(_2510_),
    .B1(_2516_),
    .C1(_2519_),
    .X(_0226_));
 sky130_fd_sc_hd__nand2_1 _6078_ (.A(_2517_),
    .B(_0653_),
    .Y(_2520_));
 sky130_fd_sc_hd__o211a_1 _6079_ (.A1(_2995_),
    .A2(_2510_),
    .B1(_2516_),
    .C1(_2520_),
    .X(_0225_));
 sky130_fd_sc_hd__nand2_1 _6080_ (.A(_2517_),
    .B(_0883_),
    .Y(_2521_));
 sky130_fd_sc_hd__o211a_1 _6081_ (.A1(_2998_),
    .A2(_2510_),
    .B1(_2516_),
    .C1(_2521_),
    .X(_0224_));
 sky130_fd_sc_hd__nand2_1 _6082_ (.A(_2517_),
    .B(_0965_),
    .Y(_2522_));
 sky130_fd_sc_hd__o211a_1 _6083_ (.A1(_3001_),
    .A2(_2510_),
    .B1(_2516_),
    .C1(_2522_),
    .X(_0223_));
 sky130_fd_sc_hd__nand2_1 _6084_ (.A(_2517_),
    .B(_0462_),
    .Y(_2523_));
 sky130_fd_sc_hd__o211a_1 _6085_ (.A1(_3005_),
    .A2(_2510_),
    .B1(_2516_),
    .C1(_2523_),
    .X(_0222_));
 sky130_fd_sc_hd__nand2_1 _6086_ (.A(_2517_),
    .B(_0650_),
    .Y(_2524_));
 sky130_fd_sc_hd__o211a_1 _6087_ (.A1(_3008_),
    .A2(_2511_),
    .B1(_2516_),
    .C1(_2524_),
    .X(_0221_));
 sky130_fd_sc_hd__nand2_1 _6088_ (.A(_2517_),
    .B(_0448_),
    .Y(_2525_));
 sky130_fd_sc_hd__o211a_1 _6089_ (.A1(_3011_),
    .A2(_2511_),
    .B1(_2516_),
    .C1(_2525_),
    .X(_0220_));
 sky130_fd_sc_hd__nand2_1 _6090_ (.A(_2517_),
    .B(_0647_),
    .Y(_2526_));
 sky130_fd_sc_hd__o211a_1 _6091_ (.A1(_3014_),
    .A2(_2511_),
    .B1(_2516_),
    .C1(_2526_),
    .X(_0219_));
 sky130_fd_sc_hd__nand2_1 _6092_ (.A(_2517_),
    .B(_0887_),
    .Y(_2527_));
 sky130_fd_sc_hd__o211a_1 _6093_ (.A1(_3017_),
    .A2(_2511_),
    .B1(_2516_),
    .C1(_2527_),
    .X(_0218_));
 sky130_fd_sc_hd__buf_2 _6094_ (.A(_2904_),
    .X(_2528_));
 sky130_fd_sc_hd__nand2_1 _6095_ (.A(_2509_),
    .B(_0955_),
    .Y(_2529_));
 sky130_fd_sc_hd__o211a_1 _6096_ (.A1(_3020_),
    .A2(_2511_),
    .B1(_2528_),
    .C1(_2529_),
    .X(_0217_));
 sky130_fd_sc_hd__nand2_1 _6097_ (.A(_2509_),
    .B(_0474_),
    .Y(_2530_));
 sky130_fd_sc_hd__o211a_1 _6098_ (.A1(_3023_),
    .A2(_2511_),
    .B1(_2528_),
    .C1(_2530_),
    .X(_0216_));
 sky130_fd_sc_hd__nand2_2 _6099_ (.A(_2970_),
    .B(_2940_),
    .Y(_2531_));
 sky130_fd_sc_hd__buf_2 _6100_ (.A(_2531_),
    .X(_2532_));
 sky130_fd_sc_hd__buf_2 _6101_ (.A(_2531_),
    .X(_2533_));
 sky130_fd_sc_hd__nand2_1 _6102_ (.A(_2533_),
    .B(_0663_),
    .Y(_2534_));
 sky130_fd_sc_hd__o211a_1 _6103_ (.A1(_2966_),
    .A2(_2532_),
    .B1(_2528_),
    .C1(_2534_),
    .X(_0215_));
 sky130_fd_sc_hd__nand2_1 _6104_ (.A(_2533_),
    .B(_3238_),
    .Y(_2535_));
 sky130_fd_sc_hd__o211a_1 _6105_ (.A1(_2979_),
    .A2(_2532_),
    .B1(_2528_),
    .C1(_2535_),
    .X(_0214_));
 sky130_fd_sc_hd__nand2_1 _6106_ (.A(_2533_),
    .B(_1297_),
    .Y(_2536_));
 sky130_fd_sc_hd__o211a_1 _6107_ (.A1(_2982_),
    .A2(_2532_),
    .B1(_2528_),
    .C1(_2536_),
    .X(_0213_));
 sky130_fd_sc_hd__nand2_1 _6108_ (.A(_2533_),
    .B(_0829_),
    .Y(_2537_));
 sky130_fd_sc_hd__o211a_1 _6109_ (.A1(_2985_),
    .A2(_2532_),
    .B1(_2528_),
    .C1(_2537_),
    .X(_0212_));
 sky130_fd_sc_hd__buf_2 _6110_ (.A(_2531_),
    .X(_2538_));
 sky130_fd_sc_hd__nand2_1 _6111_ (.A(_2538_),
    .B(_1043_),
    .Y(_2539_));
 sky130_fd_sc_hd__o211a_1 _6112_ (.A1(_2988_),
    .A2(_2532_),
    .B1(_2528_),
    .C1(_2539_),
    .X(_0211_));
 sky130_fd_sc_hd__nand2_1 _6113_ (.A(_2538_),
    .B(_1360_),
    .Y(_2540_));
 sky130_fd_sc_hd__o211a_1 _6114_ (.A1(_2992_),
    .A2(_2532_),
    .B1(_2528_),
    .C1(_2540_),
    .X(_0210_));
 sky130_fd_sc_hd__nand2_1 _6115_ (.A(_2538_),
    .B(_0755_),
    .Y(_2541_));
 sky130_fd_sc_hd__o211a_1 _6116_ (.A1(_2995_),
    .A2(_2532_),
    .B1(_2528_),
    .C1(_2541_),
    .X(_0209_));
 sky130_fd_sc_hd__nand2_1 _6117_ (.A(_2538_),
    .B(_1430_),
    .Y(_2542_));
 sky130_fd_sc_hd__o211a_1 _6118_ (.A1(_2998_),
    .A2(_2532_),
    .B1(_2528_),
    .C1(_2542_),
    .X(_0208_));
 sky130_fd_sc_hd__buf_2 _6119_ (.A(_2904_),
    .X(_2543_));
 sky130_fd_sc_hd__nand2_1 _6120_ (.A(_2538_),
    .B(_3257_),
    .Y(_2544_));
 sky130_fd_sc_hd__o211a_1 _6121_ (.A1(_3001_),
    .A2(_2532_),
    .B1(_2543_),
    .C1(_2544_),
    .X(_0207_));
 sky130_fd_sc_hd__nand2_1 _6122_ (.A(_2538_),
    .B(_0759_),
    .Y(_2545_));
 sky130_fd_sc_hd__o211a_1 _6123_ (.A1(_3005_),
    .A2(_2532_),
    .B1(_2543_),
    .C1(_2545_),
    .X(_0206_));
 sky130_fd_sc_hd__nand2_1 _6124_ (.A(_2538_),
    .B(_0833_),
    .Y(_2546_));
 sky130_fd_sc_hd__o211a_1 _6125_ (.A1(_3008_),
    .A2(_2533_),
    .B1(_2543_),
    .C1(_2546_),
    .X(_0205_));
 sky130_fd_sc_hd__nand2_1 _6126_ (.A(_2538_),
    .B(_1144_),
    .Y(_2547_));
 sky130_fd_sc_hd__o211a_1 _6127_ (.A1(_3011_),
    .A2(_2533_),
    .B1(_2543_),
    .C1(_2547_),
    .X(_0204_));
 sky130_fd_sc_hd__nand2_1 _6128_ (.A(_2538_),
    .B(_1149_),
    .Y(_2548_));
 sky130_fd_sc_hd__o211a_1 _6129_ (.A1(_3014_),
    .A2(_2533_),
    .B1(_2543_),
    .C1(_2548_),
    .X(_0203_));
 sky130_fd_sc_hd__nand2_1 _6130_ (.A(_2538_),
    .B(_1426_),
    .Y(_2549_));
 sky130_fd_sc_hd__o211a_1 _6131_ (.A1(_3017_),
    .A2(_2533_),
    .B1(_2543_),
    .C1(_2549_),
    .X(_0202_));
 sky130_fd_sc_hd__nand2_1 _6132_ (.A(_2531_),
    .B(_1574_),
    .Y(_2550_));
 sky130_fd_sc_hd__o211a_1 _6133_ (.A1(_3020_),
    .A2(_2533_),
    .B1(_2543_),
    .C1(_2550_),
    .X(_0201_));
 sky130_fd_sc_hd__nand2_1 _6134_ (.A(_2531_),
    .B(_3277_),
    .Y(_2551_));
 sky130_fd_sc_hd__o211a_1 _6135_ (.A1(_3023_),
    .A2(_2533_),
    .B1(_2543_),
    .C1(_2551_),
    .X(_0200_));
 sky130_fd_sc_hd__and4_1 _6136_ (.A(_2970_),
    .B(\egd_top.BitStream_buffer.buffer_index[6] ),
    .C(\egd_top.BitStream_buffer.buffer_index[5] ),
    .D(_2939_),
    .X(_2552_));
 sky130_fd_sc_hd__inv_2 _6137_ (.A(_2552_),
    .Y(_2553_));
 sky130_fd_sc_hd__buf_2 _6138_ (.A(_2553_),
    .X(_2554_));
 sky130_fd_sc_hd__buf_2 _6139_ (.A(_2553_),
    .X(_2555_));
 sky130_fd_sc_hd__nand2_1 _6140_ (.A(_2555_),
    .B(_1016_),
    .Y(_2556_));
 sky130_fd_sc_hd__o211a_1 _6141_ (.A1(_2966_),
    .A2(_2554_),
    .B1(_2543_),
    .C1(_2556_),
    .X(_0199_));
 sky130_fd_sc_hd__nand2_1 _6142_ (.A(_2555_),
    .B(_1169_),
    .Y(_2557_));
 sky130_fd_sc_hd__o211a_1 _6143_ (.A1(_2979_),
    .A2(_2554_),
    .B1(_2543_),
    .C1(_2557_),
    .X(_0198_));
 sky130_fd_sc_hd__buf_2 _6144_ (.A(_2904_),
    .X(_2558_));
 sky130_fd_sc_hd__nand2_1 _6145_ (.A(_2555_),
    .B(_3049_),
    .Y(_2559_));
 sky130_fd_sc_hd__o211a_1 _6146_ (.A1(_2982_),
    .A2(_2554_),
    .B1(_2558_),
    .C1(_2559_),
    .X(_0197_));
 sky130_fd_sc_hd__nand2_1 _6147_ (.A(_2555_),
    .B(_0709_),
    .Y(_2560_));
 sky130_fd_sc_hd__o211a_1 _6148_ (.A1(_2985_),
    .A2(_2554_),
    .B1(_2558_),
    .C1(_2560_),
    .X(_0196_));
 sky130_fd_sc_hd__buf_2 _6149_ (.A(_2553_),
    .X(_2561_));
 sky130_fd_sc_hd__nand2_1 _6150_ (.A(_2561_),
    .B(_0796_),
    .Y(_2562_));
 sky130_fd_sc_hd__o211a_1 _6151_ (.A1(_2988_),
    .A2(_2554_),
    .B1(_2558_),
    .C1(_2562_),
    .X(_0195_));
 sky130_fd_sc_hd__nand2_1 _6152_ (.A(_2561_),
    .B(_3102_),
    .Y(_2563_));
 sky130_fd_sc_hd__o211a_1 _6153_ (.A1(_2992_),
    .A2(_2554_),
    .B1(_2558_),
    .C1(_2563_),
    .X(_0194_));
 sky130_fd_sc_hd__nand2_1 _6154_ (.A(_2561_),
    .B(_0713_),
    .Y(_2564_));
 sky130_fd_sc_hd__o211a_1 _6155_ (.A1(_2995_),
    .A2(_2554_),
    .B1(_2558_),
    .C1(_2564_),
    .X(_0193_));
 sky130_fd_sc_hd__nand2_1 _6156_ (.A(_2561_),
    .B(_3085_),
    .Y(_2565_));
 sky130_fd_sc_hd__o211a_1 _6157_ (.A1(_2998_),
    .A2(_2554_),
    .B1(_2558_),
    .C1(_2565_),
    .X(_0192_));
 sky130_fd_sc_hd__nand2_1 _6158_ (.A(_2561_),
    .B(_0718_),
    .Y(_2566_));
 sky130_fd_sc_hd__o211a_1 _6159_ (.A1(_3001_),
    .A2(_2554_),
    .B1(_2558_),
    .C1(_2566_),
    .X(_0191_));
 sky130_fd_sc_hd__nand2_1 _6160_ (.A(_2561_),
    .B(_3119_),
    .Y(_2567_));
 sky130_fd_sc_hd__o211a_1 _6161_ (.A1(_3005_),
    .A2(_2554_),
    .B1(_2558_),
    .C1(_2567_),
    .X(_0190_));
 sky130_fd_sc_hd__nand2_1 _6162_ (.A(_2561_),
    .B(_0721_),
    .Y(_2568_));
 sky130_fd_sc_hd__o211a_1 _6163_ (.A1(_3008_),
    .A2(_2555_),
    .B1(_2558_),
    .C1(_2568_),
    .X(_0189_));
 sky130_fd_sc_hd__nand2_1 _6164_ (.A(_2561_),
    .B(_0804_),
    .Y(_2569_));
 sky130_fd_sc_hd__o211a_1 _6165_ (.A1(_3011_),
    .A2(_2555_),
    .B1(_2558_),
    .C1(_2569_),
    .X(_0188_));
 sky130_fd_sc_hd__buf_2 _6166_ (.A(_2904_),
    .X(_2570_));
 sky130_fd_sc_hd__nand2_1 _6167_ (.A(_2561_),
    .B(_1025_),
    .Y(_2571_));
 sky130_fd_sc_hd__o211a_1 _6168_ (.A1(_3014_),
    .A2(_2555_),
    .B1(_2570_),
    .C1(_2571_),
    .X(_0187_));
 sky130_fd_sc_hd__nand2_1 _6169_ (.A(_2561_),
    .B(_0727_),
    .Y(_2572_));
 sky130_fd_sc_hd__o211a_1 _6170_ (.A1(_3017_),
    .A2(_2555_),
    .B1(_2570_),
    .C1(_2572_),
    .X(_0186_));
 sky130_fd_sc_hd__nand2_1 _6171_ (.A(_2553_),
    .B(_0808_),
    .Y(_2573_));
 sky130_fd_sc_hd__o211a_1 _6172_ (.A1(_3020_),
    .A2(_2555_),
    .B1(_2570_),
    .C1(_2573_),
    .X(_0185_));
 sky130_fd_sc_hd__nand2_1 _6173_ (.A(_2553_),
    .B(_1035_),
    .Y(_2574_));
 sky130_fd_sc_hd__o211a_1 _6174_ (.A1(_3023_),
    .A2(_2555_),
    .B1(_2570_),
    .C1(_2574_),
    .X(_0184_));
 sky130_fd_sc_hd__inv_2 _6175_ (.A(\egd_top.BitStream_buffer.pc_previous[5] ),
    .Y(_2575_));
 sky130_fd_sc_hd__or2_1 _6176_ (.A(\egd_top.BitStream_buffer.pc_previous[1] ),
    .B(\egd_top.BitStream_buffer.exp_golomb_len[1] ),
    .X(_2576_));
 sky130_fd_sc_hd__nand2_1 _6177_ (.A(\egd_top.BitStream_buffer.pc_previous[1] ),
    .B(\egd_top.BitStream_buffer.exp_golomb_len[1] ),
    .Y(_2577_));
 sky130_fd_sc_hd__nand2_2 _6178_ (.A(_2576_),
    .B(_2577_),
    .Y(_2578_));
 sky130_fd_sc_hd__o21ai_4 _6179_ (.A1(_2925_),
    .A2(_2578_),
    .B1(_2577_),
    .Y(_2579_));
 sky130_fd_sc_hd__or2_1 _6180_ (.A(\egd_top.BitStream_buffer.pc_previous[2] ),
    .B(\egd_top.BitStream_buffer.exp_golomb_len[2] ),
    .X(_2580_));
 sky130_fd_sc_hd__nand2_1 _6181_ (.A(\egd_top.BitStream_buffer.pc_previous[2] ),
    .B(\egd_top.BitStream_buffer.exp_golomb_len[2] ),
    .Y(_2581_));
 sky130_fd_sc_hd__a21bo_2 _6182_ (.A1(_2579_),
    .A2(_2580_),
    .B1_N(_2581_),
    .X(_2582_));
 sky130_fd_sc_hd__or2_1 _6183_ (.A(\egd_top.BitStream_buffer.pc_previous[3] ),
    .B(\egd_top.BitStream_buffer.exp_golomb_len[3] ),
    .X(_2583_));
 sky130_fd_sc_hd__nand2_1 _6184_ (.A(\egd_top.BitStream_buffer.pc_previous[3] ),
    .B(\egd_top.BitStream_buffer.exp_golomb_len[3] ),
    .Y(_2584_));
 sky130_fd_sc_hd__a21bo_1 _6185_ (.A1(_2582_),
    .A2(_2583_),
    .B1_N(_2584_),
    .X(_2585_));
 sky130_fd_sc_hd__nand2_1 _6186_ (.A(_2585_),
    .B(\egd_top.BitStream_buffer.pc_previous[4] ),
    .Y(_2586_));
 sky130_fd_sc_hd__nor2_2 _6187_ (.A(_2575_),
    .B(_2586_),
    .Y(_2587_));
 sky130_fd_sc_hd__xor2_4 _6188_ (.A(\egd_top.BitStream_buffer.pc_previous[6] ),
    .B(_2587_),
    .X(\egd_top.BitStream_buffer.pc[6] ));
 sky130_fd_sc_hd__nand2_1 _6189_ (.A(_2902_),
    .B(\egd_top.BitStream_buffer.pc[6] ),
    .Y(_2588_));
 sky130_fd_sc_hd__inv_2 _6190_ (.A(_2588_),
    .Y(_0183_));
 sky130_fd_sc_hd__and2_1 _6191_ (.A(_2586_),
    .B(_2575_),
    .X(_2589_));
 sky130_fd_sc_hd__nor2_2 _6192_ (.A(_2587_),
    .B(_2589_),
    .Y(\egd_top.BitStream_buffer.pc[5] ));
 sky130_fd_sc_hd__nand2_1 _6193_ (.A(_2902_),
    .B(\egd_top.BitStream_buffer.pc[5] ),
    .Y(_2590_));
 sky130_fd_sc_hd__inv_2 _6194_ (.A(_2590_),
    .Y(_0182_));
 sky130_fd_sc_hd__or2_1 _6195_ (.A(\egd_top.BitStream_buffer.pc_previous[4] ),
    .B(_2585_),
    .X(_2591_));
 sky130_fd_sc_hd__and2_1 _6196_ (.A(_2591_),
    .B(_2586_),
    .X(_2592_));
 sky130_fd_sc_hd__clkbuf_2 _6197_ (.A(_2592_),
    .X(\egd_top.BitStream_buffer.pc[4] ));
 sky130_fd_sc_hd__nand2_1 _6198_ (.A(_2902_),
    .B(\egd_top.BitStream_buffer.pc[4] ),
    .Y(_2593_));
 sky130_fd_sc_hd__inv_2 _6199_ (.A(_2593_),
    .Y(_0181_));
 sky130_fd_sc_hd__nand2_2 _6200_ (.A(_2583_),
    .B(_2584_),
    .Y(_2594_));
 sky130_fd_sc_hd__xnor2_4 _6201_ (.A(_2594_),
    .B(_2582_),
    .Y(\egd_top.BitStream_buffer.pc[3] ));
 sky130_fd_sc_hd__nand2_1 _6202_ (.A(_2902_),
    .B(\egd_top.BitStream_buffer.pc[3] ),
    .Y(_2595_));
 sky130_fd_sc_hd__inv_2 _6203_ (.A(_2595_),
    .Y(_0180_));
 sky130_fd_sc_hd__nand2_2 _6204_ (.A(_2580_),
    .B(_2581_),
    .Y(_2596_));
 sky130_fd_sc_hd__xnor2_4 _6205_ (.A(_2596_),
    .B(_2579_),
    .Y(\egd_top.BitStream_buffer.pc[2] ));
 sky130_fd_sc_hd__nand2_1 _6206_ (.A(_2902_),
    .B(\egd_top.BitStream_buffer.pc[2] ),
    .Y(_2597_));
 sky130_fd_sc_hd__inv_2 _6207_ (.A(_2597_),
    .Y(_0179_));
 sky130_fd_sc_hd__xor2_4 _6208_ (.A(_2925_),
    .B(_2578_),
    .X(\egd_top.BitStream_buffer.pc[1] ));
 sky130_fd_sc_hd__nand2_1 _6209_ (.A(_2902_),
    .B(\egd_top.BitStream_buffer.pc[1] ),
    .Y(_2598_));
 sky130_fd_sc_hd__inv_2 _6210_ (.A(_2598_),
    .Y(_0178_));
 sky130_fd_sc_hd__or2_1 _6211_ (.A(_2905_),
    .B(_2929_),
    .X(_2599_));
 sky130_fd_sc_hd__inv_2 _6212_ (.A(_2599_),
    .Y(_0177_));
 sky130_fd_sc_hd__nor3_1 _6213_ (.A(_2967_),
    .B(\egd_top.BitStream_buffer.buffer_index[5] ),
    .C(_2971_),
    .Y(_2600_));
 sky130_fd_sc_hd__inv_2 _6214_ (.A(_2600_),
    .Y(_2601_));
 sky130_fd_sc_hd__buf_2 _6215_ (.A(_2601_),
    .X(_2602_));
 sky130_fd_sc_hd__buf_2 _6216_ (.A(_2601_),
    .X(_2603_));
 sky130_fd_sc_hd__nand2_1 _6217_ (.A(_2603_),
    .B(_3296_),
    .Y(_2604_));
 sky130_fd_sc_hd__o211a_1 _6218_ (.A1(_2966_),
    .A2(_2602_),
    .B1(_2570_),
    .C1(_2604_),
    .X(_0176_));
 sky130_fd_sc_hd__nand2_1 _6219_ (.A(_2603_),
    .B(_0767_),
    .Y(_2605_));
 sky130_fd_sc_hd__o211a_1 _6220_ (.A1(_2979_),
    .A2(_2602_),
    .B1(_2570_),
    .C1(_2605_),
    .X(_0175_));
 sky130_fd_sc_hd__nand2_1 _6221_ (.A(_2603_),
    .B(_0842_),
    .Y(_2606_));
 sky130_fd_sc_hd__o211a_1 _6222_ (.A1(_2982_),
    .A2(_2602_),
    .B1(_2570_),
    .C1(_2606_),
    .X(_0174_));
 sky130_fd_sc_hd__nand2_1 _6223_ (.A(_2603_),
    .B(_1007_),
    .Y(_2607_));
 sky130_fd_sc_hd__o211a_1 _6224_ (.A1(_2985_),
    .A2(_2602_),
    .B1(_2570_),
    .C1(_2607_),
    .X(_0173_));
 sky130_fd_sc_hd__buf_2 _6225_ (.A(_2601_),
    .X(_2608_));
 sky130_fd_sc_hd__nand2_1 _6226_ (.A(_2608_),
    .B(_1158_),
    .Y(_2609_));
 sky130_fd_sc_hd__o211a_1 _6227_ (.A1(_2988_),
    .A2(_2602_),
    .B1(_2570_),
    .C1(_2609_),
    .X(_0172_));
 sky130_fd_sc_hd__nand2_1 _6228_ (.A(_2608_),
    .B(_3317_),
    .Y(_2610_));
 sky130_fd_sc_hd__o211a_1 _6229_ (.A1(_2992_),
    .A2(_2602_),
    .B1(_2570_),
    .C1(_2610_),
    .X(_0171_));
 sky130_fd_sc_hd__buf_2 _6230_ (.A(_2904_),
    .X(_2611_));
 sky130_fd_sc_hd__nand2_1 _6231_ (.A(_2608_),
    .B(_0771_),
    .Y(_2612_));
 sky130_fd_sc_hd__o211a_1 _6232_ (.A1(_2995_),
    .A2(_2602_),
    .B1(_2611_),
    .C1(_2612_),
    .X(_0170_));
 sky130_fd_sc_hd__nand2_1 _6233_ (.A(_2608_),
    .B(_3306_),
    .Y(_2613_));
 sky130_fd_sc_hd__o211a_1 _6234_ (.A1(_2998_),
    .A2(_2602_),
    .B1(_2611_),
    .C1(_2613_),
    .X(_0169_));
 sky130_fd_sc_hd__nand2_1 _6235_ (.A(_2608_),
    .B(_0776_),
    .Y(_2614_));
 sky130_fd_sc_hd__o211a_1 _6236_ (.A1(_3001_),
    .A2(_2602_),
    .B1(_2611_),
    .C1(_2614_),
    .X(_0168_));
 sky130_fd_sc_hd__nand2_1 _6237_ (.A(_2608_),
    .B(_3328_),
    .Y(_2615_));
 sky130_fd_sc_hd__o211a_1 _6238_ (.A1(_3005_),
    .A2(_2602_),
    .B1(_2611_),
    .C1(_2615_),
    .X(_0167_));
 sky130_fd_sc_hd__nand2_1 _6239_ (.A(_2608_),
    .B(_0779_),
    .Y(_2616_));
 sky130_fd_sc_hd__o211a_1 _6240_ (.A1(_3008_),
    .A2(_2603_),
    .B1(_2611_),
    .C1(_2616_),
    .X(_0166_));
 sky130_fd_sc_hd__nand2_1 _6241_ (.A(_2608_),
    .B(_0850_),
    .Y(_2617_));
 sky130_fd_sc_hd__o211a_1 _6242_ (.A1(_3011_),
    .A2(_2603_),
    .B1(_2611_),
    .C1(_2617_),
    .X(_0165_));
 sky130_fd_sc_hd__nand2_1 _6243_ (.A(_2608_),
    .B(_1003_),
    .Y(_2618_));
 sky130_fd_sc_hd__o211a_1 _6244_ (.A1(_3014_),
    .A2(_2603_),
    .B1(_2611_),
    .C1(_2618_),
    .X(_0164_));
 sky130_fd_sc_hd__nand2_1 _6245_ (.A(_2608_),
    .B(_0324_),
    .Y(_2619_));
 sky130_fd_sc_hd__o211a_1 _6246_ (.A1(_3017_),
    .A2(_2603_),
    .B1(_2611_),
    .C1(_2619_),
    .X(_0163_));
 sky130_fd_sc_hd__nand2_1 _6247_ (.A(_2601_),
    .B(_0784_),
    .Y(_2620_));
 sky130_fd_sc_hd__o211a_1 _6248_ (.A1(_3020_),
    .A2(_2603_),
    .B1(_2611_),
    .C1(_2620_),
    .X(_0162_));
 sky130_fd_sc_hd__nand2_1 _6249_ (.A(_2601_),
    .B(_0854_),
    .Y(_2621_));
 sky130_fd_sc_hd__o211a_1 _6250_ (.A1(_3023_),
    .A2(_2603_),
    .B1(_2611_),
    .C1(_2621_),
    .X(_0161_));
 sky130_fd_sc_hd__nor2_1 _6251_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[13] ),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[12] ),
    .Y(_2622_));
 sky130_fd_sc_hd__nor2_2 _6252_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_valid_n ),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[15] ),
    .Y(_2623_));
 sky130_fd_sc_hd__inv_2 _6253_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[14] ),
    .Y(_2624_));
 sky130_fd_sc_hd__and3_1 _6254_ (.A(_2622_),
    .B(_2623_),
    .C(_2624_),
    .X(_2625_));
 sky130_fd_sc_hd__inv_2 _6255_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[3] ),
    .Y(_2626_));
 sky130_fd_sc_hd__inv_2 _6256_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[2] ),
    .Y(_2627_));
 sky130_fd_sc_hd__nand2_1 _6257_ (.A(_2626_),
    .B(_2627_),
    .Y(_2628_));
 sky130_fd_sc_hd__inv_2 _6258_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[4] ),
    .Y(_2629_));
 sky130_fd_sc_hd__a311oi_1 _6259_ (.A1(_2628_),
    .A2(_1945_),
    .A3(_2629_),
    .B1(\egd_top.BitStream_buffer.BitStream_buffer_output[7] ),
    .C1(\egd_top.BitStream_buffer.BitStream_buffer_output[6] ),
    .Y(_2630_));
 sky130_fd_sc_hd__inv_2 _6260_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[11] ),
    .Y(_2631_));
 sky130_fd_sc_hd__nand2_1 _6261_ (.A(_2622_),
    .B(_2631_),
    .Y(_2632_));
 sky130_fd_sc_hd__or2_1 _6262_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[10] ),
    .B(_2632_),
    .X(_2633_));
 sky130_fd_sc_hd__inv_2 _6263_ (.A(_2633_),
    .Y(_2634_));
 sky130_fd_sc_hd__clkinv_2 _6264_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[9] ),
    .Y(_2635_));
 sky130_fd_sc_hd__and3_1 _6265_ (.A(_2634_),
    .B(_2635_),
    .C(_1586_),
    .X(_2636_));
 sky130_fd_sc_hd__clkinv_4 _6266_ (.A(_2636_),
    .Y(_2637_));
 sky130_fd_sc_hd__nand2_1 _6267_ (.A(_2633_),
    .B(_2622_),
    .Y(_2638_));
 sky130_fd_sc_hd__nand2_1 _6268_ (.A(_2623_),
    .B(_2624_),
    .Y(_2639_));
 sky130_fd_sc_hd__inv_2 _6269_ (.A(_2639_),
    .Y(_2640_));
 sky130_fd_sc_hd__nand2_1 _6270_ (.A(_2638_),
    .B(_2640_),
    .Y(_2641_));
 sky130_fd_sc_hd__inv_2 _6271_ (.A(_2641_),
    .Y(_2642_));
 sky130_fd_sc_hd__o21ai_1 _6272_ (.A1(_2630_),
    .A2(_2637_),
    .B1(_2642_),
    .Y(_2643_));
 sky130_fd_sc_hd__nor2_1 _6273_ (.A(_2625_),
    .B(_2643_),
    .Y(_2644_));
 sky130_fd_sc_hd__nand2_1 _6274_ (.A(_2627_),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[1] ),
    .Y(_2645_));
 sky130_fd_sc_hd__nand2_1 _6275_ (.A(_2645_),
    .B(_2626_),
    .Y(_2646_));
 sky130_fd_sc_hd__nand2_1 _6276_ (.A(_2646_),
    .B(_2629_),
    .Y(_2647_));
 sky130_fd_sc_hd__nand2_1 _6277_ (.A(_2647_),
    .B(_1945_),
    .Y(_2648_));
 sky130_fd_sc_hd__inv_2 _6278_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[6] ),
    .Y(_2649_));
 sky130_fd_sc_hd__nand2_1 _6279_ (.A(_2648_),
    .B(_2649_),
    .Y(_2650_));
 sky130_fd_sc_hd__nand2_1 _6280_ (.A(_2650_),
    .B(_1705_),
    .Y(_2651_));
 sky130_fd_sc_hd__nand2_1 _6281_ (.A(_2651_),
    .B(_1586_),
    .Y(_2652_));
 sky130_fd_sc_hd__nand2_1 _6282_ (.A(_2652_),
    .B(_2635_),
    .Y(_2653_));
 sky130_fd_sc_hd__nand2_1 _6283_ (.A(_2653_),
    .B(_2634_),
    .Y(_2654_));
 sky130_fd_sc_hd__inv_2 _6284_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[12] ),
    .Y(_2655_));
 sky130_fd_sc_hd__a21oi_1 _6285_ (.A1(_2655_),
    .A2(\egd_top.BitStream_buffer.BitStream_buffer_output[11] ),
    .B1(\egd_top.BitStream_buffer.BitStream_buffer_output[13] ),
    .Y(_2656_));
 sky130_fd_sc_hd__nand2_1 _6286_ (.A(_2654_),
    .B(_2656_),
    .Y(_2657_));
 sky130_fd_sc_hd__nand2_1 _6287_ (.A(_2657_),
    .B(_2624_),
    .Y(_2658_));
 sky130_fd_sc_hd__nand2_1 _6288_ (.A(_2658_),
    .B(_2623_),
    .Y(_2659_));
 sky130_fd_sc_hd__nand2_1 _6289_ (.A(_2644_),
    .B(_2659_),
    .Y(_2660_));
 sky130_fd_sc_hd__or2_1 _6290_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[11] ),
    .B(_2660_),
    .X(_2661_));
 sky130_fd_sc_hd__inv_2 _6291_ (.A(_2623_),
    .Y(_2662_));
 sky130_fd_sc_hd__a21oi_2 _6292_ (.A1(_2657_),
    .A2(_2624_),
    .B1(_2662_),
    .Y(_2663_));
 sky130_fd_sc_hd__nand2_1 _6293_ (.A(_2663_),
    .B(_2644_),
    .Y(_2664_));
 sky130_fd_sc_hd__inv_2 _6294_ (.A(_2664_),
    .Y(_2665_));
 sky130_fd_sc_hd__nand2_1 _6295_ (.A(_2665_),
    .B(_2635_),
    .Y(_2666_));
 sky130_fd_sc_hd__nand2_1 _6296_ (.A(_2637_),
    .B(_2625_),
    .Y(_2667_));
 sky130_fd_sc_hd__nor2_1 _6297_ (.A(_2642_),
    .B(_2667_),
    .Y(_2668_));
 sky130_fd_sc_hd__nand2_2 _6298_ (.A(_2659_),
    .B(_2668_),
    .Y(_2669_));
 sky130_fd_sc_hd__inv_2 _6299_ (.A(_2669_),
    .Y(_2670_));
 sky130_fd_sc_hd__nand2_1 _6300_ (.A(_2670_),
    .B(_1705_),
    .Y(_2671_));
 sky130_fd_sc_hd__nand3_1 _6301_ (.A(_2661_),
    .B(_2666_),
    .C(_2671_),
    .Y(_2672_));
 sky130_fd_sc_hd__nand2_1 _6302_ (.A(_2663_),
    .B(_2668_),
    .Y(_2673_));
 sky130_fd_sc_hd__or3_1 _6303_ (.A(_2624_),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[13] ),
    .C(_2662_),
    .X(_2674_));
 sky130_fd_sc_hd__o21a_1 _6304_ (.A1(\egd_top.BitStream_buffer.BitStream_buffer_output[5] ),
    .A2(_2673_),
    .B1(_2674_),
    .X(_2675_));
 sky130_fd_sc_hd__nor2b_2 _6305_ (.A(_2672_),
    .B_N(_2675_),
    .Y(_2676_));
 sky130_fd_sc_hd__nor2_1 _6306_ (.A(_2641_),
    .B(_2667_),
    .Y(_2677_));
 sky130_fd_sc_hd__nand3_4 _6307_ (.A(_2658_),
    .B(_2677_),
    .C(_2623_),
    .Y(_2678_));
 sky130_fd_sc_hd__nand2_1 _6308_ (.A(_2678_),
    .B(_2626_),
    .Y(_2679_));
 sky130_fd_sc_hd__o21ai_2 _6309_ (.A1(\egd_top.BitStream_buffer.BitStream_buffer_output[1] ),
    .A2(_2678_),
    .B1(_2679_),
    .Y(_2680_));
 sky130_fd_sc_hd__buf_6 _6310_ (.A(_2677_),
    .X(_2681_));
 sky130_fd_sc_hd__nand2_1 _6311_ (.A(_2680_),
    .B(_2681_),
    .Y(_2682_));
 sky130_fd_sc_hd__nand2_1 _6312_ (.A(_2676_),
    .B(_2682_),
    .Y(_2683_));
 sky130_fd_sc_hd__clkbuf_4 _6313_ (.A(_2924_),
    .X(_2684_));
 sky130_fd_sc_hd__nand2_2 _6314_ (.A(_2683_),
    .B(_2684_),
    .Y(_2685_));
 sky130_fd_sc_hd__nor2_1 _6315_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[6] ),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[5] ),
    .Y(_2686_));
 sky130_fd_sc_hd__inv_2 _6316_ (.A(_2686_),
    .Y(_2687_));
 sky130_fd_sc_hd__nor2_1 _6317_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[7] ),
    .B(_2687_),
    .Y(_2688_));
 sky130_fd_sc_hd__a21oi_1 _6318_ (.A1(_2629_),
    .A2(_2688_),
    .B1(_2637_),
    .Y(_2689_));
 sky130_fd_sc_hd__nor2b_1 _6319_ (.A(_2689_),
    .B_N(_2625_),
    .Y(_2690_));
 sky130_fd_sc_hd__or3b_1 _6320_ (.A(_2663_),
    .B(_2690_),
    .C_N(_2643_),
    .X(_2691_));
 sky130_fd_sc_hd__nand2_1 _6321_ (.A(_2636_),
    .B(_2640_),
    .Y(_2692_));
 sky130_fd_sc_hd__nand2_1 _6322_ (.A(_2691_),
    .B(_2692_),
    .Y(_2693_));
 sky130_fd_sc_hd__inv_2 _6323_ (.A(_2693_),
    .Y(_2694_));
 sky130_fd_sc_hd__nand2_2 _6324_ (.A(_2694_),
    .B(_2684_),
    .Y(_2695_));
 sky130_fd_sc_hd__nor3b_1 _6325_ (.A(net21),
    .B(\egd_top.exp_golomb_decoding.te_range[2] ),
    .C_N(net20),
    .Y(_2696_));
 sky130_fd_sc_hd__nand2_1 _6326_ (.A(net18),
    .B(net17),
    .Y(_2697_));
 sky130_fd_sc_hd__inv_2 _6327_ (.A(_2697_),
    .Y(_2698_));
 sky130_fd_sc_hd__and2_1 _6328_ (.A(_2696_),
    .B(_2698_),
    .X(_2699_));
 sky130_fd_sc_hd__inv_2 _6329_ (.A(_2699_),
    .Y(_2700_));
 sky130_fd_sc_hd__a21oi_4 _6330_ (.A1(_2676_),
    .A2(_2682_),
    .B1(_2926_),
    .Y(_2701_));
 sky130_fd_sc_hd__nor2_1 _6331_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[8] ),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[7] ),
    .Y(_2702_));
 sky130_fd_sc_hd__inv_2 _6332_ (.A(_2702_),
    .Y(_2703_));
 sky130_fd_sc_hd__nand2_1 _6333_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[8] ),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[7] ),
    .Y(_2704_));
 sky130_fd_sc_hd__a21o_1 _6334_ (.A1(_2703_),
    .A2(_2704_),
    .B1(_2669_),
    .X(_2705_));
 sky130_fd_sc_hd__or3_1 _6335_ (.A(_2624_),
    .B(_0933_),
    .C(_2662_),
    .X(_2706_));
 sky130_fd_sc_hd__nand2_1 _6336_ (.A(_2705_),
    .B(_2706_),
    .Y(_2707_));
 sky130_fd_sc_hd__nand2_1 _6337_ (.A(_2655_),
    .B(_2631_),
    .Y(_2708_));
 sky130_fd_sc_hd__nand2_1 _6338_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[12] ),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[11] ),
    .Y(_2709_));
 sky130_fd_sc_hd__and2_1 _6339_ (.A(_2708_),
    .B(_2709_),
    .X(_2710_));
 sky130_fd_sc_hd__or2_1 _6340_ (.A(_2710_),
    .B(_2660_),
    .X(_2711_));
 sky130_fd_sc_hd__nor2_1 _6341_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[10] ),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[9] ),
    .Y(_2712_));
 sky130_fd_sc_hd__inv_2 _6342_ (.A(_2712_),
    .Y(_2713_));
 sky130_fd_sc_hd__nand2_1 _6343_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[10] ),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[9] ),
    .Y(_2714_));
 sky130_fd_sc_hd__nand2_1 _6344_ (.A(_2713_),
    .B(_2714_),
    .Y(_2715_));
 sky130_fd_sc_hd__nand2_1 _6345_ (.A(_2665_),
    .B(_2715_),
    .Y(_2716_));
 sky130_fd_sc_hd__inv_2 _6346_ (.A(_2673_),
    .Y(_2717_));
 sky130_fd_sc_hd__nand2_1 _6347_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[6] ),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[5] ),
    .Y(_2718_));
 sky130_fd_sc_hd__nand2_1 _6348_ (.A(_2687_),
    .B(_2718_),
    .Y(_2719_));
 sky130_fd_sc_hd__nand2_1 _6349_ (.A(_2717_),
    .B(_2719_),
    .Y(_2720_));
 sky130_fd_sc_hd__nand3_1 _6350_ (.A(_2711_),
    .B(_2716_),
    .C(_2720_),
    .Y(_2721_));
 sky130_fd_sc_hd__nor2_1 _6351_ (.A(_2707_),
    .B(_2721_),
    .Y(_2722_));
 sky130_fd_sc_hd__buf_6 _6352_ (.A(_2678_),
    .X(_2723_));
 sky130_fd_sc_hd__nand2_1 _6353_ (.A(_2723_),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[4] ),
    .Y(_2724_));
 sky130_fd_sc_hd__o21ai_1 _6354_ (.A1(_2627_),
    .A2(_2723_),
    .B1(_2724_),
    .Y(_2725_));
 sky130_fd_sc_hd__nand2_1 _6355_ (.A(_2680_),
    .B(_2725_),
    .Y(_2726_));
 sky130_fd_sc_hd__nand3_1 _6356_ (.A(_2663_),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[1] ),
    .C(_2681_),
    .Y(_2727_));
 sky130_fd_sc_hd__nand2_1 _6357_ (.A(_2678_),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[3] ),
    .Y(_2728_));
 sky130_fd_sc_hd__nand2_1 _6358_ (.A(_2727_),
    .B(_2728_),
    .Y(_2729_));
 sky130_fd_sc_hd__nand3_1 _6359_ (.A(_2663_),
    .B(_2627_),
    .C(_2681_),
    .Y(_2730_));
 sky130_fd_sc_hd__nand2_1 _6360_ (.A(_2678_),
    .B(_2629_),
    .Y(_2731_));
 sky130_fd_sc_hd__nand2_1 _6361_ (.A(_2730_),
    .B(_2731_),
    .Y(_2732_));
 sky130_fd_sc_hd__nand2_1 _6362_ (.A(_2729_),
    .B(_2732_),
    .Y(_2733_));
 sky130_fd_sc_hd__nand3_1 _6363_ (.A(_2726_),
    .B(_2733_),
    .C(_2681_),
    .Y(_2734_));
 sky130_fd_sc_hd__nand2_1 _6364_ (.A(_2722_),
    .B(_2734_),
    .Y(_2735_));
 sky130_fd_sc_hd__nor2_1 _6365_ (.A(net17),
    .B(_2922_),
    .Y(_2736_));
 sky130_fd_sc_hd__inv_2 _6366_ (.A(_2736_),
    .Y(_2737_));
 sky130_fd_sc_hd__nand2_1 _6367_ (.A(_2735_),
    .B(_2684_),
    .Y(_2738_));
 sky130_fd_sc_hd__inv_2 _6368_ (.A(_2738_),
    .Y(_2739_));
 sky130_fd_sc_hd__nor2_1 _6369_ (.A(_2739_),
    .B(_2701_),
    .Y(_2740_));
 sky130_fd_sc_hd__a211o_1 _6370_ (.A1(_2701_),
    .A2(_2735_),
    .B1(_2737_),
    .C1(_2740_),
    .X(_2741_));
 sky130_fd_sc_hd__o221ai_4 _6371_ (.A1(_2923_),
    .A2(_2685_),
    .B1(_2695_),
    .B2(_2700_),
    .C1(_2741_),
    .Y(net20));
 sky130_fd_sc_hd__nand2_1 _6372_ (.A(_2680_),
    .B(_2732_),
    .Y(_2742_));
 sky130_fd_sc_hd__nand3_1 _6373_ (.A(_2663_),
    .B(_2626_),
    .C(_2681_),
    .Y(_2743_));
 sky130_fd_sc_hd__nand2_1 _6374_ (.A(_2678_),
    .B(_1945_),
    .Y(_2744_));
 sky130_fd_sc_hd__nand2_1 _6375_ (.A(_2743_),
    .B(_2744_),
    .Y(_2745_));
 sky130_fd_sc_hd__nand2_1 _6376_ (.A(_2742_),
    .B(_2745_),
    .Y(_2746_));
 sky130_fd_sc_hd__nand2_1 _6377_ (.A(_2723_),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[5] ),
    .Y(_2747_));
 sky130_fd_sc_hd__o21ai_1 _6378_ (.A1(_2626_),
    .A2(_2723_),
    .B1(_2747_),
    .Y(_2748_));
 sky130_fd_sc_hd__nand3_1 _6379_ (.A(_2680_),
    .B(_2748_),
    .C(_2732_),
    .Y(_2749_));
 sky130_fd_sc_hd__nand3_1 _6380_ (.A(_2746_),
    .B(_2749_),
    .C(_2681_),
    .Y(_2750_));
 sky130_fd_sc_hd__nor2_1 _6381_ (.A(_1705_),
    .B(_2686_),
    .Y(_2751_));
 sky130_fd_sc_hd__o21ai_1 _6382_ (.A1(_2688_),
    .A2(_2751_),
    .B1(_2717_),
    .Y(_2752_));
 sky130_fd_sc_hd__nor2_1 _6383_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[9] ),
    .B(_2703_),
    .Y(_2753_));
 sky130_fd_sc_hd__nor2_1 _6384_ (.A(_2635_),
    .B(_2702_),
    .Y(_2754_));
 sky130_fd_sc_hd__o21ai_1 _6385_ (.A1(_2753_),
    .A2(_2754_),
    .B1(_2670_),
    .Y(_2755_));
 sky130_fd_sc_hd__nand2_1 _6386_ (.A(_2752_),
    .B(_2755_),
    .Y(_2756_));
 sky130_fd_sc_hd__nand2_1 _6387_ (.A(_2712_),
    .B(_2631_),
    .Y(_2757_));
 sky130_fd_sc_hd__nand2_1 _6388_ (.A(_2713_),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[11] ),
    .Y(_2758_));
 sky130_fd_sc_hd__a21o_1 _6389_ (.A1(_2757_),
    .A2(_2758_),
    .B1(_2664_),
    .X(_2759_));
 sky130_fd_sc_hd__nand2_1 _6390_ (.A(_2708_),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[13] ),
    .Y(_2760_));
 sky130_fd_sc_hd__a21o_1 _6391_ (.A1(_2632_),
    .A2(_2760_),
    .B1(_2660_),
    .X(_2761_));
 sky130_fd_sc_hd__nand2_1 _6392_ (.A(_2759_),
    .B(_2761_),
    .Y(_2762_));
 sky130_fd_sc_hd__nor2_1 _6393_ (.A(_2756_),
    .B(_2762_),
    .Y(_2763_));
 sky130_fd_sc_hd__nand2_1 _6394_ (.A(_2750_),
    .B(_2763_),
    .Y(_2764_));
 sky130_fd_sc_hd__nand2_1 _6395_ (.A(_2739_),
    .B(_2764_),
    .Y(_2765_));
 sky130_fd_sc_hd__nand2_1 _6396_ (.A(_2764_),
    .B(_2684_),
    .Y(_2766_));
 sky130_fd_sc_hd__nand2_1 _6397_ (.A(_2766_),
    .B(_2738_),
    .Y(_2767_));
 sky130_fd_sc_hd__and3_1 _6398_ (.A(_2765_),
    .B(_2767_),
    .C(_2736_),
    .X(_2768_));
 sky130_fd_sc_hd__a31o_2 _6399_ (.A1(net17),
    .A2(_2700_),
    .A3(_2739_),
    .B1(_2768_),
    .X(net21));
 sky130_fd_sc_hd__nand2_1 _6400_ (.A(_2767_),
    .B(_2685_),
    .Y(_2769_));
 sky130_fd_sc_hd__nand2_1 _6401_ (.A(_2769_),
    .B(_2765_),
    .Y(_2770_));
 sky130_fd_sc_hd__nor2_1 _6402_ (.A(_2729_),
    .B(_2725_),
    .Y(_2771_));
 sky130_fd_sc_hd__nand2_1 _6403_ (.A(_2723_),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[6] ),
    .Y(_2772_));
 sky130_fd_sc_hd__o21ai_1 _6404_ (.A1(_2629_),
    .A2(_2723_),
    .B1(_2772_),
    .Y(_2773_));
 sky130_fd_sc_hd__nand3_1 _6405_ (.A(_2771_),
    .B(_2745_),
    .C(_2773_),
    .Y(_2774_));
 sky130_fd_sc_hd__nand3_1 _6406_ (.A(_2680_),
    .B(_2732_),
    .C(_2745_),
    .Y(_2775_));
 sky130_fd_sc_hd__nand2_1 _6407_ (.A(_2723_),
    .B(_2649_),
    .Y(_2776_));
 sky130_fd_sc_hd__o21ai_1 _6408_ (.A1(\egd_top.BitStream_buffer.BitStream_buffer_output[4] ),
    .A2(_2723_),
    .B1(_2776_),
    .Y(_2777_));
 sky130_fd_sc_hd__nand2_1 _6409_ (.A(_2775_),
    .B(_2777_),
    .Y(_2778_));
 sky130_fd_sc_hd__nand3_1 _6410_ (.A(_2774_),
    .B(_2778_),
    .C(_2681_),
    .Y(_2779_));
 sky130_fd_sc_hd__xnor2_1 _6411_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[10] ),
    .B(_2753_),
    .Y(_2780_));
 sky130_fd_sc_hd__nor2_1 _6412_ (.A(_2687_),
    .B(_2703_),
    .Y(_2781_));
 sky130_fd_sc_hd__nor2_1 _6413_ (.A(_1586_),
    .B(_2688_),
    .Y(_2782_));
 sky130_fd_sc_hd__o21ai_1 _6414_ (.A1(_2781_),
    .A2(_2782_),
    .B1(_2717_),
    .Y(_2783_));
 sky130_fd_sc_hd__nand3_1 _6415_ (.A(_2665_),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[12] ),
    .C(_2757_),
    .Y(_2784_));
 sky130_fd_sc_hd__o211a_1 _6416_ (.A1(_2669_),
    .A2(_2780_),
    .B1(_2783_),
    .C1(_2784_),
    .X(_2785_));
 sky130_fd_sc_hd__a21oi_1 _6417_ (.A1(_2779_),
    .A2(_2785_),
    .B1(_2926_),
    .Y(_2786_));
 sky130_fd_sc_hd__nand2_1 _6418_ (.A(_2770_),
    .B(_2786_),
    .Y(_2787_));
 sky130_fd_sc_hd__nand2_1 _6419_ (.A(_2779_),
    .B(_2785_),
    .Y(_2788_));
 sky130_fd_sc_hd__nand2_1 _6420_ (.A(_2788_),
    .B(_2684_),
    .Y(_2789_));
 sky130_fd_sc_hd__nand3_1 _6421_ (.A(_2769_),
    .B(_2765_),
    .C(_2789_),
    .Y(_2790_));
 sky130_fd_sc_hd__nand3_1 _6422_ (.A(_2787_),
    .B(_2736_),
    .C(_2790_),
    .Y(_2791_));
 sky130_fd_sc_hd__or3_1 _6423_ (.A(_2923_),
    .B(_2699_),
    .C(_2766_),
    .X(_2792_));
 sky130_fd_sc_hd__nand2_2 _6424_ (.A(_2791_),
    .B(_2792_),
    .Y(net22));
 sky130_fd_sc_hd__nand2_1 _6425_ (.A(net20),
    .B(net21),
    .Y(_2793_));
 sky130_fd_sc_hd__inv_2 _6426_ (.A(_2793_),
    .Y(_2794_));
 sky130_fd_sc_hd__nand2_1 _6427_ (.A(net22),
    .B(_2794_),
    .Y(_2795_));
 sky130_fd_sc_hd__nand3_1 _6428_ (.A(_2791_),
    .B(_2793_),
    .C(_2792_),
    .Y(_2796_));
 sky130_fd_sc_hd__nand3_1 _6429_ (.A(_2795_),
    .B(_2698_),
    .C(_2796_),
    .Y(_2797_));
 sky130_fd_sc_hd__inv_2 _6430_ (.A(_2797_),
    .Y(\egd_top.exp_golomb_decoding.te_range[2] ));
 sky130_fd_sc_hd__nand2_1 _6431_ (.A(_2700_),
    .B(_2684_),
    .Y(_2798_));
 sky130_fd_sc_hd__or2_1 _6432_ (.A(_2798_),
    .B(_2659_),
    .X(_2799_));
 sky130_fd_sc_hd__inv_2 _6433_ (.A(_2799_),
    .Y(\egd_top.BitStream_buffer.exp_golomb_len[1] ));
 sky130_fd_sc_hd__nor2_1 _6434_ (.A(_2798_),
    .B(_2643_),
    .Y(\egd_top.BitStream_buffer.exp_golomb_len[2] ));
 sky130_fd_sc_hd__and3_1 _6435_ (.A(_2690_),
    .B(_2684_),
    .C(_2700_),
    .X(_2800_));
 sky130_fd_sc_hd__clkbuf_1 _6436_ (.A(_2800_),
    .X(\egd_top.BitStream_buffer.exp_golomb_len[3] ));
 sky130_fd_sc_hd__nand2_1 _6437_ (.A(_2777_),
    .B(_2745_),
    .Y(_2801_));
 sky130_fd_sc_hd__nor2_1 _6438_ (.A(_2742_),
    .B(_2801_),
    .Y(_2802_));
 sky130_fd_sc_hd__nand2_1 _6439_ (.A(_2678_),
    .B(_1705_),
    .Y(_2803_));
 sky130_fd_sc_hd__o21ai_2 _6440_ (.A1(\egd_top.BitStream_buffer.BitStream_buffer_output[5] ),
    .A2(_2678_),
    .B1(_2803_),
    .Y(_2804_));
 sky130_fd_sc_hd__inv_2 _6441_ (.A(_2804_),
    .Y(_2805_));
 sky130_fd_sc_hd__nand2_1 _6442_ (.A(_2802_),
    .B(_2805_),
    .Y(_2806_));
 sky130_fd_sc_hd__nor2_1 _6443_ (.A(_2748_),
    .B(_2773_),
    .Y(_2807_));
 sky130_fd_sc_hd__nand2_1 _6444_ (.A(_2807_),
    .B(_2771_),
    .Y(_2808_));
 sky130_fd_sc_hd__nand2_1 _6445_ (.A(_2808_),
    .B(_2804_),
    .Y(_2809_));
 sky130_fd_sc_hd__nand3_1 _6446_ (.A(_2806_),
    .B(_2809_),
    .C(_2681_),
    .Y(_2810_));
 sky130_fd_sc_hd__inv_2 _6447_ (.A(_2781_),
    .Y(_2811_));
 sky130_fd_sc_hd__nor2_1 _6448_ (.A(_2635_),
    .B(_2811_),
    .Y(_2812_));
 sky130_fd_sc_hd__nor2_1 _6449_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[9] ),
    .B(_2781_),
    .Y(_2813_));
 sky130_fd_sc_hd__a21o_1 _6450_ (.A1(_2712_),
    .A2(_2702_),
    .B1(_2631_),
    .X(_2814_));
 sky130_fd_sc_hd__o32a_1 _6451_ (.A1(_2812_),
    .A2(_2813_),
    .A3(_2673_),
    .B1(_2669_),
    .B2(_2814_),
    .X(_2815_));
 sky130_fd_sc_hd__nand2_1 _6452_ (.A(_2810_),
    .B(_2815_),
    .Y(_2816_));
 sky130_fd_sc_hd__nand2_1 _6453_ (.A(_2816_),
    .B(_2701_),
    .Y(_2817_));
 sky130_fd_sc_hd__nand3_1 _6454_ (.A(_2739_),
    .B(_2788_),
    .C(_2764_),
    .Y(_2818_));
 sky130_fd_sc_hd__nor2_1 _6455_ (.A(_2817_),
    .B(_2818_),
    .Y(_2819_));
 sky130_fd_sc_hd__inv_2 _6456_ (.A(_2816_),
    .Y(_2820_));
 sky130_fd_sc_hd__a31o_1 _6457_ (.A1(_2818_),
    .A2(_2820_),
    .A3(_2701_),
    .B1(_2737_),
    .X(_2821_));
 sky130_fd_sc_hd__nor2_1 _6458_ (.A(_2819_),
    .B(_2821_),
    .Y(_2822_));
 sky130_fd_sc_hd__nand2_1 _6459_ (.A(_2816_),
    .B(_2684_),
    .Y(_2823_));
 sky130_fd_sc_hd__inv_2 _6460_ (.A(_2823_),
    .Y(_2824_));
 sky130_fd_sc_hd__o21ai_1 _6461_ (.A1(_2735_),
    .A2(_2764_),
    .B1(_2684_),
    .Y(_2825_));
 sky130_fd_sc_hd__nand2_1 _6462_ (.A(_2825_),
    .B(_2789_),
    .Y(_2826_));
 sky130_fd_sc_hd__nor2_1 _6463_ (.A(_2824_),
    .B(_2826_),
    .Y(_2827_));
 sky130_fd_sc_hd__nor2_1 _6464_ (.A(_2767_),
    .B(_2786_),
    .Y(_2828_));
 sky130_fd_sc_hd__nor2_1 _6465_ (.A(_2823_),
    .B(_2828_),
    .Y(_2829_));
 sky130_fd_sc_hd__o21ai_1 _6466_ (.A1(_2827_),
    .A2(_2829_),
    .B1(_2685_),
    .Y(_2830_));
 sky130_fd_sc_hd__nand2_1 _6467_ (.A(_2822_),
    .B(_2830_),
    .Y(_2831_));
 sky130_fd_sc_hd__or3_2 _6468_ (.A(_2923_),
    .B(_2699_),
    .C(_2693_),
    .X(_2832_));
 sky130_fd_sc_hd__inv_2 _6469_ (.A(_2832_),
    .Y(_2833_));
 sky130_fd_sc_hd__nand2_1 _6470_ (.A(_2833_),
    .B(_2788_),
    .Y(_2834_));
 sky130_fd_sc_hd__nand2_1 _6471_ (.A(_2831_),
    .B(_2834_),
    .Y(net23));
 sky130_fd_sc_hd__nand2_1 _6472_ (.A(_2827_),
    .B(_2685_),
    .Y(_2835_));
 sky130_fd_sc_hd__o21ai_1 _6473_ (.A1(_2820_),
    .A2(_2818_),
    .B1(_2701_),
    .Y(_2836_));
 sky130_fd_sc_hd__nand2_1 _6474_ (.A(_2835_),
    .B(_2836_),
    .Y(_2837_));
 sky130_fd_sc_hd__nand3_1 _6475_ (.A(_2807_),
    .B(_2771_),
    .C(_2804_),
    .Y(_2838_));
 sky130_fd_sc_hd__nor2_1 _6476_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[6] ),
    .B(_2723_),
    .Y(_2839_));
 sky130_fd_sc_hd__nor2_1 _6477_ (.A(_1586_),
    .B(_2839_),
    .Y(_2840_));
 sky130_fd_sc_hd__inv_2 _6478_ (.A(_2840_),
    .Y(_2841_));
 sky130_fd_sc_hd__nand2_1 _6479_ (.A(_2838_),
    .B(_2841_),
    .Y(_2842_));
 sky130_fd_sc_hd__nand3_1 _6480_ (.A(_2802_),
    .B(_2804_),
    .C(_2840_),
    .Y(_2843_));
 sky130_fd_sc_hd__nand3_1 _6481_ (.A(_2842_),
    .B(_2843_),
    .C(_2681_),
    .Y(_2844_));
 sky130_fd_sc_hd__o21ai_1 _6482_ (.A1(_2715_),
    .A2(_2811_),
    .B1(_2717_),
    .Y(_2845_));
 sky130_fd_sc_hd__nand2_1 _6483_ (.A(_2844_),
    .B(_2845_),
    .Y(_2846_));
 sky130_fd_sc_hd__nand2_1 _6484_ (.A(_2846_),
    .B(_2684_),
    .Y(_2847_));
 sky130_fd_sc_hd__nand2_1 _6485_ (.A(_2837_),
    .B(_2847_),
    .Y(_2848_));
 sky130_fd_sc_hd__a21oi_2 _6486_ (.A1(_2844_),
    .A2(_2845_),
    .B1(_2926_),
    .Y(_2849_));
 sky130_fd_sc_hd__nand3_1 _6487_ (.A(_2835_),
    .B(_2849_),
    .C(_2836_),
    .Y(_2850_));
 sky130_fd_sc_hd__nand3_1 _6488_ (.A(_2848_),
    .B(_2923_),
    .C(_2850_),
    .Y(_2851_));
 sky130_fd_sc_hd__o21ai_2 _6489_ (.A1(_2820_),
    .A2(_2832_),
    .B1(_2851_),
    .Y(net24));
 sky130_fd_sc_hd__nand3_1 _6490_ (.A(_2828_),
    .B(_2823_),
    .C(_2847_),
    .Y(_2852_));
 sky130_fd_sc_hd__nor2_1 _6491_ (.A(_2840_),
    .B(_2805_),
    .Y(_2853_));
 sky130_fd_sc_hd__nand2_1 _6492_ (.A(_2802_),
    .B(_2853_),
    .Y(_2854_));
 sky130_fd_sc_hd__inv_2 _6493_ (.A(_2723_),
    .Y(_2855_));
 sky130_fd_sc_hd__nand2_1 _6494_ (.A(_2855_),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[7] ),
    .Y(_2856_));
 sky130_fd_sc_hd__nand3_1 _6495_ (.A(_2854_),
    .B(_2635_),
    .C(_2856_),
    .Y(_2857_));
 sky130_fd_sc_hd__nand2_1 _6496_ (.A(_2856_),
    .B(_2635_),
    .Y(_2858_));
 sky130_fd_sc_hd__nand3_1 _6497_ (.A(_2802_),
    .B(_2853_),
    .C(_2858_),
    .Y(_2859_));
 sky130_fd_sc_hd__nand3_2 _6498_ (.A(_2857_),
    .B(_2681_),
    .C(_2859_),
    .Y(_2860_));
 sky130_fd_sc_hd__nor2_1 _6499_ (.A(_2695_),
    .B(_2860_),
    .Y(_2861_));
 sky130_fd_sc_hd__nand2_1 _6500_ (.A(_2852_),
    .B(_2861_),
    .Y(_2862_));
 sky130_fd_sc_hd__nor2_1 _6501_ (.A(_2926_),
    .B(_2860_),
    .Y(_2863_));
 sky130_fd_sc_hd__nor2_1 _6502_ (.A(_2863_),
    .B(_2849_),
    .Y(_2864_));
 sky130_fd_sc_hd__nand2_1 _6503_ (.A(_2864_),
    .B(_2827_),
    .Y(_2865_));
 sky130_fd_sc_hd__nand3_1 _6504_ (.A(_2862_),
    .B(_2685_),
    .C(_2865_),
    .Y(_2866_));
 sky130_fd_sc_hd__nand2_1 _6505_ (.A(_2819_),
    .B(_2849_),
    .Y(_2867_));
 sky130_fd_sc_hd__nand2_1 _6506_ (.A(_2867_),
    .B(_2860_),
    .Y(_2868_));
 sky130_fd_sc_hd__inv_2 _6507_ (.A(_2860_),
    .Y(_2869_));
 sky130_fd_sc_hd__nand3_1 _6508_ (.A(_2819_),
    .B(_2849_),
    .C(_2869_),
    .Y(_2870_));
 sky130_fd_sc_hd__nand3_1 _6509_ (.A(_2868_),
    .B(_2701_),
    .C(_2870_),
    .Y(_2871_));
 sky130_fd_sc_hd__nand2_1 _6510_ (.A(_2866_),
    .B(_2871_),
    .Y(_2872_));
 sky130_fd_sc_hd__nand2_1 _6511_ (.A(_2872_),
    .B(_2923_),
    .Y(_2873_));
 sky130_fd_sc_hd__nand2_1 _6512_ (.A(_2833_),
    .B(_2846_),
    .Y(_2874_));
 sky130_fd_sc_hd__nand2_1 _6513_ (.A(_2873_),
    .B(_2874_),
    .Y(net25));
 sky130_fd_sc_hd__o21ai_1 _6514_ (.A1(_2858_),
    .A2(_2854_),
    .B1(_2855_),
    .Y(_2875_));
 sky130_fd_sc_hd__or2_1 _6515_ (.A(_2695_),
    .B(_2875_),
    .X(_2876_));
 sky130_fd_sc_hd__nand3_1 _6516_ (.A(_2870_),
    .B(_2701_),
    .C(_2876_),
    .Y(_2877_));
 sky130_fd_sc_hd__nor2_1 _6517_ (.A(_2737_),
    .B(_2695_),
    .Y(_2878_));
 sky130_fd_sc_hd__nor2_1 _6518_ (.A(_2701_),
    .B(_2876_),
    .Y(_2879_));
 sky130_fd_sc_hd__nand2_1 _6519_ (.A(_2865_),
    .B(_2879_),
    .Y(_2880_));
 sky130_fd_sc_hd__nand3_1 _6520_ (.A(_2877_),
    .B(_2878_),
    .C(_2880_),
    .Y(_2881_));
 sky130_fd_sc_hd__o21ai_2 _6521_ (.A1(_2832_),
    .A2(_2860_),
    .B1(_2881_),
    .Y(net26));
 sky130_fd_sc_hd__a2bb2o_1 _6522_ (.A1_N(_2875_),
    .A2_N(_2832_),
    .B1(_2685_),
    .B2(_2878_),
    .X(net27));
 sky130_fd_sc_hd__buf_1 _6523_ (.A(wb_clk_i),
    .X(_2882_));
 sky130_fd_sc_hd__buf_1 _6524_ (.A(clknet_1_1__leaf__2882_),
    .X(_2883_));
 sky130_fd_sc_hd__buf_1 _6525_ (.A(clknet_1_1__leaf__2883_),
    .X(_2884_));
 sky130_fd_sc_hd__inv_2 _6526__72 (.A(clknet_1_0__leaf__2884_),
    .Y(net106));
 sky130_fd_sc_hd__inv_2 _6527__73 (.A(clknet_1_1__leaf__2884_),
    .Y(net107));
 sky130_fd_sc_hd__inv_2 _6528__74 (.A(clknet_1_1__leaf__2884_),
    .Y(net108));
 sky130_fd_sc_hd__inv_2 _6529__75 (.A(clknet_1_1__leaf__2884_),
    .Y(net109));
 sky130_fd_sc_hd__inv_2 _6530__76 (.A(clknet_1_1__leaf__2884_),
    .Y(net110));
 sky130_fd_sc_hd__inv_2 _6531__77 (.A(clknet_1_0__leaf__2884_),
    .Y(net111));
 sky130_fd_sc_hd__inv_2 _6532__78 (.A(clknet_1_0__leaf__2884_),
    .Y(net112));
 sky130_fd_sc_hd__inv_2 _6533__79 (.A(clknet_1_0__leaf__2884_),
    .Y(net113));
 sky130_fd_sc_hd__inv_2 _6534__80 (.A(clknet_1_0__leaf__2884_),
    .Y(net114));
 sky130_fd_sc_hd__inv_2 _6535__81 (.A(clknet_1_1__leaf__2884_),
    .Y(net115));
 sky130_fd_sc_hd__buf_1 _6536_ (.A(clknet_1_1__leaf__2883_),
    .X(_2885_));
 sky130_fd_sc_hd__inv_2 _6537__82 (.A(clknet_1_0__leaf__2885_),
    .Y(net116));
 sky130_fd_sc_hd__inv_2 _6538__83 (.A(clknet_1_1__leaf__2885_),
    .Y(net117));
 sky130_fd_sc_hd__inv_2 _6539__84 (.A(clknet_1_1__leaf__2885_),
    .Y(net118));
 sky130_fd_sc_hd__inv_2 _6540__85 (.A(clknet_1_0__leaf__2885_),
    .Y(net119));
 sky130_fd_sc_hd__inv_2 _6541__86 (.A(clknet_1_0__leaf__2885_),
    .Y(net120));
 sky130_fd_sc_hd__inv_2 _6542__87 (.A(clknet_1_1__leaf__2885_),
    .Y(net121));
 sky130_fd_sc_hd__inv_2 _6543__88 (.A(clknet_1_1__leaf__2885_),
    .Y(net122));
 sky130_fd_sc_hd__inv_2 _6544__89 (.A(clknet_1_0__leaf__2885_),
    .Y(net123));
 sky130_fd_sc_hd__inv_2 _6545__90 (.A(clknet_1_0__leaf__2885_),
    .Y(net124));
 sky130_fd_sc_hd__inv_2 _6546__91 (.A(clknet_1_0__leaf__2885_),
    .Y(net125));
 sky130_fd_sc_hd__buf_1 _6547_ (.A(clknet_1_0__leaf__2883_),
    .X(_2886_));
 sky130_fd_sc_hd__inv_2 _6548__92 (.A(clknet_1_0__leaf__2886_),
    .Y(net126));
 sky130_fd_sc_hd__inv_2 _6549__93 (.A(clknet_1_1__leaf__2886_),
    .Y(net127));
 sky130_fd_sc_hd__inv_2 _6550__94 (.A(clknet_1_1__leaf__2886_),
    .Y(net128));
 sky130_fd_sc_hd__inv_2 _6551__95 (.A(clknet_1_1__leaf__2886_),
    .Y(net129));
 sky130_fd_sc_hd__inv_2 _6552__96 (.A(clknet_1_1__leaf__2886_),
    .Y(net130));
 sky130_fd_sc_hd__inv_2 _6553__97 (.A(clknet_1_1__leaf__2886_),
    .Y(net131));
 sky130_fd_sc_hd__inv_2 _6554__98 (.A(clknet_1_0__leaf__2886_),
    .Y(net132));
 sky130_fd_sc_hd__inv_2 _6555__99 (.A(clknet_1_0__leaf__2886_),
    .Y(net133));
 sky130_fd_sc_hd__inv_2 _6556__100 (.A(clknet_1_0__leaf__2886_),
    .Y(net134));
 sky130_fd_sc_hd__inv_2 _6557__101 (.A(clknet_1_0__leaf__2886_),
    .Y(net135));
 sky130_fd_sc_hd__buf_1 _6558_ (.A(clknet_1_0__leaf__2883_),
    .X(_2887_));
 sky130_fd_sc_hd__inv_2 _6559__102 (.A(clknet_1_0__leaf__2887_),
    .Y(net136));
 sky130_fd_sc_hd__inv_2 _6560__103 (.A(clknet_1_0__leaf__2887_),
    .Y(net137));
 sky130_fd_sc_hd__inv_2 _6561__104 (.A(clknet_1_1__leaf__2887_),
    .Y(net138));
 sky130_fd_sc_hd__inv_2 _6562__105 (.A(clknet_1_1__leaf__2887_),
    .Y(net139));
 sky130_fd_sc_hd__inv_2 _6563__106 (.A(clknet_1_1__leaf__2887_),
    .Y(net140));
 sky130_fd_sc_hd__inv_2 _6564__107 (.A(clknet_1_1__leaf__2887_),
    .Y(net141));
 sky130_fd_sc_hd__inv_2 _6565__108 (.A(clknet_1_0__leaf__2887_),
    .Y(net142));
 sky130_fd_sc_hd__inv_2 _6566__109 (.A(clknet_1_0__leaf__2887_),
    .Y(net143));
 sky130_fd_sc_hd__inv_2 _6567__110 (.A(clknet_1_1__leaf__2887_),
    .Y(net144));
 sky130_fd_sc_hd__inv_2 _6568__111 (.A(clknet_1_0__leaf__2887_),
    .Y(net145));
 sky130_fd_sc_hd__buf_1 _6569_ (.A(clknet_1_1__leaf__2883_),
    .X(_2888_));
 sky130_fd_sc_hd__inv_2 _6570__112 (.A(clknet_1_0__leaf__2888_),
    .Y(net146));
 sky130_fd_sc_hd__inv_2 _6571__113 (.A(clknet_1_0__leaf__2888_),
    .Y(net147));
 sky130_fd_sc_hd__inv_2 _6572__114 (.A(clknet_1_1__leaf__2888_),
    .Y(net148));
 sky130_fd_sc_hd__inv_2 _6573__115 (.A(clknet_1_0__leaf__2888_),
    .Y(net149));
 sky130_fd_sc_hd__inv_2 _6574__116 (.A(clknet_1_0__leaf__2888_),
    .Y(net150));
 sky130_fd_sc_hd__inv_2 _6575__117 (.A(clknet_1_1__leaf__2888_),
    .Y(net151));
 sky130_fd_sc_hd__inv_2 _6576__118 (.A(clknet_1_1__leaf__2888_),
    .Y(net152));
 sky130_fd_sc_hd__inv_2 _6577__119 (.A(clknet_1_1__leaf__2888_),
    .Y(net153));
 sky130_fd_sc_hd__inv_2 _6578__120 (.A(clknet_1_1__leaf__2888_),
    .Y(net154));
 sky130_fd_sc_hd__inv_2 _6579__121 (.A(clknet_1_1__leaf__2888_),
    .Y(net155));
 sky130_fd_sc_hd__buf_1 _6580_ (.A(clknet_1_1__leaf__2883_),
    .X(_2889_));
 sky130_fd_sc_hd__inv_2 _6581__122 (.A(clknet_1_0__leaf__2889_),
    .Y(net156));
 sky130_fd_sc_hd__inv_2 _6582__123 (.A(clknet_1_0__leaf__2889_),
    .Y(net157));
 sky130_fd_sc_hd__inv_2 _6583__124 (.A(clknet_1_0__leaf__2889_),
    .Y(net158));
 sky130_fd_sc_hd__inv_2 _6584__125 (.A(clknet_1_0__leaf__2889_),
    .Y(net159));
 sky130_fd_sc_hd__inv_2 _6585__126 (.A(clknet_1_0__leaf__2889_),
    .Y(net160));
 sky130_fd_sc_hd__inv_2 _6586__127 (.A(clknet_1_1__leaf__2889_),
    .Y(net161));
 sky130_fd_sc_hd__inv_2 _6587__128 (.A(clknet_1_1__leaf__2889_),
    .Y(net162));
 sky130_fd_sc_hd__inv_2 _6588__129 (.A(clknet_1_1__leaf__2889_),
    .Y(net163));
 sky130_fd_sc_hd__inv_2 _6589__130 (.A(clknet_1_1__leaf__2889_),
    .Y(net164));
 sky130_fd_sc_hd__inv_2 _6590__131 (.A(clknet_1_1__leaf__2889_),
    .Y(net165));
 sky130_fd_sc_hd__buf_1 _6591_ (.A(clknet_1_1__leaf__2883_),
    .X(_2890_));
 sky130_fd_sc_hd__inv_2 _6592__132 (.A(clknet_1_1__leaf__2890_),
    .Y(net166));
 sky130_fd_sc_hd__inv_2 _6593__133 (.A(clknet_1_0__leaf__2890_),
    .Y(net167));
 sky130_fd_sc_hd__inv_2 _6594__134 (.A(clknet_1_1__leaf__2890_),
    .Y(net168));
 sky130_fd_sc_hd__inv_2 _6595__135 (.A(clknet_1_0__leaf__2890_),
    .Y(net169));
 sky130_fd_sc_hd__inv_2 _6596__136 (.A(clknet_1_1__leaf__2890_),
    .Y(net170));
 sky130_fd_sc_hd__inv_2 _6597__137 (.A(clknet_1_1__leaf__2890_),
    .Y(net171));
 sky130_fd_sc_hd__inv_2 _6598__138 (.A(clknet_1_0__leaf__2890_),
    .Y(net172));
 sky130_fd_sc_hd__inv_2 _6599__139 (.A(clknet_1_0__leaf__2890_),
    .Y(net173));
 sky130_fd_sc_hd__inv_2 _6600__140 (.A(clknet_1_0__leaf__2890_),
    .Y(net174));
 sky130_fd_sc_hd__inv_2 _6601__141 (.A(clknet_1_0__leaf__2890_),
    .Y(net175));
 sky130_fd_sc_hd__buf_1 _6602_ (.A(clknet_1_1__leaf__2883_),
    .X(_2891_));
 sky130_fd_sc_hd__inv_2 _6603__142 (.A(clknet_1_0__leaf__2891_),
    .Y(net176));
 sky130_fd_sc_hd__inv_2 _6604__143 (.A(clknet_1_1__leaf__2891_),
    .Y(net177));
 sky130_fd_sc_hd__inv_2 _6605__144 (.A(clknet_1_1__leaf__2891_),
    .Y(net178));
 sky130_fd_sc_hd__inv_2 _6606__145 (.A(clknet_1_1__leaf__2891_),
    .Y(net179));
 sky130_fd_sc_hd__inv_2 _6607__146 (.A(clknet_1_1__leaf__2891_),
    .Y(net180));
 sky130_fd_sc_hd__inv_2 _6608__147 (.A(clknet_1_0__leaf__2891_),
    .Y(net181));
 sky130_fd_sc_hd__inv_2 _6609__148 (.A(clknet_1_0__leaf__2891_),
    .Y(net182));
 sky130_fd_sc_hd__inv_2 _6610__149 (.A(clknet_1_0__leaf__2891_),
    .Y(net183));
 sky130_fd_sc_hd__inv_2 _6611__150 (.A(clknet_1_0__leaf__2891_),
    .Y(net184));
 sky130_fd_sc_hd__inv_2 _6612__151 (.A(clknet_1_1__leaf__2891_),
    .Y(net185));
 sky130_fd_sc_hd__buf_1 _6613_ (.A(clknet_1_0__leaf__2883_),
    .X(_2892_));
 sky130_fd_sc_hd__inv_2 _6614__152 (.A(clknet_1_1__leaf__2892_),
    .Y(net186));
 sky130_fd_sc_hd__inv_2 _6615__153 (.A(clknet_1_1__leaf__2892_),
    .Y(net187));
 sky130_fd_sc_hd__inv_2 _6616__154 (.A(clknet_1_1__leaf__2892_),
    .Y(net188));
 sky130_fd_sc_hd__inv_2 _6617__155 (.A(clknet_1_1__leaf__2892_),
    .Y(net189));
 sky130_fd_sc_hd__inv_2 _6618__156 (.A(clknet_1_1__leaf__2892_),
    .Y(net190));
 sky130_fd_sc_hd__inv_2 _6619__157 (.A(clknet_1_1__leaf__2892_),
    .Y(net191));
 sky130_fd_sc_hd__inv_2 _6620__158 (.A(clknet_1_0__leaf__2892_),
    .Y(net192));
 sky130_fd_sc_hd__inv_2 _6621__159 (.A(clknet_1_0__leaf__2892_),
    .Y(net193));
 sky130_fd_sc_hd__inv_2 _6622__160 (.A(clknet_1_0__leaf__2892_),
    .Y(net194));
 sky130_fd_sc_hd__inv_2 _6623__161 (.A(clknet_1_0__leaf__2892_),
    .Y(net195));
 sky130_fd_sc_hd__buf_1 _6624_ (.A(clknet_1_1__leaf__2882_),
    .X(_2893_));
 sky130_fd_sc_hd__inv_2 _6625__2 (.A(clknet_1_1__leaf__2893_),
    .Y(net36));
 sky130_fd_sc_hd__inv_2 _6626__3 (.A(clknet_1_1__leaf__2893_),
    .Y(net37));
 sky130_fd_sc_hd__inv_2 _6627__4 (.A(clknet_1_0__leaf__2893_),
    .Y(net38));
 sky130_fd_sc_hd__inv_2 _6628__5 (.A(clknet_1_0__leaf__2893_),
    .Y(net39));
 sky130_fd_sc_hd__inv_2 _6629__6 (.A(clknet_1_0__leaf__2893_),
    .Y(net40));
 sky130_fd_sc_hd__inv_2 _6630__7 (.A(clknet_1_0__leaf__2893_),
    .Y(net41));
 sky130_fd_sc_hd__inv_2 _6631__8 (.A(clknet_1_0__leaf__2893_),
    .Y(net42));
 sky130_fd_sc_hd__inv_2 _6632__9 (.A(clknet_1_1__leaf__2893_),
    .Y(net43));
 sky130_fd_sc_hd__inv_2 _6633__10 (.A(clknet_1_1__leaf__2893_),
    .Y(net44));
 sky130_fd_sc_hd__inv_2 _6634__11 (.A(clknet_1_1__leaf__2893_),
    .Y(net45));
 sky130_fd_sc_hd__buf_1 _6635_ (.A(clknet_1_1__leaf__2882_),
    .X(_2894_));
 sky130_fd_sc_hd__inv_2 _6636__12 (.A(clknet_1_1__leaf__2894_),
    .Y(net46));
 sky130_fd_sc_hd__inv_2 _6637__13 (.A(clknet_1_1__leaf__2894_),
    .Y(net47));
 sky130_fd_sc_hd__inv_2 _6638__14 (.A(clknet_1_1__leaf__2894_),
    .Y(net48));
 sky130_fd_sc_hd__inv_2 _6639__15 (.A(clknet_1_1__leaf__2894_),
    .Y(net49));
 sky130_fd_sc_hd__inv_2 _6640__16 (.A(clknet_1_0__leaf__2894_),
    .Y(net50));
 sky130_fd_sc_hd__inv_2 _6641__17 (.A(clknet_1_0__leaf__2894_),
    .Y(net51));
 sky130_fd_sc_hd__inv_2 _6642__18 (.A(clknet_1_1__leaf__2894_),
    .Y(net52));
 sky130_fd_sc_hd__inv_2 _6643__19 (.A(clknet_1_0__leaf__2894_),
    .Y(net53));
 sky130_fd_sc_hd__inv_2 _6644__20 (.A(clknet_1_0__leaf__2894_),
    .Y(net54));
 sky130_fd_sc_hd__inv_2 _6645__21 (.A(clknet_1_0__leaf__2894_),
    .Y(net55));
 sky130_fd_sc_hd__buf_1 _6646_ (.A(clknet_1_0__leaf__2882_),
    .X(_2895_));
 sky130_fd_sc_hd__inv_2 _6647__22 (.A(clknet_1_1__leaf__2895_),
    .Y(net56));
 sky130_fd_sc_hd__inv_2 _6648__23 (.A(clknet_1_0__leaf__2895_),
    .Y(net57));
 sky130_fd_sc_hd__inv_2 _6649__24 (.A(clknet_1_1__leaf__2895_),
    .Y(net58));
 sky130_fd_sc_hd__inv_2 _6650__25 (.A(clknet_1_1__leaf__2895_),
    .Y(net59));
 sky130_fd_sc_hd__inv_2 _6651__26 (.A(clknet_1_1__leaf__2895_),
    .Y(net60));
 sky130_fd_sc_hd__inv_2 _6652__27 (.A(clknet_1_1__leaf__2895_),
    .Y(net61));
 sky130_fd_sc_hd__inv_2 _6653__28 (.A(clknet_1_0__leaf__2895_),
    .Y(net62));
 sky130_fd_sc_hd__inv_2 _6654__29 (.A(clknet_1_0__leaf__2895_),
    .Y(net63));
 sky130_fd_sc_hd__inv_2 _6655__30 (.A(clknet_1_0__leaf__2895_),
    .Y(net64));
 sky130_fd_sc_hd__inv_2 _6656__31 (.A(clknet_1_0__leaf__2895_),
    .Y(net65));
 sky130_fd_sc_hd__buf_1 _6657_ (.A(clknet_1_1__leaf__2882_),
    .X(_2896_));
 sky130_fd_sc_hd__inv_2 _6658__32 (.A(clknet_1_0__leaf__2896_),
    .Y(net66));
 sky130_fd_sc_hd__inv_2 _6659__33 (.A(clknet_1_1__leaf__2896_),
    .Y(net67));
 sky130_fd_sc_hd__inv_2 _6660__34 (.A(clknet_1_0__leaf__2896_),
    .Y(net68));
 sky130_fd_sc_hd__inv_2 _6661__35 (.A(clknet_1_0__leaf__2896_),
    .Y(net69));
 sky130_fd_sc_hd__inv_2 _6662__36 (.A(clknet_1_0__leaf__2896_),
    .Y(net70));
 sky130_fd_sc_hd__inv_2 _6663__37 (.A(clknet_1_1__leaf__2896_),
    .Y(net71));
 sky130_fd_sc_hd__inv_2 _6664__38 (.A(clknet_1_1__leaf__2896_),
    .Y(net72));
 sky130_fd_sc_hd__inv_2 _6665__39 (.A(clknet_1_0__leaf__2896_),
    .Y(net73));
 sky130_fd_sc_hd__inv_2 _6666__40 (.A(clknet_1_1__leaf__2896_),
    .Y(net74));
 sky130_fd_sc_hd__inv_2 _6667__41 (.A(clknet_1_1__leaf__2896_),
    .Y(net75));
 sky130_fd_sc_hd__buf_1 _6668_ (.A(clknet_1_0__leaf__2882_),
    .X(_2897_));
 sky130_fd_sc_hd__inv_2 _6669__42 (.A(clknet_1_1__leaf__2897_),
    .Y(net76));
 sky130_fd_sc_hd__inv_2 _6670__43 (.A(clknet_1_1__leaf__2897_),
    .Y(net77));
 sky130_fd_sc_hd__inv_2 _6671__44 (.A(clknet_1_0__leaf__2897_),
    .Y(net78));
 sky130_fd_sc_hd__inv_2 _6672__45 (.A(clknet_1_0__leaf__2897_),
    .Y(net79));
 sky130_fd_sc_hd__inv_2 _6673__46 (.A(clknet_1_0__leaf__2897_),
    .Y(net80));
 sky130_fd_sc_hd__inv_2 _6674__47 (.A(clknet_1_1__leaf__2897_),
    .Y(net81));
 sky130_fd_sc_hd__inv_2 _6675__48 (.A(clknet_1_1__leaf__2897_),
    .Y(net82));
 sky130_fd_sc_hd__inv_2 _6676__49 (.A(clknet_1_1__leaf__2897_),
    .Y(net83));
 sky130_fd_sc_hd__inv_2 _6677__50 (.A(clknet_1_0__leaf__2897_),
    .Y(net84));
 sky130_fd_sc_hd__inv_2 _6678__51 (.A(clknet_1_1__leaf__2897_),
    .Y(net85));
 sky130_fd_sc_hd__buf_1 _6679_ (.A(clknet_1_0__leaf__2882_),
    .X(_2898_));
 sky130_fd_sc_hd__inv_2 _6680__52 (.A(clknet_1_1__leaf__2898_),
    .Y(net86));
 sky130_fd_sc_hd__inv_2 _6681__53 (.A(clknet_1_1__leaf__2898_),
    .Y(net87));
 sky130_fd_sc_hd__inv_2 _6682__54 (.A(clknet_1_1__leaf__2898_),
    .Y(net88));
 sky130_fd_sc_hd__inv_2 _6683__55 (.A(clknet_1_1__leaf__2898_),
    .Y(net89));
 sky130_fd_sc_hd__inv_2 _6684__56 (.A(clknet_1_1__leaf__2898_),
    .Y(net90));
 sky130_fd_sc_hd__inv_2 _6685__57 (.A(clknet_1_0__leaf__2898_),
    .Y(net91));
 sky130_fd_sc_hd__inv_2 _6686__58 (.A(clknet_1_0__leaf__2898_),
    .Y(net92));
 sky130_fd_sc_hd__inv_2 _6687__59 (.A(clknet_1_0__leaf__2898_),
    .Y(net93));
 sky130_fd_sc_hd__inv_2 _6688__60 (.A(clknet_1_0__leaf__2898_),
    .Y(net94));
 sky130_fd_sc_hd__inv_2 _6689__61 (.A(clknet_1_0__leaf__2898_),
    .Y(net95));
 sky130_fd_sc_hd__buf_1 _6690_ (.A(clknet_1_0__leaf__2882_),
    .X(_2899_));
 sky130_fd_sc_hd__inv_2 _6691__62 (.A(clknet_1_1__leaf__2899_),
    .Y(net96));
 sky130_fd_sc_hd__inv_2 _6692__63 (.A(clknet_1_1__leaf__2899_),
    .Y(net97));
 sky130_fd_sc_hd__inv_2 _6693__64 (.A(clknet_1_1__leaf__2899_),
    .Y(net98));
 sky130_fd_sc_hd__inv_2 _6694__65 (.A(clknet_1_0__leaf__2899_),
    .Y(net99));
 sky130_fd_sc_hd__inv_2 _6695__66 (.A(clknet_1_0__leaf__2899_),
    .Y(net100));
 sky130_fd_sc_hd__inv_2 _6696__67 (.A(clknet_1_0__leaf__2899_),
    .Y(net101));
 sky130_fd_sc_hd__inv_2 _6697__68 (.A(clknet_1_0__leaf__2899_),
    .Y(net102));
 sky130_fd_sc_hd__inv_2 _6698__69 (.A(clknet_1_0__leaf__2899_),
    .Y(net103));
 sky130_fd_sc_hd__inv_2 _6699__70 (.A(clknet_1_1__leaf__2899_),
    .Y(net104));
 sky130_fd_sc_hd__inv_2 _6700__71 (.A(clknet_1_1__leaf__2899_),
    .Y(net105));
 sky130_fd_sc_hd__inv_2 _6701__1 (.A(clknet_1_0__leaf__2883_),
    .Y(net35));
 sky130_fd_sc_hd__dfxtp_1 _6702_ (.CLK(net106),
    .D(_0161_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[95] ));
 sky130_fd_sc_hd__dfxtp_1 _6703_ (.CLK(net107),
    .D(_0162_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[94] ));
 sky130_fd_sc_hd__dfxtp_1 _6704_ (.CLK(net108),
    .D(_0163_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[93] ));
 sky130_fd_sc_hd__dfxtp_1 _6705_ (.CLK(net109),
    .D(_0164_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[92] ));
 sky130_fd_sc_hd__dfxtp_1 _6706_ (.CLK(net110),
    .D(_0165_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[91] ));
 sky130_fd_sc_hd__dfxtp_1 _6707_ (.CLK(net111),
    .D(_0166_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[90] ));
 sky130_fd_sc_hd__dfxtp_1 _6708_ (.CLK(net112),
    .D(_0167_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[89] ));
 sky130_fd_sc_hd__dfxtp_1 _6709_ (.CLK(net113),
    .D(_0168_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[88] ));
 sky130_fd_sc_hd__dfxtp_1 _6710_ (.CLK(net114),
    .D(_0169_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[87] ));
 sky130_fd_sc_hd__dfxtp_1 _6711_ (.CLK(net115),
    .D(_0170_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[86] ));
 sky130_fd_sc_hd__dfxtp_1 _6712_ (.CLK(net116),
    .D(_0171_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[85] ));
 sky130_fd_sc_hd__dfxtp_1 _6713_ (.CLK(net117),
    .D(_0172_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[84] ));
 sky130_fd_sc_hd__dfxtp_1 _6714_ (.CLK(net118),
    .D(_0173_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[83] ));
 sky130_fd_sc_hd__dfxtp_1 _6715_ (.CLK(net119),
    .D(_0174_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[82] ));
 sky130_fd_sc_hd__dfxtp_1 _6716_ (.CLK(net120),
    .D(_0175_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[81] ));
 sky130_fd_sc_hd__dfxtp_1 _6717_ (.CLK(net121),
    .D(_0176_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[80] ));
 sky130_fd_sc_hd__dfxtp_2 _6718_ (.CLK(net122),
    .D(_0177_),
    .Q(\egd_top.BitStream_buffer.pc_previous[0] ));
 sky130_fd_sc_hd__dfxtp_1 _6719_ (.CLK(net123),
    .D(_0178_),
    .Q(\egd_top.BitStream_buffer.pc_previous[1] ));
 sky130_fd_sc_hd__dfxtp_1 _6720_ (.CLK(net124),
    .D(_0179_),
    .Q(\egd_top.BitStream_buffer.pc_previous[2] ));
 sky130_fd_sc_hd__dfxtp_1 _6721_ (.CLK(net125),
    .D(_0180_),
    .Q(\egd_top.BitStream_buffer.pc_previous[3] ));
 sky130_fd_sc_hd__dfxtp_1 _6722_ (.CLK(net126),
    .D(_0181_),
    .Q(\egd_top.BitStream_buffer.pc_previous[4] ));
 sky130_fd_sc_hd__dfxtp_1 _6723_ (.CLK(net127),
    .D(_0182_),
    .Q(\egd_top.BitStream_buffer.pc_previous[5] ));
 sky130_fd_sc_hd__dfxtp_2 _6724_ (.CLK(net128),
    .D(_0183_),
    .Q(\egd_top.BitStream_buffer.pc_previous[6] ));
 sky130_fd_sc_hd__dfxtp_1 _6725_ (.CLK(net129),
    .D(_0184_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[111] ));
 sky130_fd_sc_hd__dfxtp_1 _6726_ (.CLK(net130),
    .D(_0185_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[110] ));
 sky130_fd_sc_hd__dfxtp_1 _6727_ (.CLK(net131),
    .D(_0186_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[109] ));
 sky130_fd_sc_hd__dfxtp_1 _6728_ (.CLK(net132),
    .D(_0187_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[108] ));
 sky130_fd_sc_hd__dfxtp_1 _6729_ (.CLK(net133),
    .D(_0188_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[107] ));
 sky130_fd_sc_hd__dfxtp_1 _6730_ (.CLK(net134),
    .D(_0189_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[106] ));
 sky130_fd_sc_hd__dfxtp_1 _6731_ (.CLK(net135),
    .D(_0190_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[105] ));
 sky130_fd_sc_hd__dfxtp_1 _6732_ (.CLK(net136),
    .D(_0191_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[104] ));
 sky130_fd_sc_hd__dfxtp_1 _6733_ (.CLK(net137),
    .D(_0192_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[103] ));
 sky130_fd_sc_hd__dfxtp_1 _6734_ (.CLK(net138),
    .D(_0193_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[102] ));
 sky130_fd_sc_hd__dfxtp_1 _6735_ (.CLK(net139),
    .D(_0194_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[101] ));
 sky130_fd_sc_hd__dfxtp_1 _6736_ (.CLK(net140),
    .D(_0195_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[100] ));
 sky130_fd_sc_hd__dfxtp_1 _6737_ (.CLK(net141),
    .D(_0196_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[99] ));
 sky130_fd_sc_hd__dfxtp_1 _6738_ (.CLK(net142),
    .D(_0197_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[98] ));
 sky130_fd_sc_hd__dfxtp_1 _6739_ (.CLK(net143),
    .D(_0198_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[97] ));
 sky130_fd_sc_hd__dfxtp_1 _6740_ (.CLK(net144),
    .D(_0199_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[96] ));
 sky130_fd_sc_hd__dfxtp_1 _6741_ (.CLK(net145),
    .D(_0200_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[79] ));
 sky130_fd_sc_hd__dfxtp_1 _6742_ (.CLK(net146),
    .D(_0201_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[78] ));
 sky130_fd_sc_hd__dfxtp_1 _6743_ (.CLK(net147),
    .D(_0202_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[77] ));
 sky130_fd_sc_hd__dfxtp_1 _6744_ (.CLK(net148),
    .D(_0203_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[76] ));
 sky130_fd_sc_hd__dfxtp_1 _6745_ (.CLK(net149),
    .D(_0204_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[75] ));
 sky130_fd_sc_hd__dfxtp_1 _6746_ (.CLK(net150),
    .D(_0205_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[74] ));
 sky130_fd_sc_hd__dfxtp_1 _6747_ (.CLK(net151),
    .D(_0206_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[73] ));
 sky130_fd_sc_hd__dfxtp_1 _6748_ (.CLK(net152),
    .D(_0207_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[72] ));
 sky130_fd_sc_hd__dfxtp_1 _6749_ (.CLK(net153),
    .D(_0208_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[71] ));
 sky130_fd_sc_hd__dfxtp_1 _6750_ (.CLK(net154),
    .D(_0209_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[70] ));
 sky130_fd_sc_hd__dfxtp_1 _6751_ (.CLK(net155),
    .D(_0210_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[69] ));
 sky130_fd_sc_hd__dfxtp_1 _6752_ (.CLK(net156),
    .D(_0211_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[68] ));
 sky130_fd_sc_hd__dfxtp_1 _6753_ (.CLK(net157),
    .D(_0212_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[67] ));
 sky130_fd_sc_hd__dfxtp_1 _6754_ (.CLK(net158),
    .D(_0213_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[66] ));
 sky130_fd_sc_hd__dfxtp_1 _6755_ (.CLK(net159),
    .D(_0214_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[65] ));
 sky130_fd_sc_hd__dfxtp_1 _6756_ (.CLK(net160),
    .D(_0215_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[64] ));
 sky130_fd_sc_hd__dfxtp_1 _6757_ (.CLK(net161),
    .D(_0216_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[63] ));
 sky130_fd_sc_hd__dfxtp_1 _6758_ (.CLK(net162),
    .D(_0217_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[62] ));
 sky130_fd_sc_hd__dfxtp_1 _6759_ (.CLK(net163),
    .D(_0218_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[61] ));
 sky130_fd_sc_hd__dfxtp_1 _6760_ (.CLK(net164),
    .D(_0219_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[60] ));
 sky130_fd_sc_hd__dfxtp_1 _6761_ (.CLK(net165),
    .D(_0220_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[59] ));
 sky130_fd_sc_hd__dfxtp_1 _6762_ (.CLK(net166),
    .D(_0221_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[58] ));
 sky130_fd_sc_hd__dfxtp_1 _6763_ (.CLK(net167),
    .D(_0222_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[57] ));
 sky130_fd_sc_hd__dfxtp_1 _6764_ (.CLK(net168),
    .D(_0223_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[56] ));
 sky130_fd_sc_hd__dfxtp_1 _6765_ (.CLK(net169),
    .D(_0224_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[55] ));
 sky130_fd_sc_hd__dfxtp_1 _6766_ (.CLK(net170),
    .D(_0225_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[54] ));
 sky130_fd_sc_hd__dfxtp_1 _6767_ (.CLK(net171),
    .D(_0226_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[53] ));
 sky130_fd_sc_hd__dfxtp_1 _6768_ (.CLK(net172),
    .D(_0227_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[52] ));
 sky130_fd_sc_hd__dfxtp_1 _6769_ (.CLK(net173),
    .D(_0228_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[51] ));
 sky130_fd_sc_hd__dfxtp_1 _6770_ (.CLK(net174),
    .D(_0229_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[50] ));
 sky130_fd_sc_hd__dfxtp_1 _6771_ (.CLK(net175),
    .D(_0230_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[49] ));
 sky130_fd_sc_hd__dfxtp_1 _6772_ (.CLK(net176),
    .D(_0231_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[48] ));
 sky130_fd_sc_hd__dfxtp_1 _6773_ (.CLK(net177),
    .D(_0232_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[47] ));
 sky130_fd_sc_hd__dfxtp_2 _6774_ (.CLK(net178),
    .D(_0233_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[46] ));
 sky130_fd_sc_hd__dfxtp_1 _6775_ (.CLK(net179),
    .D(_0234_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[45] ));
 sky130_fd_sc_hd__dfxtp_1 _6776_ (.CLK(net180),
    .D(_0235_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[44] ));
 sky130_fd_sc_hd__dfxtp_1 _6777_ (.CLK(net181),
    .D(_0236_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[43] ));
 sky130_fd_sc_hd__dfxtp_1 _6778_ (.CLK(net182),
    .D(_0237_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[42] ));
 sky130_fd_sc_hd__dfxtp_1 _6779_ (.CLK(net183),
    .D(_0238_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[41] ));
 sky130_fd_sc_hd__dfxtp_1 _6780_ (.CLK(net184),
    .D(_0239_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[40] ));
 sky130_fd_sc_hd__dfxtp_1 _6781_ (.CLK(net185),
    .D(_0240_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[39] ));
 sky130_fd_sc_hd__dfxtp_1 _6782_ (.CLK(net186),
    .D(_0241_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[38] ));
 sky130_fd_sc_hd__dfxtp_1 _6783_ (.CLK(net187),
    .D(_0242_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[37] ));
 sky130_fd_sc_hd__dfxtp_1 _6784_ (.CLK(net188),
    .D(_0243_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[36] ));
 sky130_fd_sc_hd__dfxtp_1 _6785_ (.CLK(net189),
    .D(_0244_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[35] ));
 sky130_fd_sc_hd__dfxtp_2 _6786_ (.CLK(net190),
    .D(_0245_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[34] ));
 sky130_fd_sc_hd__dfxtp_1 _6787_ (.CLK(net191),
    .D(_0246_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[33] ));
 sky130_fd_sc_hd__dfxtp_4 _6788_ (.CLK(net192),
    .D(_0247_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[32] ));
 sky130_fd_sc_hd__dfxtp_1 _6789_ (.CLK(net193),
    .D(_0248_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[31] ));
 sky130_fd_sc_hd__dfxtp_1 _6790_ (.CLK(net194),
    .D(_0249_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[30] ));
 sky130_fd_sc_hd__dfxtp_2 _6791_ (.CLK(net195),
    .D(_0250_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[29] ));
 sky130_fd_sc_hd__dfxtp_4 _6792_ (.CLK(net36),
    .D(_0251_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[28] ));
 sky130_fd_sc_hd__dfxtp_2 _6793_ (.CLK(net37),
    .D(_0252_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[27] ));
 sky130_fd_sc_hd__dfxtp_1 _6794_ (.CLK(net38),
    .D(_0253_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[26] ));
 sky130_fd_sc_hd__dfxtp_1 _6795_ (.CLK(net39),
    .D(_0254_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[25] ));
 sky130_fd_sc_hd__dfxtp_1 _6796_ (.CLK(net40),
    .D(_0255_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[24] ));
 sky130_fd_sc_hd__dfxtp_1 _6797_ (.CLK(net41),
    .D(_0256_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[23] ));
 sky130_fd_sc_hd__dfxtp_1 _6798_ (.CLK(net42),
    .D(_0257_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[22] ));
 sky130_fd_sc_hd__dfxtp_1 _6799_ (.CLK(net43),
    .D(_0258_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[21] ));
 sky130_fd_sc_hd__dfxtp_1 _6800_ (.CLK(net44),
    .D(_0259_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[20] ));
 sky130_fd_sc_hd__dfxtp_1 _6801_ (.CLK(net45),
    .D(_0260_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[19] ));
 sky130_fd_sc_hd__dfxtp_1 _6802_ (.CLK(net46),
    .D(_0261_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[18] ));
 sky130_fd_sc_hd__dfxtp_4 _6803_ (.CLK(net47),
    .D(_0262_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[17] ));
 sky130_fd_sc_hd__dfxtp_2 _6804_ (.CLK(net48),
    .D(_0263_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[16] ));
 sky130_fd_sc_hd__dfxtp_2 _6805_ (.CLK(net49),
    .D(_0264_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[15] ));
 sky130_fd_sc_hd__dfxtp_2 _6806_ (.CLK(net50),
    .D(_0265_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[14] ));
 sky130_fd_sc_hd__dfxtp_2 _6807_ (.CLK(net51),
    .D(_0266_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[13] ));
 sky130_fd_sc_hd__dfxtp_2 _6808_ (.CLK(net52),
    .D(_0267_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[12] ));
 sky130_fd_sc_hd__dfxtp_2 _6809_ (.CLK(net53),
    .D(_0268_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[11] ));
 sky130_fd_sc_hd__dfxtp_1 _6810_ (.CLK(net54),
    .D(_0269_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[10] ));
 sky130_fd_sc_hd__dfxtp_1 _6811_ (.CLK(net55),
    .D(_0270_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[9] ));
 sky130_fd_sc_hd__dfxtp_1 _6812_ (.CLK(net56),
    .D(_0271_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[8] ));
 sky130_fd_sc_hd__dfxtp_1 _6813_ (.CLK(net57),
    .D(_0272_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[7] ));
 sky130_fd_sc_hd__dfxtp_1 _6814_ (.CLK(net58),
    .D(_0273_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[6] ));
 sky130_fd_sc_hd__dfxtp_1 _6815_ (.CLK(net59),
    .D(_0274_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[5] ));
 sky130_fd_sc_hd__dfxtp_1 _6816_ (.CLK(net60),
    .D(_0275_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[4] ));
 sky130_fd_sc_hd__dfxtp_1 _6817_ (.CLK(net61),
    .D(_0276_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[3] ));
 sky130_fd_sc_hd__dfxtp_1 _6818_ (.CLK(net62),
    .D(_0277_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[2] ));
 sky130_fd_sc_hd__dfxtp_1 _6819_ (.CLK(net63),
    .D(_0278_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[1] ));
 sky130_fd_sc_hd__dfxtp_1 _6820_ (.CLK(net64),
    .D(_0279_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _6821_ (.CLK(net65),
    .D(_0280_),
    .Q(\egd_top.BitStream_buffer.buffer_index[4] ));
 sky130_fd_sc_hd__dfxtp_1 _6822_ (.CLK(net66),
    .D(_0281_),
    .Q(\egd_top.BitStream_buffer.buffer_index[5] ));
 sky130_fd_sc_hd__dfxtp_1 _6823_ (.CLK(net67),
    .D(_0282_),
    .Q(\egd_top.BitStream_buffer.buffer_index[6] ));
 sky130_fd_sc_hd__dfxtp_1 _6824_ (.CLK(net68),
    .D(_0283_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[1] ));
 sky130_fd_sc_hd__dfxtp_1 _6825_ (.CLK(net69),
    .D(_0284_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[2] ));
 sky130_fd_sc_hd__dfxtp_1 _6826_ (.CLK(net70),
    .D(_0285_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[3] ));
 sky130_fd_sc_hd__dfxtp_1 _6827_ (.CLK(net71),
    .D(_0286_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[4] ));
 sky130_fd_sc_hd__dfxtp_2 _6828_ (.CLK(net72),
    .D(_0287_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[5] ));
 sky130_fd_sc_hd__dfxtp_2 _6829_ (.CLK(net73),
    .D(_0288_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[6] ));
 sky130_fd_sc_hd__dfxtp_2 _6830_ (.CLK(net74),
    .D(_0289_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[7] ));
 sky130_fd_sc_hd__dfxtp_1 _6831_ (.CLK(net75),
    .D(_0290_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[8] ));
 sky130_fd_sc_hd__dfxtp_2 _6832_ (.CLK(net76),
    .D(_0291_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[9] ));
 sky130_fd_sc_hd__dfxtp_2 _6833_ (.CLK(net77),
    .D(_0292_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[10] ));
 sky130_fd_sc_hd__dfxtp_2 _6834_ (.CLK(net78),
    .D(_0293_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[11] ));
 sky130_fd_sc_hd__dfxtp_2 _6835_ (.CLK(net79),
    .D(_0294_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[12] ));
 sky130_fd_sc_hd__dfxtp_1 _6836_ (.CLK(net80),
    .D(_0295_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[13] ));
 sky130_fd_sc_hd__dfxtp_1 _6837_ (.CLK(net81),
    .D(_0296_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[14] ));
 sky130_fd_sc_hd__dfxtp_1 _6838_ (.CLK(net82),
    .D(_0297_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[15] ));
 sky130_fd_sc_hd__dfxtp_1 _6839_ (.CLK(net83),
    .D(_0298_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[127] ));
 sky130_fd_sc_hd__dfxtp_2 _6840_ (.CLK(net84),
    .D(_0299_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[126] ));
 sky130_fd_sc_hd__dfxtp_2 _6841_ (.CLK(net85),
    .D(_0300_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[125] ));
 sky130_fd_sc_hd__dfxtp_2 _6842_ (.CLK(net86),
    .D(_0301_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[124] ));
 sky130_fd_sc_hd__dfxtp_2 _6843_ (.CLK(net87),
    .D(_0302_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[123] ));
 sky130_fd_sc_hd__dfxtp_1 _6844_ (.CLK(net88),
    .D(_0303_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[122] ));
 sky130_fd_sc_hd__dfxtp_2 _6845_ (.CLK(net89),
    .D(_0304_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[121] ));
 sky130_fd_sc_hd__dfxtp_2 _6846_ (.CLK(net90),
    .D(_0305_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[120] ));
 sky130_fd_sc_hd__dfxtp_1 _6847_ (.CLK(net91),
    .D(_0306_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[119] ));
 sky130_fd_sc_hd__dfxtp_2 _6848_ (.CLK(net92),
    .D(_0307_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[118] ));
 sky130_fd_sc_hd__dfxtp_1 _6849_ (.CLK(net93),
    .D(_0308_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[117] ));
 sky130_fd_sc_hd__dfxtp_1 _6850_ (.CLK(net94),
    .D(_0309_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[116] ));
 sky130_fd_sc_hd__dfxtp_1 _6851_ (.CLK(net95),
    .D(_0310_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[115] ));
 sky130_fd_sc_hd__dfxtp_1 _6852_ (.CLK(net96),
    .D(_0311_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[114] ));
 sky130_fd_sc_hd__dfxtp_1 _6853_ (.CLK(net97),
    .D(_0312_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[113] ));
 sky130_fd_sc_hd__dfxtp_1 _6854_ (.CLK(net98),
    .D(_0313_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[112] ));
 sky130_fd_sc_hd__dfxtp_1 _6855_ (.CLK(net99),
    .D(_0314_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_valid_n ));
 sky130_fd_sc_hd__dfxtp_2 _6856_ (.CLK(net100),
    .D(_0315_),
    .Q(net28));
 sky130_fd_sc_hd__dfxtp_2 _6857_ (.CLK(net101),
    .D(_0316_),
    .Q(net29));
 sky130_fd_sc_hd__dfxtp_4 _6858_ (.CLK(net102),
    .D(_0317_),
    .Q(net30));
 sky130_fd_sc_hd__dfxtp_2 _6859_ (.CLK(net103),
    .D(_0318_),
    .Q(net31));
 sky130_fd_sc_hd__dfxtp_2 _6860_ (.CLK(net104),
    .D(_0319_),
    .Q(net32));
 sky130_fd_sc_hd__dfxtp_2 _6861_ (.CLK(net105),
    .D(_0320_),
    .Q(net33));
 sky130_fd_sc_hd__dfxtp_4 _6862_ (.CLK(net35),
    .D(_0321_),
    .Q(net34));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2882_ (.A(_2882_),
    .X(clknet_0__2882_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2883_ (.A(_2883_),
    .X(clknet_0__2883_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2884_ (.A(_2884_),
    .X(clknet_0__2884_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2885_ (.A(_2885_),
    .X(clknet_0__2885_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2886_ (.A(_2886_),
    .X(clknet_0__2886_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2887_ (.A(_2887_),
    .X(clknet_0__2887_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2888_ (.A(_2888_),
    .X(clknet_0__2888_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2889_ (.A(_2889_),
    .X(clknet_0__2889_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2890_ (.A(_2890_),
    .X(clknet_0__2890_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2891_ (.A(_2891_),
    .X(clknet_0__2891_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2892_ (.A(_2892_),
    .X(clknet_0__2892_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2893_ (.A(_2893_),
    .X(clknet_0__2893_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2894_ (.A(_2894_),
    .X(clknet_0__2894_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2895_ (.A(_2895_),
    .X(clknet_0__2895_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2896_ (.A(_2896_),
    .X(clknet_0__2896_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2897_ (.A(_2897_),
    .X(clknet_0__2897_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2898_ (.A(_2898_),
    .X(clknet_0__2898_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2899_ (.A(_2899_),
    .X(clknet_0__2899_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2882_ (.A(clknet_0__2882_),
    .X(clknet_1_0__leaf__2882_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2883_ (.A(clknet_0__2883_),
    .X(clknet_1_0__leaf__2883_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2884_ (.A(clknet_0__2884_),
    .X(clknet_1_0__leaf__2884_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2885_ (.A(clknet_0__2885_),
    .X(clknet_1_0__leaf__2885_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2886_ (.A(clknet_0__2886_),
    .X(clknet_1_0__leaf__2886_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2887_ (.A(clknet_0__2887_),
    .X(clknet_1_0__leaf__2887_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2888_ (.A(clknet_0__2888_),
    .X(clknet_1_0__leaf__2888_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2889_ (.A(clknet_0__2889_),
    .X(clknet_1_0__leaf__2889_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2890_ (.A(clknet_0__2890_),
    .X(clknet_1_0__leaf__2890_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2891_ (.A(clknet_0__2891_),
    .X(clknet_1_0__leaf__2891_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2892_ (.A(clknet_0__2892_),
    .X(clknet_1_0__leaf__2892_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2893_ (.A(clknet_0__2893_),
    .X(clknet_1_0__leaf__2893_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2894_ (.A(clknet_0__2894_),
    .X(clknet_1_0__leaf__2894_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2895_ (.A(clknet_0__2895_),
    .X(clknet_1_0__leaf__2895_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2896_ (.A(clknet_0__2896_),
    .X(clknet_1_0__leaf__2896_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2897_ (.A(clknet_0__2897_),
    .X(clknet_1_0__leaf__2897_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2898_ (.A(clknet_0__2898_),
    .X(clknet_1_0__leaf__2898_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2899_ (.A(clknet_0__2899_),
    .X(clknet_1_0__leaf__2899_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2882_ (.A(clknet_0__2882_),
    .X(clknet_1_1__leaf__2882_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2883_ (.A(clknet_0__2883_),
    .X(clknet_1_1__leaf__2883_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2884_ (.A(clknet_0__2884_),
    .X(clknet_1_1__leaf__2884_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2885_ (.A(clknet_0__2885_),
    .X(clknet_1_1__leaf__2885_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2886_ (.A(clknet_0__2886_),
    .X(clknet_1_1__leaf__2886_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2887_ (.A(clknet_0__2887_),
    .X(clknet_1_1__leaf__2887_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2888_ (.A(clknet_0__2888_),
    .X(clknet_1_1__leaf__2888_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2889_ (.A(clknet_0__2889_),
    .X(clknet_1_1__leaf__2889_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2890_ (.A(clknet_0__2890_),
    .X(clknet_1_1__leaf__2890_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2891_ (.A(clknet_0__2891_),
    .X(clknet_1_1__leaf__2891_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2892_ (.A(clknet_0__2892_),
    .X(clknet_1_1__leaf__2892_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2893_ (.A(clknet_0__2893_),
    .X(clknet_1_1__leaf__2893_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2894_ (.A(clknet_0__2894_),
    .X(clknet_1_1__leaf__2894_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2895_ (.A(clknet_0__2895_),
    .X(clknet_1_1__leaf__2895_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2896_ (.A(clknet_0__2896_),
    .X(clknet_1_1__leaf__2896_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2897_ (.A(clknet_0__2897_),
    .X(clknet_1_1__leaf__2897_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2898_ (.A(clknet_0__2898_),
    .X(clknet_1_1__leaf__2898_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2899_ (.A(clknet_0__2899_),
    .X(clknet_1_1__leaf__2899_));
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(la_data_in_58_43[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(la_data_in_58_43[3]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(la_data_in_58_43[4]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(la_data_in_58_43[5]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(la_data_in_58_43[6]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(la_data_in_58_43[7]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(la_data_in_58_43[8]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(la_data_in_58_43[9]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_4 input17 (.A(la_data_in_60_59[0]),
    .X(net17));
 sky130_fd_sc_hd__buf_2 input18 (.A(la_data_in_60_59[1]),
    .X(net18));
 sky130_fd_sc_hd__buf_2 input19 (.A(la_data_in_65),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(la_data_in_58_43[10]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(la_data_in_58_43[11]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(la_data_in_58_43[12]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(la_data_in_58_43[13]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(la_data_in_58_43[14]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(la_data_in_58_43[15]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(la_data_in_58_43[1]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(la_data_in_58_43[2]),
    .X(net9));
 sky130_fd_sc_hd__buf_12 output20 (.A(net20),
    .X(la_data_out_23_16[0]));
 sky130_fd_sc_hd__buf_12 output21 (.A(net21),
    .X(la_data_out_23_16[1]));
 sky130_fd_sc_hd__buf_12 output22 (.A(net22),
    .X(la_data_out_23_16[2]));
 sky130_fd_sc_hd__buf_12 output23 (.A(net23),
    .X(la_data_out_23_16[3]));
 sky130_fd_sc_hd__buf_12 output24 (.A(net24),
    .X(la_data_out_23_16[4]));
 sky130_fd_sc_hd__buf_12 output25 (.A(net25),
    .X(la_data_out_23_16[5]));
 sky130_fd_sc_hd__buf_12 output26 (.A(net26),
    .X(la_data_out_23_16[6]));
 sky130_fd_sc_hd__buf_12 output27 (.A(net27),
    .X(la_data_out_23_16[7]));
 sky130_fd_sc_hd__buf_12 output28 (.A(net28),
    .X(la_data_out_26_24[0]));
 sky130_fd_sc_hd__buf_12 output29 (.A(net29),
    .X(la_data_out_26_24[1]));
 sky130_fd_sc_hd__buf_12 output30 (.A(net30),
    .X(la_data_out_26_24[2]));
 sky130_fd_sc_hd__buf_12 output31 (.A(net31),
    .X(la_data_out_30_27[0]));
 sky130_fd_sc_hd__buf_12 output32 (.A(net32),
    .X(la_data_out_30_27[1]));
 sky130_fd_sc_hd__buf_12 output33 (.A(net33),
    .X(la_data_out_30_27[2]));
 sky130_fd_sc_hd__buf_12 output34 (.A(net34),
    .X(la_data_out_30_27[3]));
endmodule

