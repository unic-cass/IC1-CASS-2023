magic
tech sky130B
magscale 1 2
timestamp 1676037725
<< nwell >>
rect -38 331 134 704
<< pwell >>
rect 5 49 91 255
rect 0 0 96 49
<< psubdiff >>
rect 31 205 65 229
rect 31 137 65 171
rect 31 79 65 103
<< nsubdiff >>
rect 31 575 65 599
rect 31 492 65 541
rect 31 434 65 458
<< psubdiffcont >>
rect 31 171 65 205
rect 31 103 65 137
<< nsubdiffcont >>
rect 31 541 65 575
rect 31 458 65 492
<< locali >>
rect 0 649 31 683
rect 65 649 96 683
rect 18 575 78 613
rect 18 541 31 575
rect 65 541 78 575
rect 18 492 78 541
rect 18 458 31 492
rect 65 458 78 492
rect 18 378 78 458
rect 18 205 78 288
rect 18 171 31 205
rect 65 171 78 205
rect 18 137 78 171
rect 18 103 31 137
rect 65 103 78 137
rect 18 53 78 103
rect 0 -17 31 17
rect 65 -17 96 17
<< viali >>
rect 31 649 65 683
rect 31 -17 65 17
<< metal1 >>
rect 0 683 96 715
rect 0 649 31 683
rect 65 649 96 683
rect 0 617 96 649
rect 0 17 96 49
rect 0 -17 31 17
rect 65 -17 96 17
rect 0 -49 96 -17
<< labels >>
flabel pwell s 0 0 96 49 0 FreeSans 200 0 0 0 VNB
port 1 nsew
flabel nwell s 0 617 96 666 0 FreeSans 200 0 0 0 VPB
port 2 nsew
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 VNB
port 1 nsew
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 VNB
port 1 nsew
flabel locali s 31 94 65 128 0 FreeSans 340 0 0 0 VNB
port 1 nsew
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 VPB
port 2 nsew
flabel locali s 31 464 65 498 0 FreeSans 340 0 0 0 VPB
port 2 nsew
flabel locali s 31 538 65 572 0 FreeSans 340 0 0 0 VPB
port 2 nsew
rlabel comment s 0 0 0 0 4 SKY130_FD_IO__TAP_1
flabel metal1 s 0 617 96 666 0 FreeSans 200 0 0 0 VPWR
port 3 nsew
flabel metal1 s 0 0 96 49 0 FreeSans 200 0 0 0 VGND
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 96 666
string GDS_END 269468
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 266434
<< end >>
