magic
tech sky130B
magscale 1 2
timestamp 1676037725
<< locali >>
rect 266 1369 616 1388
rect 266 1263 280 1369
rect 602 1263 616 1369
rect 266 1249 616 1263
rect 266 125 616 139
rect 266 19 280 125
rect 602 19 616 125
rect 266 0 616 19
<< viali >>
rect 280 1263 602 1369
rect 280 19 602 125
<< obsli1 >>
rect 120 1225 186 1291
rect 696 1225 762 1291
rect 120 1203 160 1225
rect 722 1203 762 1225
rect 41 1179 160 1203
rect 41 1145 60 1179
rect 94 1145 160 1179
rect 41 1107 160 1145
rect 41 1073 60 1107
rect 94 1073 160 1107
rect 41 1035 160 1073
rect 41 1001 60 1035
rect 94 1001 160 1035
rect 41 963 160 1001
rect 41 929 60 963
rect 94 929 160 963
rect 41 891 160 929
rect 41 857 60 891
rect 94 857 160 891
rect 41 819 160 857
rect 41 785 60 819
rect 94 785 160 819
rect 41 747 160 785
rect 41 713 60 747
rect 94 713 160 747
rect 41 675 160 713
rect 41 641 60 675
rect 94 641 160 675
rect 41 603 160 641
rect 41 569 60 603
rect 94 569 160 603
rect 41 531 160 569
rect 41 497 60 531
rect 94 497 160 531
rect 41 459 160 497
rect 41 425 60 459
rect 94 425 160 459
rect 41 387 160 425
rect 41 353 60 387
rect 94 353 160 387
rect 41 315 160 353
rect 41 281 60 315
rect 94 281 160 315
rect 41 243 160 281
rect 41 209 60 243
rect 94 209 160 243
rect 41 185 160 209
rect 212 185 246 1203
rect 318 185 352 1203
rect 424 185 458 1203
rect 530 185 564 1203
rect 636 185 670 1203
rect 722 1179 841 1203
rect 722 1145 788 1179
rect 822 1145 841 1179
rect 722 1107 841 1145
rect 722 1073 788 1107
rect 822 1073 841 1107
rect 722 1035 841 1073
rect 722 1001 788 1035
rect 822 1001 841 1035
rect 722 963 841 1001
rect 722 929 788 963
rect 822 929 841 963
rect 722 891 841 929
rect 722 857 788 891
rect 822 857 841 891
rect 722 819 841 857
rect 722 785 788 819
rect 822 785 841 819
rect 722 747 841 785
rect 722 713 788 747
rect 822 713 841 747
rect 722 675 841 713
rect 722 641 788 675
rect 822 641 841 675
rect 722 603 841 641
rect 722 569 788 603
rect 822 569 841 603
rect 722 531 841 569
rect 722 497 788 531
rect 822 497 841 531
rect 722 459 841 497
rect 722 425 788 459
rect 822 425 841 459
rect 722 387 841 425
rect 722 353 788 387
rect 822 353 841 387
rect 722 315 841 353
rect 722 281 788 315
rect 822 281 841 315
rect 722 243 841 281
rect 722 209 788 243
rect 822 209 841 243
rect 722 185 841 209
rect 120 163 160 185
rect 722 163 762 185
rect 120 97 186 163
rect 696 97 762 163
<< obsli1c >>
rect 60 1145 94 1179
rect 60 1073 94 1107
rect 60 1001 94 1035
rect 60 929 94 963
rect 60 857 94 891
rect 60 785 94 819
rect 60 713 94 747
rect 60 641 94 675
rect 60 569 94 603
rect 60 497 94 531
rect 60 425 94 459
rect 60 353 94 387
rect 60 281 94 315
rect 60 209 94 243
rect 788 1145 822 1179
rect 788 1073 822 1107
rect 788 1001 822 1035
rect 788 929 822 963
rect 788 857 822 891
rect 788 785 822 819
rect 788 713 822 747
rect 788 641 822 675
rect 788 569 822 603
rect 788 497 822 531
rect 788 425 822 459
rect 788 353 822 387
rect 788 281 822 315
rect 788 209 822 243
<< metal1 >>
rect 264 1369 618 1388
rect 264 1263 280 1369
rect 602 1263 618 1369
rect 264 1251 618 1263
rect 41 1179 100 1191
rect 41 1145 60 1179
rect 94 1145 100 1179
rect 41 1107 100 1145
rect 41 1073 60 1107
rect 94 1073 100 1107
rect 41 1035 100 1073
rect 41 1001 60 1035
rect 94 1001 100 1035
rect 41 963 100 1001
rect 41 929 60 963
rect 94 929 100 963
rect 41 891 100 929
rect 41 857 60 891
rect 94 857 100 891
rect 41 819 100 857
rect 41 785 60 819
rect 94 785 100 819
rect 41 747 100 785
rect 41 713 60 747
rect 94 713 100 747
rect 41 675 100 713
rect 41 641 60 675
rect 94 641 100 675
rect 41 603 100 641
rect 41 569 60 603
rect 94 569 100 603
rect 41 531 100 569
rect 41 497 60 531
rect 94 497 100 531
rect 41 459 100 497
rect 41 425 60 459
rect 94 425 100 459
rect 41 387 100 425
rect 41 353 60 387
rect 94 353 100 387
rect 41 315 100 353
rect 41 281 60 315
rect 94 281 100 315
rect 41 243 100 281
rect 41 209 60 243
rect 94 209 100 243
rect 41 197 100 209
rect 782 1179 841 1191
rect 782 1145 788 1179
rect 822 1145 841 1179
rect 782 1107 841 1145
rect 782 1073 788 1107
rect 822 1073 841 1107
rect 782 1035 841 1073
rect 782 1001 788 1035
rect 822 1001 841 1035
rect 782 963 841 1001
rect 782 929 788 963
rect 822 929 841 963
rect 782 891 841 929
rect 782 857 788 891
rect 822 857 841 891
rect 782 819 841 857
rect 782 785 788 819
rect 822 785 841 819
rect 782 747 841 785
rect 782 713 788 747
rect 822 713 841 747
rect 782 675 841 713
rect 782 641 788 675
rect 822 641 841 675
rect 782 603 841 641
rect 782 569 788 603
rect 822 569 841 603
rect 782 531 841 569
rect 782 497 788 531
rect 822 497 841 531
rect 782 459 841 497
rect 782 425 788 459
rect 822 425 841 459
rect 782 387 841 425
rect 782 353 788 387
rect 822 353 841 387
rect 782 315 841 353
rect 782 281 788 315
rect 822 281 841 315
rect 782 243 841 281
rect 782 209 788 243
rect 822 209 841 243
rect 782 197 841 209
rect 264 125 618 137
rect 264 19 280 125
rect 602 19 618 125
rect 264 0 618 19
<< obsm1 >>
rect 203 197 255 1191
rect 309 197 361 1191
rect 415 197 467 1191
rect 521 197 573 1191
rect 627 197 679 1191
<< metal2 >>
rect 14 719 868 1191
rect 14 197 868 669
<< labels >>
rlabel metal2 s 14 719 868 1191 6 DRAIN
port 1 nsew
rlabel viali s 280 1263 602 1369 6 GATE
port 2 nsew
rlabel viali s 280 19 602 125 6 GATE
port 2 nsew
rlabel locali s 266 1249 616 1388 6 GATE
port 2 nsew
rlabel locali s 266 0 616 139 6 GATE
port 2 nsew
rlabel metal1 s 264 1251 618 1388 6 GATE
port 2 nsew
rlabel metal1 s 264 0 618 137 6 GATE
port 2 nsew
rlabel metal2 s 14 197 868 669 6 SOURCE
port 3 nsew
rlabel metal1 s 41 197 100 1191 6 SUBSTRATE
port 4 nsew
rlabel metal1 s 782 197 841 1191 6 SUBSTRATE
port 4 nsew
<< properties >>
string FIXED_BBOX 14 0 868 1388
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 3193000
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 3164878
string device primitive
<< end >>
