magic
tech sky130A
magscale 1 2
timestamp 1676037725
<< nwell >>
rect 0 1331 3633 2349
rect 2202 1178 3633 1331
<< pwell >>
rect 181 1100 970 1240
rect 181 988 3592 1100
rect 235 846 3592 988
rect 235 101 3633 846
rect 123 10 3633 101
<< mvnmos >>
rect 260 1014 380 1214
rect 483 914 583 1214
rect 637 914 737 1214
rect 791 914 891 1214
rect 1057 990 1857 1074
rect 1913 990 3513 1074
rect 314 220 414 820
rect 470 220 570 820
rect 626 220 726 820
rect 782 220 882 820
rect 1048 220 1148 820
rect 1204 220 1304 820
rect 1360 220 1460 820
rect 1516 220 1616 820
rect 1672 220 1772 820
rect 1828 220 1928 820
rect 1984 220 2084 820
rect 2140 220 2240 820
rect 2296 220 2396 820
rect 2452 220 2552 820
rect 2608 220 2708 820
rect 2874 220 2974 820
rect 3030 220 3130 820
rect 3186 220 3286 820
rect 3342 220 3442 820
<< mvpmos >>
rect 150 1898 250 2098
rect 306 1898 406 2098
rect 462 1898 562 2098
rect 618 1898 718 2098
rect 821 2014 2421 2098
rect 150 1397 250 1597
rect 306 1397 406 1597
rect 483 1397 643 1597
rect 699 1397 859 1597
rect 915 1397 1075 1597
rect 1131 1397 1291 1597
rect 1347 1397 1507 1597
rect 1563 1397 1723 1597
rect 1779 1397 1939 1597
rect 1995 1397 2155 1597
rect 2321 1244 2421 1844
rect 2587 1244 2687 1844
rect 2743 1244 2843 1844
rect 2899 1244 2999 1844
rect 3055 1244 3155 1844
rect 3258 1244 3358 2244
rect 3414 1244 3514 2244
<< mvndiff >>
rect 207 1196 260 1214
rect 207 1162 215 1196
rect 249 1162 260 1196
rect 207 1128 260 1162
rect 207 1094 215 1128
rect 249 1094 260 1128
rect 207 1060 260 1094
rect 207 1026 215 1060
rect 249 1026 260 1060
rect 207 1014 260 1026
rect 380 1164 483 1214
rect 380 1130 438 1164
rect 472 1130 483 1164
rect 380 1096 483 1130
rect 380 1062 438 1096
rect 472 1062 483 1096
rect 380 1028 483 1062
rect 380 1014 438 1028
rect 430 994 438 1014
rect 472 994 483 1028
rect 430 960 483 994
rect 430 926 438 960
rect 472 926 483 960
rect 430 914 483 926
rect 583 914 637 1214
rect 737 914 791 1214
rect 891 1164 944 1214
rect 891 1130 902 1164
rect 936 1130 944 1164
rect 891 1096 944 1130
rect 891 1062 902 1096
rect 936 1062 944 1096
rect 891 1028 944 1062
rect 891 994 902 1028
rect 936 994 944 1028
rect 891 960 944 994
rect 1004 1062 1057 1074
rect 1004 1028 1012 1062
rect 1046 1028 1057 1062
rect 1004 990 1057 1028
rect 1857 1062 1913 1074
rect 1857 1028 1868 1062
rect 1902 1028 1913 1062
rect 1857 990 1913 1028
rect 3513 1062 3566 1074
rect 3513 1028 3524 1062
rect 3558 1028 3566 1062
rect 3513 990 3566 1028
rect 891 926 902 960
rect 936 926 944 960
rect 891 914 944 926
rect 261 742 314 820
rect 261 708 269 742
rect 303 708 314 742
rect 261 674 314 708
rect 261 640 269 674
rect 303 640 314 674
rect 261 606 314 640
rect 261 572 269 606
rect 303 572 314 606
rect 261 538 314 572
rect 261 504 269 538
rect 303 504 314 538
rect 261 470 314 504
rect 261 436 269 470
rect 303 436 314 470
rect 261 402 314 436
rect 261 368 269 402
rect 303 368 314 402
rect 261 334 314 368
rect 261 300 269 334
rect 303 300 314 334
rect 261 266 314 300
rect 261 232 269 266
rect 303 232 314 266
rect 261 220 314 232
rect 414 742 470 820
rect 414 708 425 742
rect 459 708 470 742
rect 414 674 470 708
rect 414 640 425 674
rect 459 640 470 674
rect 414 606 470 640
rect 414 572 425 606
rect 459 572 470 606
rect 414 538 470 572
rect 414 504 425 538
rect 459 504 470 538
rect 414 470 470 504
rect 414 436 425 470
rect 459 436 470 470
rect 414 402 470 436
rect 414 368 425 402
rect 459 368 470 402
rect 414 334 470 368
rect 414 300 425 334
rect 459 300 470 334
rect 414 266 470 300
rect 414 232 425 266
rect 459 232 470 266
rect 414 220 470 232
rect 570 742 626 820
rect 570 708 581 742
rect 615 708 626 742
rect 570 674 626 708
rect 570 640 581 674
rect 615 640 626 674
rect 570 606 626 640
rect 570 572 581 606
rect 615 572 626 606
rect 570 538 626 572
rect 570 504 581 538
rect 615 504 626 538
rect 570 470 626 504
rect 570 436 581 470
rect 615 436 626 470
rect 570 402 626 436
rect 570 368 581 402
rect 615 368 626 402
rect 570 334 626 368
rect 570 300 581 334
rect 615 300 626 334
rect 570 266 626 300
rect 570 232 581 266
rect 615 232 626 266
rect 570 220 626 232
rect 726 742 782 820
rect 726 708 737 742
rect 771 708 782 742
rect 726 674 782 708
rect 726 640 737 674
rect 771 640 782 674
rect 726 606 782 640
rect 726 572 737 606
rect 771 572 782 606
rect 726 538 782 572
rect 726 504 737 538
rect 771 504 782 538
rect 726 470 782 504
rect 726 436 737 470
rect 771 436 782 470
rect 726 402 782 436
rect 726 368 737 402
rect 771 368 782 402
rect 726 334 782 368
rect 726 300 737 334
rect 771 300 782 334
rect 726 266 782 300
rect 726 232 737 266
rect 771 232 782 266
rect 726 220 782 232
rect 882 742 935 820
rect 882 708 893 742
rect 927 708 935 742
rect 882 674 935 708
rect 882 640 893 674
rect 927 640 935 674
rect 882 606 935 640
rect 882 572 893 606
rect 927 572 935 606
rect 882 538 935 572
rect 882 504 893 538
rect 927 504 935 538
rect 882 470 935 504
rect 882 436 893 470
rect 927 436 935 470
rect 882 402 935 436
rect 882 368 893 402
rect 927 368 935 402
rect 882 334 935 368
rect 882 300 893 334
rect 927 300 935 334
rect 882 266 935 300
rect 882 232 893 266
rect 927 232 935 266
rect 882 220 935 232
rect 995 742 1048 820
rect 995 708 1003 742
rect 1037 708 1048 742
rect 995 674 1048 708
rect 995 640 1003 674
rect 1037 640 1048 674
rect 995 606 1048 640
rect 995 572 1003 606
rect 1037 572 1048 606
rect 995 538 1048 572
rect 995 504 1003 538
rect 1037 504 1048 538
rect 995 470 1048 504
rect 995 436 1003 470
rect 1037 436 1048 470
rect 995 402 1048 436
rect 995 368 1003 402
rect 1037 368 1048 402
rect 995 334 1048 368
rect 995 300 1003 334
rect 1037 300 1048 334
rect 995 266 1048 300
rect 995 232 1003 266
rect 1037 232 1048 266
rect 995 220 1048 232
rect 1148 742 1204 820
rect 1148 708 1159 742
rect 1193 708 1204 742
rect 1148 674 1204 708
rect 1148 640 1159 674
rect 1193 640 1204 674
rect 1148 606 1204 640
rect 1148 572 1159 606
rect 1193 572 1204 606
rect 1148 538 1204 572
rect 1148 504 1159 538
rect 1193 504 1204 538
rect 1148 470 1204 504
rect 1148 436 1159 470
rect 1193 436 1204 470
rect 1148 402 1204 436
rect 1148 368 1159 402
rect 1193 368 1204 402
rect 1148 334 1204 368
rect 1148 300 1159 334
rect 1193 300 1204 334
rect 1148 266 1204 300
rect 1148 232 1159 266
rect 1193 232 1204 266
rect 1148 220 1204 232
rect 1304 742 1360 820
rect 1304 708 1315 742
rect 1349 708 1360 742
rect 1304 674 1360 708
rect 1304 640 1315 674
rect 1349 640 1360 674
rect 1304 606 1360 640
rect 1304 572 1315 606
rect 1349 572 1360 606
rect 1304 538 1360 572
rect 1304 504 1315 538
rect 1349 504 1360 538
rect 1304 470 1360 504
rect 1304 436 1315 470
rect 1349 436 1360 470
rect 1304 402 1360 436
rect 1304 368 1315 402
rect 1349 368 1360 402
rect 1304 334 1360 368
rect 1304 300 1315 334
rect 1349 300 1360 334
rect 1304 266 1360 300
rect 1304 232 1315 266
rect 1349 232 1360 266
rect 1304 220 1360 232
rect 1460 742 1516 820
rect 1460 708 1471 742
rect 1505 708 1516 742
rect 1460 674 1516 708
rect 1460 640 1471 674
rect 1505 640 1516 674
rect 1460 606 1516 640
rect 1460 572 1471 606
rect 1505 572 1516 606
rect 1460 538 1516 572
rect 1460 504 1471 538
rect 1505 504 1516 538
rect 1460 470 1516 504
rect 1460 436 1471 470
rect 1505 436 1516 470
rect 1460 402 1516 436
rect 1460 368 1471 402
rect 1505 368 1516 402
rect 1460 334 1516 368
rect 1460 300 1471 334
rect 1505 300 1516 334
rect 1460 266 1516 300
rect 1460 232 1471 266
rect 1505 232 1516 266
rect 1460 220 1516 232
rect 1616 742 1672 820
rect 1616 708 1627 742
rect 1661 708 1672 742
rect 1616 674 1672 708
rect 1616 640 1627 674
rect 1661 640 1672 674
rect 1616 606 1672 640
rect 1616 572 1627 606
rect 1661 572 1672 606
rect 1616 538 1672 572
rect 1616 504 1627 538
rect 1661 504 1672 538
rect 1616 470 1672 504
rect 1616 436 1627 470
rect 1661 436 1672 470
rect 1616 402 1672 436
rect 1616 368 1627 402
rect 1661 368 1672 402
rect 1616 334 1672 368
rect 1616 300 1627 334
rect 1661 300 1672 334
rect 1616 266 1672 300
rect 1616 232 1627 266
rect 1661 232 1672 266
rect 1616 220 1672 232
rect 1772 742 1828 820
rect 1772 708 1783 742
rect 1817 708 1828 742
rect 1772 674 1828 708
rect 1772 640 1783 674
rect 1817 640 1828 674
rect 1772 606 1828 640
rect 1772 572 1783 606
rect 1817 572 1828 606
rect 1772 538 1828 572
rect 1772 504 1783 538
rect 1817 504 1828 538
rect 1772 470 1828 504
rect 1772 436 1783 470
rect 1817 436 1828 470
rect 1772 402 1828 436
rect 1772 368 1783 402
rect 1817 368 1828 402
rect 1772 334 1828 368
rect 1772 300 1783 334
rect 1817 300 1828 334
rect 1772 266 1828 300
rect 1772 232 1783 266
rect 1817 232 1828 266
rect 1772 220 1828 232
rect 1928 742 1984 820
rect 1928 708 1939 742
rect 1973 708 1984 742
rect 1928 674 1984 708
rect 1928 640 1939 674
rect 1973 640 1984 674
rect 1928 606 1984 640
rect 1928 572 1939 606
rect 1973 572 1984 606
rect 1928 538 1984 572
rect 1928 504 1939 538
rect 1973 504 1984 538
rect 1928 470 1984 504
rect 1928 436 1939 470
rect 1973 436 1984 470
rect 1928 402 1984 436
rect 1928 368 1939 402
rect 1973 368 1984 402
rect 1928 334 1984 368
rect 1928 300 1939 334
rect 1973 300 1984 334
rect 1928 266 1984 300
rect 1928 232 1939 266
rect 1973 232 1984 266
rect 1928 220 1984 232
rect 2084 742 2140 820
rect 2084 708 2095 742
rect 2129 708 2140 742
rect 2084 674 2140 708
rect 2084 640 2095 674
rect 2129 640 2140 674
rect 2084 606 2140 640
rect 2084 572 2095 606
rect 2129 572 2140 606
rect 2084 538 2140 572
rect 2084 504 2095 538
rect 2129 504 2140 538
rect 2084 470 2140 504
rect 2084 436 2095 470
rect 2129 436 2140 470
rect 2084 402 2140 436
rect 2084 368 2095 402
rect 2129 368 2140 402
rect 2084 334 2140 368
rect 2084 300 2095 334
rect 2129 300 2140 334
rect 2084 266 2140 300
rect 2084 232 2095 266
rect 2129 232 2140 266
rect 2084 220 2140 232
rect 2240 742 2296 820
rect 2240 708 2251 742
rect 2285 708 2296 742
rect 2240 674 2296 708
rect 2240 640 2251 674
rect 2285 640 2296 674
rect 2240 606 2296 640
rect 2240 572 2251 606
rect 2285 572 2296 606
rect 2240 538 2296 572
rect 2240 504 2251 538
rect 2285 504 2296 538
rect 2240 470 2296 504
rect 2240 436 2251 470
rect 2285 436 2296 470
rect 2240 402 2296 436
rect 2240 368 2251 402
rect 2285 368 2296 402
rect 2240 334 2296 368
rect 2240 300 2251 334
rect 2285 300 2296 334
rect 2240 266 2296 300
rect 2240 232 2251 266
rect 2285 232 2296 266
rect 2240 220 2296 232
rect 2396 742 2452 820
rect 2396 708 2407 742
rect 2441 708 2452 742
rect 2396 674 2452 708
rect 2396 640 2407 674
rect 2441 640 2452 674
rect 2396 606 2452 640
rect 2396 572 2407 606
rect 2441 572 2452 606
rect 2396 538 2452 572
rect 2396 504 2407 538
rect 2441 504 2452 538
rect 2396 470 2452 504
rect 2396 436 2407 470
rect 2441 436 2452 470
rect 2396 402 2452 436
rect 2396 368 2407 402
rect 2441 368 2452 402
rect 2396 334 2452 368
rect 2396 300 2407 334
rect 2441 300 2452 334
rect 2396 266 2452 300
rect 2396 232 2407 266
rect 2441 232 2452 266
rect 2396 220 2452 232
rect 2552 742 2608 820
rect 2552 708 2563 742
rect 2597 708 2608 742
rect 2552 674 2608 708
rect 2552 640 2563 674
rect 2597 640 2608 674
rect 2552 606 2608 640
rect 2552 572 2563 606
rect 2597 572 2608 606
rect 2552 538 2608 572
rect 2552 504 2563 538
rect 2597 504 2608 538
rect 2552 470 2608 504
rect 2552 436 2563 470
rect 2597 436 2608 470
rect 2552 402 2608 436
rect 2552 368 2563 402
rect 2597 368 2608 402
rect 2552 334 2608 368
rect 2552 300 2563 334
rect 2597 300 2608 334
rect 2552 266 2608 300
rect 2552 232 2563 266
rect 2597 232 2608 266
rect 2552 220 2608 232
rect 2708 742 2761 820
rect 2708 708 2719 742
rect 2753 708 2761 742
rect 2708 674 2761 708
rect 2708 640 2719 674
rect 2753 640 2761 674
rect 2708 606 2761 640
rect 2708 572 2719 606
rect 2753 572 2761 606
rect 2708 538 2761 572
rect 2708 504 2719 538
rect 2753 504 2761 538
rect 2708 470 2761 504
rect 2708 436 2719 470
rect 2753 436 2761 470
rect 2708 402 2761 436
rect 2708 368 2719 402
rect 2753 368 2761 402
rect 2708 334 2761 368
rect 2708 300 2719 334
rect 2753 300 2761 334
rect 2708 266 2761 300
rect 2708 232 2719 266
rect 2753 232 2761 266
rect 2708 220 2761 232
rect 2821 742 2874 820
rect 2821 708 2829 742
rect 2863 708 2874 742
rect 2821 674 2874 708
rect 2821 640 2829 674
rect 2863 640 2874 674
rect 2821 606 2874 640
rect 2821 572 2829 606
rect 2863 572 2874 606
rect 2821 538 2874 572
rect 2821 504 2829 538
rect 2863 504 2874 538
rect 2821 470 2874 504
rect 2821 436 2829 470
rect 2863 436 2874 470
rect 2821 402 2874 436
rect 2821 368 2829 402
rect 2863 368 2874 402
rect 2821 334 2874 368
rect 2821 300 2829 334
rect 2863 300 2874 334
rect 2821 266 2874 300
rect 2821 232 2829 266
rect 2863 232 2874 266
rect 2821 220 2874 232
rect 2974 742 3030 820
rect 2974 708 2985 742
rect 3019 708 3030 742
rect 2974 674 3030 708
rect 2974 640 2985 674
rect 3019 640 3030 674
rect 2974 606 3030 640
rect 2974 572 2985 606
rect 3019 572 3030 606
rect 2974 538 3030 572
rect 2974 504 2985 538
rect 3019 504 3030 538
rect 2974 470 3030 504
rect 2974 436 2985 470
rect 3019 436 3030 470
rect 2974 402 3030 436
rect 2974 368 2985 402
rect 3019 368 3030 402
rect 2974 334 3030 368
rect 2974 300 2985 334
rect 3019 300 3030 334
rect 2974 266 3030 300
rect 2974 232 2985 266
rect 3019 232 3030 266
rect 2974 220 3030 232
rect 3130 742 3186 820
rect 3130 708 3141 742
rect 3175 708 3186 742
rect 3130 674 3186 708
rect 3130 640 3141 674
rect 3175 640 3186 674
rect 3130 606 3186 640
rect 3130 572 3141 606
rect 3175 572 3186 606
rect 3130 538 3186 572
rect 3130 504 3141 538
rect 3175 504 3186 538
rect 3130 470 3186 504
rect 3130 436 3141 470
rect 3175 436 3186 470
rect 3130 402 3186 436
rect 3130 368 3141 402
rect 3175 368 3186 402
rect 3130 334 3186 368
rect 3130 300 3141 334
rect 3175 300 3186 334
rect 3130 266 3186 300
rect 3130 232 3141 266
rect 3175 232 3186 266
rect 3130 220 3186 232
rect 3286 742 3342 820
rect 3286 708 3297 742
rect 3331 708 3342 742
rect 3286 674 3342 708
rect 3286 640 3297 674
rect 3331 640 3342 674
rect 3286 606 3342 640
rect 3286 572 3297 606
rect 3331 572 3342 606
rect 3286 538 3342 572
rect 3286 504 3297 538
rect 3331 504 3342 538
rect 3286 470 3342 504
rect 3286 436 3297 470
rect 3331 436 3342 470
rect 3286 402 3342 436
rect 3286 368 3297 402
rect 3331 368 3342 402
rect 3286 334 3342 368
rect 3286 300 3297 334
rect 3331 300 3342 334
rect 3286 266 3342 300
rect 3286 232 3297 266
rect 3331 232 3342 266
rect 3286 220 3342 232
rect 3442 742 3495 820
rect 3442 708 3453 742
rect 3487 708 3495 742
rect 3442 674 3495 708
rect 3442 640 3453 674
rect 3487 640 3495 674
rect 3442 606 3495 640
rect 3442 572 3453 606
rect 3487 572 3495 606
rect 3442 538 3495 572
rect 3442 504 3453 538
rect 3487 504 3495 538
rect 3442 470 3495 504
rect 3442 436 3453 470
rect 3487 436 3495 470
rect 3442 402 3495 436
rect 3442 368 3453 402
rect 3487 368 3495 402
rect 3442 334 3495 368
rect 3442 300 3453 334
rect 3487 300 3495 334
rect 3442 266 3495 300
rect 3442 232 3453 266
rect 3487 232 3495 266
rect 3442 220 3495 232
<< mvpdiff >>
rect 97 2080 150 2098
rect 97 2046 105 2080
rect 139 2046 150 2080
rect 97 2012 150 2046
rect 97 1978 105 2012
rect 139 1978 150 2012
rect 97 1944 150 1978
rect 97 1910 105 1944
rect 139 1910 150 1944
rect 97 1898 150 1910
rect 250 2080 306 2098
rect 250 2046 261 2080
rect 295 2046 306 2080
rect 250 2012 306 2046
rect 250 1978 261 2012
rect 295 1978 306 2012
rect 250 1944 306 1978
rect 250 1910 261 1944
rect 295 1910 306 1944
rect 250 1898 306 1910
rect 406 2080 462 2098
rect 406 2046 417 2080
rect 451 2046 462 2080
rect 406 2012 462 2046
rect 406 1978 417 2012
rect 451 1978 462 2012
rect 406 1944 462 1978
rect 406 1910 417 1944
rect 451 1910 462 1944
rect 406 1898 462 1910
rect 562 2080 618 2098
rect 562 2046 573 2080
rect 607 2046 618 2080
rect 562 2012 618 2046
rect 562 1978 573 2012
rect 607 1978 618 2012
rect 562 1944 618 1978
rect 562 1910 573 1944
rect 607 1910 618 1944
rect 562 1898 618 1910
rect 718 2080 821 2098
rect 718 2046 729 2080
rect 763 2046 821 2080
rect 718 2014 821 2046
rect 2421 2060 2474 2098
rect 2421 2026 2432 2060
rect 2466 2026 2474 2060
rect 2421 2014 2474 2026
rect 718 2012 771 2014
rect 718 1978 729 2012
rect 763 1978 771 2012
rect 718 1944 771 1978
rect 718 1910 729 1944
rect 763 1910 771 1944
rect 3205 2174 3258 2244
rect 3205 2140 3213 2174
rect 3247 2140 3258 2174
rect 3205 2106 3258 2140
rect 3205 2072 3213 2106
rect 3247 2072 3258 2106
rect 3205 2038 3258 2072
rect 3205 2004 3213 2038
rect 3247 2004 3258 2038
rect 3205 1970 3258 2004
rect 718 1898 771 1910
rect 3205 1936 3213 1970
rect 3247 1936 3258 1970
rect 3205 1902 3258 1936
rect 3205 1868 3213 1902
rect 3247 1868 3258 1902
rect 3205 1844 3258 1868
rect 2268 1766 2321 1844
rect 2268 1732 2276 1766
rect 2310 1732 2321 1766
rect 2268 1698 2321 1732
rect 2268 1664 2276 1698
rect 2310 1664 2321 1698
rect 2268 1630 2321 1664
rect 97 1579 150 1597
rect 97 1545 105 1579
rect 139 1545 150 1579
rect 97 1511 150 1545
rect 97 1477 105 1511
rect 139 1477 150 1511
rect 97 1443 150 1477
rect 97 1409 105 1443
rect 139 1409 150 1443
rect 97 1397 150 1409
rect 250 1579 306 1597
rect 250 1545 261 1579
rect 295 1545 306 1579
rect 250 1511 306 1545
rect 250 1477 261 1511
rect 295 1477 306 1511
rect 250 1443 306 1477
rect 250 1409 261 1443
rect 295 1409 306 1443
rect 250 1397 306 1409
rect 406 1579 483 1597
rect 406 1545 438 1579
rect 472 1545 483 1579
rect 406 1511 483 1545
rect 406 1477 438 1511
rect 472 1477 483 1511
rect 406 1443 483 1477
rect 406 1409 438 1443
rect 472 1409 483 1443
rect 406 1397 483 1409
rect 643 1579 699 1597
rect 643 1545 654 1579
rect 688 1545 699 1579
rect 643 1511 699 1545
rect 643 1477 654 1511
rect 688 1477 699 1511
rect 643 1443 699 1477
rect 643 1409 654 1443
rect 688 1409 699 1443
rect 643 1397 699 1409
rect 859 1579 915 1597
rect 859 1545 870 1579
rect 904 1545 915 1579
rect 859 1511 915 1545
rect 859 1477 870 1511
rect 904 1477 915 1511
rect 859 1443 915 1477
rect 859 1409 870 1443
rect 904 1409 915 1443
rect 859 1397 915 1409
rect 1075 1579 1131 1597
rect 1075 1545 1086 1579
rect 1120 1545 1131 1579
rect 1075 1511 1131 1545
rect 1075 1477 1086 1511
rect 1120 1477 1131 1511
rect 1075 1443 1131 1477
rect 1075 1409 1086 1443
rect 1120 1409 1131 1443
rect 1075 1397 1131 1409
rect 1291 1579 1347 1597
rect 1291 1545 1302 1579
rect 1336 1545 1347 1579
rect 1291 1511 1347 1545
rect 1291 1477 1302 1511
rect 1336 1477 1347 1511
rect 1291 1443 1347 1477
rect 1291 1409 1302 1443
rect 1336 1409 1347 1443
rect 1291 1397 1347 1409
rect 1507 1579 1563 1597
rect 1507 1545 1518 1579
rect 1552 1545 1563 1579
rect 1507 1511 1563 1545
rect 1507 1477 1518 1511
rect 1552 1477 1563 1511
rect 1507 1443 1563 1477
rect 1507 1409 1518 1443
rect 1552 1409 1563 1443
rect 1507 1397 1563 1409
rect 1723 1579 1779 1597
rect 1723 1545 1734 1579
rect 1768 1545 1779 1579
rect 1723 1511 1779 1545
rect 1723 1477 1734 1511
rect 1768 1477 1779 1511
rect 1723 1443 1779 1477
rect 1723 1409 1734 1443
rect 1768 1409 1779 1443
rect 1723 1397 1779 1409
rect 1939 1579 1995 1597
rect 1939 1545 1950 1579
rect 1984 1545 1995 1579
rect 1939 1511 1995 1545
rect 1939 1477 1950 1511
rect 1984 1477 1995 1511
rect 1939 1443 1995 1477
rect 1939 1409 1950 1443
rect 1984 1409 1995 1443
rect 1939 1397 1995 1409
rect 2155 1579 2208 1597
rect 2155 1545 2166 1579
rect 2200 1545 2208 1579
rect 2155 1511 2208 1545
rect 2155 1477 2166 1511
rect 2200 1477 2208 1511
rect 2155 1443 2208 1477
rect 2155 1409 2166 1443
rect 2200 1409 2208 1443
rect 2155 1397 2208 1409
rect 2268 1596 2276 1630
rect 2310 1596 2321 1630
rect 2268 1562 2321 1596
rect 2268 1528 2276 1562
rect 2310 1528 2321 1562
rect 2268 1494 2321 1528
rect 2268 1460 2276 1494
rect 2310 1460 2321 1494
rect 2268 1426 2321 1460
rect 2268 1392 2276 1426
rect 2310 1392 2321 1426
rect 2268 1358 2321 1392
rect 2268 1324 2276 1358
rect 2310 1324 2321 1358
rect 2268 1290 2321 1324
rect 2268 1256 2276 1290
rect 2310 1256 2321 1290
rect 2268 1244 2321 1256
rect 2421 1766 2474 1844
rect 2421 1732 2432 1766
rect 2466 1732 2474 1766
rect 2421 1698 2474 1732
rect 2421 1664 2432 1698
rect 2466 1664 2474 1698
rect 2421 1630 2474 1664
rect 2421 1596 2432 1630
rect 2466 1596 2474 1630
rect 2421 1562 2474 1596
rect 2421 1528 2432 1562
rect 2466 1528 2474 1562
rect 2421 1494 2474 1528
rect 2421 1460 2432 1494
rect 2466 1460 2474 1494
rect 2421 1426 2474 1460
rect 2421 1392 2432 1426
rect 2466 1392 2474 1426
rect 2421 1358 2474 1392
rect 2421 1324 2432 1358
rect 2466 1324 2474 1358
rect 2421 1290 2474 1324
rect 2421 1256 2432 1290
rect 2466 1256 2474 1290
rect 2421 1244 2474 1256
rect 2534 1766 2587 1844
rect 2534 1732 2542 1766
rect 2576 1732 2587 1766
rect 2534 1698 2587 1732
rect 2534 1664 2542 1698
rect 2576 1664 2587 1698
rect 2534 1630 2587 1664
rect 2534 1596 2542 1630
rect 2576 1596 2587 1630
rect 2534 1562 2587 1596
rect 2534 1528 2542 1562
rect 2576 1528 2587 1562
rect 2534 1494 2587 1528
rect 2534 1460 2542 1494
rect 2576 1460 2587 1494
rect 2534 1426 2587 1460
rect 2534 1392 2542 1426
rect 2576 1392 2587 1426
rect 2534 1358 2587 1392
rect 2534 1324 2542 1358
rect 2576 1324 2587 1358
rect 2534 1290 2587 1324
rect 2534 1256 2542 1290
rect 2576 1256 2587 1290
rect 2534 1244 2587 1256
rect 2687 1766 2743 1844
rect 2687 1732 2698 1766
rect 2732 1732 2743 1766
rect 2687 1698 2743 1732
rect 2687 1664 2698 1698
rect 2732 1664 2743 1698
rect 2687 1630 2743 1664
rect 2687 1596 2698 1630
rect 2732 1596 2743 1630
rect 2687 1562 2743 1596
rect 2687 1528 2698 1562
rect 2732 1528 2743 1562
rect 2687 1494 2743 1528
rect 2687 1460 2698 1494
rect 2732 1460 2743 1494
rect 2687 1426 2743 1460
rect 2687 1392 2698 1426
rect 2732 1392 2743 1426
rect 2687 1358 2743 1392
rect 2687 1324 2698 1358
rect 2732 1324 2743 1358
rect 2687 1290 2743 1324
rect 2687 1256 2698 1290
rect 2732 1256 2743 1290
rect 2687 1244 2743 1256
rect 2843 1766 2899 1844
rect 2843 1732 2854 1766
rect 2888 1732 2899 1766
rect 2843 1698 2899 1732
rect 2843 1664 2854 1698
rect 2888 1664 2899 1698
rect 2843 1630 2899 1664
rect 2843 1596 2854 1630
rect 2888 1596 2899 1630
rect 2843 1562 2899 1596
rect 2843 1528 2854 1562
rect 2888 1528 2899 1562
rect 2843 1494 2899 1528
rect 2843 1460 2854 1494
rect 2888 1460 2899 1494
rect 2843 1426 2899 1460
rect 2843 1392 2854 1426
rect 2888 1392 2899 1426
rect 2843 1358 2899 1392
rect 2843 1324 2854 1358
rect 2888 1324 2899 1358
rect 2843 1290 2899 1324
rect 2843 1256 2854 1290
rect 2888 1256 2899 1290
rect 2843 1244 2899 1256
rect 2999 1766 3055 1844
rect 2999 1732 3010 1766
rect 3044 1732 3055 1766
rect 2999 1698 3055 1732
rect 2999 1664 3010 1698
rect 3044 1664 3055 1698
rect 2999 1630 3055 1664
rect 2999 1596 3010 1630
rect 3044 1596 3055 1630
rect 2999 1562 3055 1596
rect 2999 1528 3010 1562
rect 3044 1528 3055 1562
rect 2999 1494 3055 1528
rect 2999 1460 3010 1494
rect 3044 1460 3055 1494
rect 2999 1426 3055 1460
rect 2999 1392 3010 1426
rect 3044 1392 3055 1426
rect 2999 1358 3055 1392
rect 2999 1324 3010 1358
rect 3044 1324 3055 1358
rect 2999 1290 3055 1324
rect 2999 1256 3010 1290
rect 3044 1256 3055 1290
rect 2999 1244 3055 1256
rect 3155 1834 3258 1844
rect 3155 1800 3213 1834
rect 3247 1800 3258 1834
rect 3155 1766 3258 1800
rect 3155 1732 3213 1766
rect 3247 1732 3258 1766
rect 3155 1698 3258 1732
rect 3155 1664 3213 1698
rect 3247 1664 3258 1698
rect 3155 1630 3258 1664
rect 3155 1596 3213 1630
rect 3247 1596 3258 1630
rect 3155 1562 3258 1596
rect 3155 1528 3213 1562
rect 3247 1528 3258 1562
rect 3155 1494 3258 1528
rect 3155 1460 3213 1494
rect 3247 1460 3258 1494
rect 3155 1426 3258 1460
rect 3155 1392 3213 1426
rect 3247 1392 3258 1426
rect 3155 1358 3258 1392
rect 3155 1324 3213 1358
rect 3247 1324 3258 1358
rect 3155 1290 3258 1324
rect 3155 1256 3213 1290
rect 3247 1256 3258 1290
rect 3155 1244 3258 1256
rect 3358 2174 3414 2244
rect 3358 2140 3369 2174
rect 3403 2140 3414 2174
rect 3358 2106 3414 2140
rect 3358 2072 3369 2106
rect 3403 2072 3414 2106
rect 3358 2038 3414 2072
rect 3358 2004 3369 2038
rect 3403 2004 3414 2038
rect 3358 1970 3414 2004
rect 3358 1936 3369 1970
rect 3403 1936 3414 1970
rect 3358 1902 3414 1936
rect 3358 1868 3369 1902
rect 3403 1868 3414 1902
rect 3358 1834 3414 1868
rect 3358 1800 3369 1834
rect 3403 1800 3414 1834
rect 3358 1766 3414 1800
rect 3358 1732 3369 1766
rect 3403 1732 3414 1766
rect 3358 1698 3414 1732
rect 3358 1664 3369 1698
rect 3403 1664 3414 1698
rect 3358 1630 3414 1664
rect 3358 1596 3369 1630
rect 3403 1596 3414 1630
rect 3358 1562 3414 1596
rect 3358 1528 3369 1562
rect 3403 1528 3414 1562
rect 3358 1494 3414 1528
rect 3358 1460 3369 1494
rect 3403 1460 3414 1494
rect 3358 1426 3414 1460
rect 3358 1392 3369 1426
rect 3403 1392 3414 1426
rect 3358 1358 3414 1392
rect 3358 1324 3369 1358
rect 3403 1324 3414 1358
rect 3358 1290 3414 1324
rect 3358 1256 3369 1290
rect 3403 1256 3414 1290
rect 3358 1244 3414 1256
rect 3514 2174 3567 2244
rect 3514 2140 3525 2174
rect 3559 2140 3567 2174
rect 3514 2106 3567 2140
rect 3514 2072 3525 2106
rect 3559 2072 3567 2106
rect 3514 2038 3567 2072
rect 3514 2004 3525 2038
rect 3559 2004 3567 2038
rect 3514 1970 3567 2004
rect 3514 1936 3525 1970
rect 3559 1936 3567 1970
rect 3514 1902 3567 1936
rect 3514 1868 3525 1902
rect 3559 1868 3567 1902
rect 3514 1834 3567 1868
rect 3514 1800 3525 1834
rect 3559 1800 3567 1834
rect 3514 1766 3567 1800
rect 3514 1732 3525 1766
rect 3559 1732 3567 1766
rect 3514 1698 3567 1732
rect 3514 1664 3525 1698
rect 3559 1664 3567 1698
rect 3514 1630 3567 1664
rect 3514 1596 3525 1630
rect 3559 1596 3567 1630
rect 3514 1562 3567 1596
rect 3514 1528 3525 1562
rect 3559 1528 3567 1562
rect 3514 1494 3567 1528
rect 3514 1460 3525 1494
rect 3559 1460 3567 1494
rect 3514 1426 3567 1460
rect 3514 1392 3525 1426
rect 3559 1392 3567 1426
rect 3514 1358 3567 1392
rect 3514 1324 3525 1358
rect 3559 1324 3567 1358
rect 3514 1290 3567 1324
rect 3514 1256 3525 1290
rect 3559 1256 3567 1290
rect 3514 1244 3567 1256
<< mvndiffc >>
rect 215 1162 249 1196
rect 215 1094 249 1128
rect 215 1026 249 1060
rect 438 1130 472 1164
rect 438 1062 472 1096
rect 438 994 472 1028
rect 438 926 472 960
rect 902 1130 936 1164
rect 902 1062 936 1096
rect 902 994 936 1028
rect 1012 1028 1046 1062
rect 1868 1028 1902 1062
rect 3524 1028 3558 1062
rect 902 926 936 960
rect 269 708 303 742
rect 269 640 303 674
rect 269 572 303 606
rect 269 504 303 538
rect 269 436 303 470
rect 269 368 303 402
rect 269 300 303 334
rect 269 232 303 266
rect 425 708 459 742
rect 425 640 459 674
rect 425 572 459 606
rect 425 504 459 538
rect 425 436 459 470
rect 425 368 459 402
rect 425 300 459 334
rect 425 232 459 266
rect 581 708 615 742
rect 581 640 615 674
rect 581 572 615 606
rect 581 504 615 538
rect 581 436 615 470
rect 581 368 615 402
rect 581 300 615 334
rect 581 232 615 266
rect 737 708 771 742
rect 737 640 771 674
rect 737 572 771 606
rect 737 504 771 538
rect 737 436 771 470
rect 737 368 771 402
rect 737 300 771 334
rect 737 232 771 266
rect 893 708 927 742
rect 893 640 927 674
rect 893 572 927 606
rect 893 504 927 538
rect 893 436 927 470
rect 893 368 927 402
rect 893 300 927 334
rect 893 232 927 266
rect 1003 708 1037 742
rect 1003 640 1037 674
rect 1003 572 1037 606
rect 1003 504 1037 538
rect 1003 436 1037 470
rect 1003 368 1037 402
rect 1003 300 1037 334
rect 1003 232 1037 266
rect 1159 708 1193 742
rect 1159 640 1193 674
rect 1159 572 1193 606
rect 1159 504 1193 538
rect 1159 436 1193 470
rect 1159 368 1193 402
rect 1159 300 1193 334
rect 1159 232 1193 266
rect 1315 708 1349 742
rect 1315 640 1349 674
rect 1315 572 1349 606
rect 1315 504 1349 538
rect 1315 436 1349 470
rect 1315 368 1349 402
rect 1315 300 1349 334
rect 1315 232 1349 266
rect 1471 708 1505 742
rect 1471 640 1505 674
rect 1471 572 1505 606
rect 1471 504 1505 538
rect 1471 436 1505 470
rect 1471 368 1505 402
rect 1471 300 1505 334
rect 1471 232 1505 266
rect 1627 708 1661 742
rect 1627 640 1661 674
rect 1627 572 1661 606
rect 1627 504 1661 538
rect 1627 436 1661 470
rect 1627 368 1661 402
rect 1627 300 1661 334
rect 1627 232 1661 266
rect 1783 708 1817 742
rect 1783 640 1817 674
rect 1783 572 1817 606
rect 1783 504 1817 538
rect 1783 436 1817 470
rect 1783 368 1817 402
rect 1783 300 1817 334
rect 1783 232 1817 266
rect 1939 708 1973 742
rect 1939 640 1973 674
rect 1939 572 1973 606
rect 1939 504 1973 538
rect 1939 436 1973 470
rect 1939 368 1973 402
rect 1939 300 1973 334
rect 1939 232 1973 266
rect 2095 708 2129 742
rect 2095 640 2129 674
rect 2095 572 2129 606
rect 2095 504 2129 538
rect 2095 436 2129 470
rect 2095 368 2129 402
rect 2095 300 2129 334
rect 2095 232 2129 266
rect 2251 708 2285 742
rect 2251 640 2285 674
rect 2251 572 2285 606
rect 2251 504 2285 538
rect 2251 436 2285 470
rect 2251 368 2285 402
rect 2251 300 2285 334
rect 2251 232 2285 266
rect 2407 708 2441 742
rect 2407 640 2441 674
rect 2407 572 2441 606
rect 2407 504 2441 538
rect 2407 436 2441 470
rect 2407 368 2441 402
rect 2407 300 2441 334
rect 2407 232 2441 266
rect 2563 708 2597 742
rect 2563 640 2597 674
rect 2563 572 2597 606
rect 2563 504 2597 538
rect 2563 436 2597 470
rect 2563 368 2597 402
rect 2563 300 2597 334
rect 2563 232 2597 266
rect 2719 708 2753 742
rect 2719 640 2753 674
rect 2719 572 2753 606
rect 2719 504 2753 538
rect 2719 436 2753 470
rect 2719 368 2753 402
rect 2719 300 2753 334
rect 2719 232 2753 266
rect 2829 708 2863 742
rect 2829 640 2863 674
rect 2829 572 2863 606
rect 2829 504 2863 538
rect 2829 436 2863 470
rect 2829 368 2863 402
rect 2829 300 2863 334
rect 2829 232 2863 266
rect 2985 708 3019 742
rect 2985 640 3019 674
rect 2985 572 3019 606
rect 2985 504 3019 538
rect 2985 436 3019 470
rect 2985 368 3019 402
rect 2985 300 3019 334
rect 2985 232 3019 266
rect 3141 708 3175 742
rect 3141 640 3175 674
rect 3141 572 3175 606
rect 3141 504 3175 538
rect 3141 436 3175 470
rect 3141 368 3175 402
rect 3141 300 3175 334
rect 3141 232 3175 266
rect 3297 708 3331 742
rect 3297 640 3331 674
rect 3297 572 3331 606
rect 3297 504 3331 538
rect 3297 436 3331 470
rect 3297 368 3331 402
rect 3297 300 3331 334
rect 3297 232 3331 266
rect 3453 708 3487 742
rect 3453 640 3487 674
rect 3453 572 3487 606
rect 3453 504 3487 538
rect 3453 436 3487 470
rect 3453 368 3487 402
rect 3453 300 3487 334
rect 3453 232 3487 266
<< mvpdiffc >>
rect 105 2046 139 2080
rect 105 1978 139 2012
rect 105 1910 139 1944
rect 261 2046 295 2080
rect 261 1978 295 2012
rect 261 1910 295 1944
rect 417 2046 451 2080
rect 417 1978 451 2012
rect 417 1910 451 1944
rect 573 2046 607 2080
rect 573 1978 607 2012
rect 573 1910 607 1944
rect 729 2046 763 2080
rect 2432 2026 2466 2060
rect 729 1978 763 2012
rect 729 1910 763 1944
rect 3213 2140 3247 2174
rect 3213 2072 3247 2106
rect 3213 2004 3247 2038
rect 3213 1936 3247 1970
rect 3213 1868 3247 1902
rect 2276 1732 2310 1766
rect 2276 1664 2310 1698
rect 105 1545 139 1579
rect 105 1477 139 1511
rect 105 1409 139 1443
rect 261 1545 295 1579
rect 261 1477 295 1511
rect 261 1409 295 1443
rect 438 1545 472 1579
rect 438 1477 472 1511
rect 438 1409 472 1443
rect 654 1545 688 1579
rect 654 1477 688 1511
rect 654 1409 688 1443
rect 870 1545 904 1579
rect 870 1477 904 1511
rect 870 1409 904 1443
rect 1086 1545 1120 1579
rect 1086 1477 1120 1511
rect 1086 1409 1120 1443
rect 1302 1545 1336 1579
rect 1302 1477 1336 1511
rect 1302 1409 1336 1443
rect 1518 1545 1552 1579
rect 1518 1477 1552 1511
rect 1518 1409 1552 1443
rect 1734 1545 1768 1579
rect 1734 1477 1768 1511
rect 1734 1409 1768 1443
rect 1950 1545 1984 1579
rect 1950 1477 1984 1511
rect 1950 1409 1984 1443
rect 2166 1545 2200 1579
rect 2166 1477 2200 1511
rect 2166 1409 2200 1443
rect 2276 1596 2310 1630
rect 2276 1528 2310 1562
rect 2276 1460 2310 1494
rect 2276 1392 2310 1426
rect 2276 1324 2310 1358
rect 2276 1256 2310 1290
rect 2432 1732 2466 1766
rect 2432 1664 2466 1698
rect 2432 1596 2466 1630
rect 2432 1528 2466 1562
rect 2432 1460 2466 1494
rect 2432 1392 2466 1426
rect 2432 1324 2466 1358
rect 2432 1256 2466 1290
rect 2542 1732 2576 1766
rect 2542 1664 2576 1698
rect 2542 1596 2576 1630
rect 2542 1528 2576 1562
rect 2542 1460 2576 1494
rect 2542 1392 2576 1426
rect 2542 1324 2576 1358
rect 2542 1256 2576 1290
rect 2698 1732 2732 1766
rect 2698 1664 2732 1698
rect 2698 1596 2732 1630
rect 2698 1528 2732 1562
rect 2698 1460 2732 1494
rect 2698 1392 2732 1426
rect 2698 1324 2732 1358
rect 2698 1256 2732 1290
rect 2854 1732 2888 1766
rect 2854 1664 2888 1698
rect 2854 1596 2888 1630
rect 2854 1528 2888 1562
rect 2854 1460 2888 1494
rect 2854 1392 2888 1426
rect 2854 1324 2888 1358
rect 2854 1256 2888 1290
rect 3010 1732 3044 1766
rect 3010 1664 3044 1698
rect 3010 1596 3044 1630
rect 3010 1528 3044 1562
rect 3010 1460 3044 1494
rect 3010 1392 3044 1426
rect 3010 1324 3044 1358
rect 3010 1256 3044 1290
rect 3213 1800 3247 1834
rect 3213 1732 3247 1766
rect 3213 1664 3247 1698
rect 3213 1596 3247 1630
rect 3213 1528 3247 1562
rect 3213 1460 3247 1494
rect 3213 1392 3247 1426
rect 3213 1324 3247 1358
rect 3213 1256 3247 1290
rect 3369 2140 3403 2174
rect 3369 2072 3403 2106
rect 3369 2004 3403 2038
rect 3369 1936 3403 1970
rect 3369 1868 3403 1902
rect 3369 1800 3403 1834
rect 3369 1732 3403 1766
rect 3369 1664 3403 1698
rect 3369 1596 3403 1630
rect 3369 1528 3403 1562
rect 3369 1460 3403 1494
rect 3369 1392 3403 1426
rect 3369 1324 3403 1358
rect 3369 1256 3403 1290
rect 3525 2140 3559 2174
rect 3525 2072 3559 2106
rect 3525 2004 3559 2038
rect 3525 1936 3559 1970
rect 3525 1868 3559 1902
rect 3525 1800 3559 1834
rect 3525 1732 3559 1766
rect 3525 1664 3559 1698
rect 3525 1596 3559 1630
rect 3525 1528 3559 1562
rect 3525 1460 3559 1494
rect 3525 1392 3559 1426
rect 3525 1324 3559 1358
rect 3525 1256 3559 1290
<< mvpsubdiff >>
rect 3569 796 3607 820
rect 3569 762 3571 796
rect 3605 762 3607 796
rect 3569 728 3607 762
rect 3569 694 3571 728
rect 3605 694 3607 728
rect 3569 660 3607 694
rect 3569 626 3571 660
rect 3605 626 3607 660
rect 3569 592 3607 626
rect 3569 558 3571 592
rect 3605 558 3607 592
rect 3569 524 3607 558
rect 3569 490 3571 524
rect 3605 490 3607 524
rect 3569 456 3607 490
rect 3569 422 3571 456
rect 3605 422 3607 456
rect 3569 388 3607 422
rect 3569 354 3571 388
rect 3605 354 3607 388
rect 3569 320 3607 354
rect 3569 286 3571 320
rect 3605 286 3607 320
rect 3569 252 3607 286
rect 3569 218 3571 252
rect 3605 218 3607 252
rect 3569 184 3607 218
rect 3569 150 3571 184
rect 3605 150 3607 184
rect 3569 75 3607 150
rect 149 72 3607 75
rect 149 38 193 72
rect 227 38 261 72
rect 295 38 329 72
rect 363 38 397 72
rect 431 38 465 72
rect 499 38 533 72
rect 567 38 601 72
rect 635 38 669 72
rect 703 38 737 72
rect 771 38 805 72
rect 839 38 873 72
rect 907 38 941 72
rect 975 38 1009 72
rect 1043 38 1077 72
rect 1111 38 1145 72
rect 1179 38 1213 72
rect 1247 38 1281 72
rect 1315 38 1349 72
rect 1383 38 1417 72
rect 1451 38 1485 72
rect 1519 38 1553 72
rect 1587 38 1621 72
rect 1655 38 1689 72
rect 1723 38 1757 72
rect 1791 38 1825 72
rect 1859 38 1893 72
rect 1927 38 1961 72
rect 1995 38 2029 72
rect 2063 38 2097 72
rect 2131 38 2165 72
rect 2199 38 2233 72
rect 2267 38 2301 72
rect 2335 38 2369 72
rect 2403 38 2437 72
rect 2471 38 2505 72
rect 2539 38 2573 72
rect 2607 38 2641 72
rect 2675 38 2709 72
rect 2743 38 2777 72
rect 2811 38 2845 72
rect 2879 38 2913 72
rect 2947 38 2981 72
rect 3015 38 3049 72
rect 3083 38 3117 72
rect 3151 38 3185 72
rect 3219 38 3253 72
rect 3287 38 3321 72
rect 3355 38 3389 72
rect 3423 38 3457 72
rect 3491 38 3525 72
rect 3559 38 3607 72
rect 149 36 3607 38
<< mvnsubdiff >>
rect 92 2281 3098 2283
rect 92 2247 116 2281
rect 150 2247 184 2281
rect 218 2247 252 2281
rect 286 2247 320 2281
rect 354 2247 388 2281
rect 422 2247 456 2281
rect 490 2247 524 2281
rect 558 2247 592 2281
rect 626 2247 660 2281
rect 694 2247 728 2281
rect 762 2247 796 2281
rect 830 2247 864 2281
rect 898 2247 932 2281
rect 966 2247 1000 2281
rect 1034 2247 1068 2281
rect 1102 2247 1136 2281
rect 1170 2247 1204 2281
rect 1238 2247 1272 2281
rect 1306 2247 1340 2281
rect 1374 2247 1408 2281
rect 1442 2247 1476 2281
rect 1510 2247 1544 2281
rect 1578 2247 1612 2281
rect 1646 2247 1680 2281
rect 1714 2247 1748 2281
rect 1782 2247 1816 2281
rect 1850 2247 1884 2281
rect 1918 2247 1952 2281
rect 1986 2247 2020 2281
rect 2054 2247 2088 2281
rect 2122 2247 2156 2281
rect 2190 2247 2224 2281
rect 2258 2247 2292 2281
rect 2326 2247 2360 2281
rect 2394 2247 2428 2281
rect 2462 2247 2496 2281
rect 2530 2247 2564 2281
rect 2598 2247 2632 2281
rect 2666 2247 2700 2281
rect 2734 2247 2768 2281
rect 2802 2247 2836 2281
rect 2870 2247 2904 2281
rect 2938 2247 2972 2281
rect 3006 2247 3040 2281
rect 3074 2247 3098 2281
rect 92 2245 3098 2247
rect 2608 2158 3098 2245
rect 2608 1988 2632 2158
rect 3074 1988 3098 2158
rect 2608 1964 3098 1988
rect 867 1864 1561 1888
rect 867 1762 891 1864
rect 1537 1762 1561 1864
rect 867 1738 1561 1762
<< mvpsubdiffcont >>
rect 3571 762 3605 796
rect 3571 694 3605 728
rect 3571 626 3605 660
rect 3571 558 3605 592
rect 3571 490 3605 524
rect 3571 422 3605 456
rect 3571 354 3605 388
rect 3571 286 3605 320
rect 3571 218 3605 252
rect 3571 150 3605 184
rect 193 38 227 72
rect 261 38 295 72
rect 329 38 363 72
rect 397 38 431 72
rect 465 38 499 72
rect 533 38 567 72
rect 601 38 635 72
rect 669 38 703 72
rect 737 38 771 72
rect 805 38 839 72
rect 873 38 907 72
rect 941 38 975 72
rect 1009 38 1043 72
rect 1077 38 1111 72
rect 1145 38 1179 72
rect 1213 38 1247 72
rect 1281 38 1315 72
rect 1349 38 1383 72
rect 1417 38 1451 72
rect 1485 38 1519 72
rect 1553 38 1587 72
rect 1621 38 1655 72
rect 1689 38 1723 72
rect 1757 38 1791 72
rect 1825 38 1859 72
rect 1893 38 1927 72
rect 1961 38 1995 72
rect 2029 38 2063 72
rect 2097 38 2131 72
rect 2165 38 2199 72
rect 2233 38 2267 72
rect 2301 38 2335 72
rect 2369 38 2403 72
rect 2437 38 2471 72
rect 2505 38 2539 72
rect 2573 38 2607 72
rect 2641 38 2675 72
rect 2709 38 2743 72
rect 2777 38 2811 72
rect 2845 38 2879 72
rect 2913 38 2947 72
rect 2981 38 3015 72
rect 3049 38 3083 72
rect 3117 38 3151 72
rect 3185 38 3219 72
rect 3253 38 3287 72
rect 3321 38 3355 72
rect 3389 38 3423 72
rect 3457 38 3491 72
rect 3525 38 3559 72
<< mvnsubdiffcont >>
rect 116 2247 150 2281
rect 184 2247 218 2281
rect 252 2247 286 2281
rect 320 2247 354 2281
rect 388 2247 422 2281
rect 456 2247 490 2281
rect 524 2247 558 2281
rect 592 2247 626 2281
rect 660 2247 694 2281
rect 728 2247 762 2281
rect 796 2247 830 2281
rect 864 2247 898 2281
rect 932 2247 966 2281
rect 1000 2247 1034 2281
rect 1068 2247 1102 2281
rect 1136 2247 1170 2281
rect 1204 2247 1238 2281
rect 1272 2247 1306 2281
rect 1340 2247 1374 2281
rect 1408 2247 1442 2281
rect 1476 2247 1510 2281
rect 1544 2247 1578 2281
rect 1612 2247 1646 2281
rect 1680 2247 1714 2281
rect 1748 2247 1782 2281
rect 1816 2247 1850 2281
rect 1884 2247 1918 2281
rect 1952 2247 1986 2281
rect 2020 2247 2054 2281
rect 2088 2247 2122 2281
rect 2156 2247 2190 2281
rect 2224 2247 2258 2281
rect 2292 2247 2326 2281
rect 2360 2247 2394 2281
rect 2428 2247 2462 2281
rect 2496 2247 2530 2281
rect 2564 2247 2598 2281
rect 2632 2247 2666 2281
rect 2700 2247 2734 2281
rect 2768 2247 2802 2281
rect 2836 2247 2870 2281
rect 2904 2247 2938 2281
rect 2972 2247 3006 2281
rect 3040 2247 3074 2281
rect 2632 1988 3074 2158
rect 891 1762 1537 1864
<< poly >>
rect 445 2191 579 2207
rect 445 2157 461 2191
rect 495 2157 529 2191
rect 563 2157 579 2191
rect 445 2141 579 2157
rect 3258 2244 3358 2270
rect 3414 2244 3514 2270
rect 150 2098 250 2124
rect 306 2098 406 2124
rect 462 2098 562 2141
rect 618 2098 718 2124
rect 821 2098 2421 2124
rect 821 1988 2421 2014
rect 821 1966 2187 1988
rect 821 1932 841 1966
rect 875 1932 909 1966
rect 943 1932 977 1966
rect 1011 1932 1045 1966
rect 1079 1932 1113 1966
rect 1147 1932 1181 1966
rect 1215 1932 1249 1966
rect 1283 1932 1317 1966
rect 1351 1932 1385 1966
rect 1419 1932 1453 1966
rect 1487 1932 1521 1966
rect 1555 1932 1589 1966
rect 1623 1932 1657 1966
rect 1691 1932 1725 1966
rect 1759 1932 1793 1966
rect 1827 1932 1861 1966
rect 1895 1932 1929 1966
rect 1963 1932 1997 1966
rect 2031 1932 2065 1966
rect 2099 1932 2133 1966
rect 2167 1932 2187 1966
rect 821 1912 2187 1932
rect 2280 1926 2421 1942
rect 150 1850 250 1898
rect 150 1816 184 1850
rect 218 1816 250 1850
rect 150 1782 250 1816
rect 150 1748 184 1782
rect 218 1748 250 1782
rect 150 1714 250 1748
rect 306 1850 406 1898
rect 462 1872 562 1898
rect 306 1816 340 1850
rect 374 1816 406 1850
rect 618 1847 718 1898
rect 2280 1892 2296 1926
rect 2330 1892 2364 1926
rect 2398 1892 2421 1926
rect 2280 1876 2421 1892
rect 306 1782 406 1816
rect 306 1748 340 1782
rect 374 1748 406 1782
rect 600 1831 734 1847
rect 600 1797 616 1831
rect 650 1797 684 1831
rect 718 1797 734 1831
rect 600 1781 734 1797
rect 306 1732 406 1748
rect 2321 1844 2421 1876
rect 2587 1926 3155 1946
rect 2587 1892 2614 1926
rect 2648 1892 2682 1926
rect 2716 1892 2750 1926
rect 2784 1892 2818 1926
rect 2852 1892 2886 1926
rect 2920 1892 2954 1926
rect 2988 1892 3022 1926
rect 3056 1892 3090 1926
rect 3124 1892 3155 1926
rect 2587 1870 3155 1892
rect 2587 1844 2687 1870
rect 2743 1844 2843 1870
rect 2899 1844 2999 1870
rect 3055 1844 3155 1870
rect 150 1680 184 1714
rect 218 1690 250 1714
rect 218 1680 406 1690
rect 150 1623 406 1680
rect 150 1597 250 1623
rect 306 1597 406 1623
rect 483 1679 2155 1695
rect 483 1645 527 1679
rect 561 1645 595 1679
rect 629 1645 663 1679
rect 697 1645 731 1679
rect 765 1645 982 1679
rect 1016 1645 1050 1679
rect 1084 1645 1118 1679
rect 1152 1645 1186 1679
rect 1220 1645 1483 1679
rect 1517 1645 1551 1679
rect 1585 1645 2155 1679
rect 483 1623 2155 1645
rect 483 1597 643 1623
rect 699 1597 859 1623
rect 915 1597 1075 1623
rect 1131 1597 1291 1623
rect 1347 1597 1507 1623
rect 1563 1597 1723 1623
rect 1779 1597 1939 1623
rect 1995 1597 2155 1623
rect 150 1371 250 1397
rect 306 1371 406 1397
rect 483 1371 643 1397
rect 699 1371 859 1397
rect 915 1371 1075 1397
rect 1131 1371 1291 1397
rect 1347 1371 1507 1397
rect 1563 1371 1723 1397
rect 1779 1371 1939 1397
rect 1995 1371 2155 1397
rect 150 1240 380 1371
rect 620 1313 754 1329
rect 423 1296 578 1312
rect 423 1262 460 1296
rect 494 1262 528 1296
rect 562 1262 578 1296
rect 620 1279 636 1313
rect 670 1279 704 1313
rect 738 1279 754 1313
rect 620 1263 754 1279
rect 796 1296 951 1312
rect 423 1240 578 1262
rect 260 1214 380 1240
rect 483 1214 583 1240
rect 637 1214 737 1263
rect 796 1262 812 1296
rect 846 1262 880 1296
rect 914 1262 951 1296
rect 796 1240 951 1262
rect 1131 1303 1833 1371
rect 1131 1269 1294 1303
rect 1328 1269 1362 1303
rect 1396 1269 1430 1303
rect 1464 1269 1498 1303
rect 1532 1269 1566 1303
rect 1600 1269 1634 1303
rect 1668 1269 1702 1303
rect 1736 1269 1770 1303
rect 1804 1269 1833 1303
rect 791 1214 891 1240
rect 1131 1224 1833 1269
rect 260 988 380 1014
rect 1131 1122 1158 1224
rect 1804 1122 1833 1224
rect 2321 1218 2421 1244
rect 2587 1218 2687 1244
rect 2743 1218 2843 1244
rect 2899 1218 2999 1244
rect 3055 1218 3155 1244
rect 3258 1218 3358 1244
rect 3414 1218 3514 1244
rect 3197 1196 3575 1218
rect 1131 1100 1833 1122
rect 1913 1156 3155 1172
rect 1913 1122 1982 1156
rect 2016 1122 2050 1156
rect 2084 1122 2118 1156
rect 2152 1122 2186 1156
rect 2220 1122 2254 1156
rect 2288 1122 2322 1156
rect 2356 1122 2390 1156
rect 2424 1122 2458 1156
rect 2492 1122 2526 1156
rect 2560 1122 3155 1156
rect 3197 1162 3217 1196
rect 3251 1162 3285 1196
rect 3319 1162 3453 1196
rect 3487 1162 3521 1196
rect 3555 1162 3575 1196
rect 3197 1142 3575 1162
rect 1913 1100 3155 1122
rect 1057 1074 1857 1100
rect 1913 1074 3513 1100
rect 1057 964 1857 990
rect 1913 964 3513 990
rect 483 888 583 914
rect 637 888 737 914
rect 791 888 891 914
rect 1672 902 2240 922
rect 1672 868 1702 902
rect 1736 868 1770 902
rect 1804 868 1838 902
rect 1872 868 1906 902
rect 1940 868 1974 902
rect 2008 868 2042 902
rect 2076 868 2110 902
rect 2144 868 2178 902
rect 2212 868 2240 902
rect 1672 846 2240 868
rect 314 820 414 846
rect 470 820 570 846
rect 626 820 726 846
rect 782 820 882 846
rect 1048 820 1148 846
rect 1204 820 1304 846
rect 1360 820 1460 846
rect 1516 820 1616 846
rect 1672 820 1772 846
rect 1828 820 1928 846
rect 1984 820 2084 846
rect 2140 820 2240 846
rect 2296 820 2396 846
rect 2452 820 2552 846
rect 2608 820 2708 846
rect 2874 820 2974 846
rect 3030 820 3130 846
rect 3186 820 3286 846
rect 3342 820 3442 846
rect 314 194 414 220
rect 470 194 570 220
rect 626 194 726 220
rect 782 194 882 220
rect 314 172 882 194
rect 314 138 344 172
rect 378 138 412 172
rect 446 138 480 172
rect 514 138 548 172
rect 582 138 616 172
rect 650 138 684 172
rect 718 138 752 172
rect 786 138 820 172
rect 854 138 882 172
rect 314 118 882 138
rect 1048 194 1148 220
rect 1204 194 1304 220
rect 1360 194 1460 220
rect 1516 194 1616 220
rect 1672 194 1772 220
rect 1828 194 1928 220
rect 1984 194 2084 220
rect 2140 194 2240 220
rect 1048 172 1616 194
rect 2296 173 2396 220
rect 2452 194 2552 220
rect 2608 194 2708 220
rect 1048 138 1078 172
rect 1112 138 1146 172
rect 1180 138 1214 172
rect 1248 138 1282 172
rect 1316 138 1350 172
rect 1384 138 1418 172
rect 1452 138 1486 172
rect 1520 138 1554 172
rect 1588 138 1616 172
rect 1048 118 1616 138
rect 2279 157 2413 173
rect 2279 123 2295 157
rect 2329 123 2363 157
rect 2397 123 2413 157
rect 2279 107 2413 123
rect 2467 172 2708 194
rect 2467 138 2491 172
rect 2525 138 2559 172
rect 2593 138 2627 172
rect 2661 138 2708 172
rect 2467 118 2708 138
rect 2874 194 2974 220
rect 3030 194 3130 220
rect 2874 172 3130 194
rect 2874 138 2910 172
rect 2944 138 2978 172
rect 3012 138 3046 172
rect 3080 138 3130 172
rect 2874 118 3130 138
rect 3186 194 3286 220
rect 3342 194 3442 220
rect 3186 172 3442 194
rect 3186 138 3222 172
rect 3256 138 3290 172
rect 3324 138 3358 172
rect 3392 138 3442 172
rect 3186 118 3442 138
<< polycont >>
rect 461 2157 495 2191
rect 529 2157 563 2191
rect 841 1932 875 1966
rect 909 1932 943 1966
rect 977 1932 1011 1966
rect 1045 1932 1079 1966
rect 1113 1932 1147 1966
rect 1181 1932 1215 1966
rect 1249 1932 1283 1966
rect 1317 1932 1351 1966
rect 1385 1932 1419 1966
rect 1453 1932 1487 1966
rect 1521 1932 1555 1966
rect 1589 1932 1623 1966
rect 1657 1932 1691 1966
rect 1725 1932 1759 1966
rect 1793 1932 1827 1966
rect 1861 1932 1895 1966
rect 1929 1932 1963 1966
rect 1997 1932 2031 1966
rect 2065 1932 2099 1966
rect 2133 1932 2167 1966
rect 184 1816 218 1850
rect 184 1748 218 1782
rect 340 1816 374 1850
rect 2296 1892 2330 1926
rect 2364 1892 2398 1926
rect 340 1748 374 1782
rect 616 1797 650 1831
rect 684 1797 718 1831
rect 2614 1892 2648 1926
rect 2682 1892 2716 1926
rect 2750 1892 2784 1926
rect 2818 1892 2852 1926
rect 2886 1892 2920 1926
rect 2954 1892 2988 1926
rect 3022 1892 3056 1926
rect 3090 1892 3124 1926
rect 184 1680 218 1714
rect 527 1645 561 1679
rect 595 1645 629 1679
rect 663 1645 697 1679
rect 731 1645 765 1679
rect 982 1645 1016 1679
rect 1050 1645 1084 1679
rect 1118 1645 1152 1679
rect 1186 1645 1220 1679
rect 1483 1645 1517 1679
rect 1551 1645 1585 1679
rect 460 1262 494 1296
rect 528 1262 562 1296
rect 636 1279 670 1313
rect 704 1279 738 1313
rect 812 1262 846 1296
rect 880 1262 914 1296
rect 1294 1269 1328 1303
rect 1362 1269 1396 1303
rect 1430 1269 1464 1303
rect 1498 1269 1532 1303
rect 1566 1269 1600 1303
rect 1634 1269 1668 1303
rect 1702 1269 1736 1303
rect 1770 1269 1804 1303
rect 1158 1122 1804 1224
rect 1982 1122 2016 1156
rect 2050 1122 2084 1156
rect 2118 1122 2152 1156
rect 2186 1122 2220 1156
rect 2254 1122 2288 1156
rect 2322 1122 2356 1156
rect 2390 1122 2424 1156
rect 2458 1122 2492 1156
rect 2526 1122 2560 1156
rect 3217 1162 3251 1196
rect 3285 1162 3319 1196
rect 3453 1162 3487 1196
rect 3521 1162 3555 1196
rect 1702 868 1736 902
rect 1770 868 1804 902
rect 1838 868 1872 902
rect 1906 868 1940 902
rect 1974 868 2008 902
rect 2042 868 2076 902
rect 2110 868 2144 902
rect 2178 868 2212 902
rect 344 138 378 172
rect 412 138 446 172
rect 480 138 514 172
rect 548 138 582 172
rect 616 138 650 172
rect 684 138 718 172
rect 752 138 786 172
rect 820 138 854 172
rect 1078 138 1112 172
rect 1146 138 1180 172
rect 1214 138 1248 172
rect 1282 138 1316 172
rect 1350 138 1384 172
rect 1418 138 1452 172
rect 1486 138 1520 172
rect 1554 138 1588 172
rect 2295 123 2329 157
rect 2363 123 2397 157
rect 2491 138 2525 172
rect 2559 138 2593 172
rect 2627 138 2661 172
rect 2910 138 2944 172
rect 2978 138 3012 172
rect 3046 138 3080 172
rect 3222 138 3256 172
rect 3290 138 3324 172
rect 3358 138 3392 172
<< locali >>
rect 100 2259 116 2281
rect 100 2247 115 2259
rect 150 2247 184 2281
rect 218 2259 252 2281
rect 286 2259 320 2281
rect 354 2259 388 2281
rect 422 2259 456 2281
rect 490 2259 524 2281
rect 558 2259 592 2281
rect 626 2259 660 2281
rect 694 2259 728 2281
rect 221 2247 252 2259
rect 105 2225 115 2247
rect 149 2225 187 2247
rect 221 2225 259 2247
rect 293 2225 305 2259
rect 437 2247 456 2259
rect 509 2247 524 2259
rect 581 2247 592 2259
rect 653 2247 660 2259
rect 725 2247 728 2259
rect 762 2259 796 2281
rect 830 2259 864 2281
rect 898 2259 932 2281
rect 966 2259 1000 2281
rect 1034 2259 1068 2281
rect 1102 2259 1136 2281
rect 1170 2259 1204 2281
rect 1238 2259 1272 2281
rect 1306 2259 1340 2281
rect 762 2247 763 2259
rect 830 2247 835 2259
rect 898 2247 907 2259
rect 966 2247 979 2259
rect 1034 2247 1051 2259
rect 1102 2247 1123 2259
rect 1170 2247 1195 2259
rect 1238 2247 1267 2259
rect 1306 2247 1339 2259
rect 1374 2247 1408 2281
rect 1442 2259 1476 2281
rect 1510 2259 1544 2281
rect 1578 2259 1612 2281
rect 1646 2259 1680 2281
rect 1714 2259 1748 2281
rect 1782 2259 1816 2281
rect 1850 2259 1884 2281
rect 1918 2259 1952 2281
rect 1445 2247 1476 2259
rect 1517 2247 1544 2259
rect 1589 2247 1612 2259
rect 1661 2247 1680 2259
rect 1733 2247 1748 2259
rect 1805 2247 1816 2259
rect 1877 2247 1884 2259
rect 1949 2247 1952 2259
rect 1986 2259 2020 2281
rect 2054 2259 2088 2281
rect 2122 2259 2156 2281
rect 2190 2259 2224 2281
rect 2258 2259 2292 2281
rect 2326 2259 2360 2281
rect 2394 2259 2428 2281
rect 2462 2259 2496 2281
rect 2530 2259 2564 2281
rect 1986 2247 1987 2259
rect 2054 2247 2059 2259
rect 2122 2247 2131 2259
rect 2190 2247 2203 2259
rect 2258 2247 2275 2259
rect 2326 2247 2347 2259
rect 2394 2247 2419 2259
rect 2462 2247 2491 2259
rect 2530 2247 2563 2259
rect 2598 2247 2632 2281
rect 2666 2259 2700 2281
rect 2734 2259 2768 2281
rect 2802 2259 2836 2281
rect 2870 2259 2904 2281
rect 2938 2259 2972 2281
rect 3006 2259 3040 2281
rect 3074 2259 3090 2281
rect 2669 2247 2700 2259
rect 2741 2247 2768 2259
rect 2813 2247 2836 2259
rect 2885 2247 2904 2259
rect 2957 2247 2972 2259
rect 3029 2247 3040 2259
rect 437 2225 475 2247
rect 509 2225 547 2247
rect 581 2225 619 2247
rect 653 2225 691 2247
rect 725 2225 763 2247
rect 797 2225 835 2247
rect 869 2225 907 2247
rect 941 2225 979 2247
rect 1013 2225 1051 2247
rect 1085 2225 1123 2247
rect 1157 2225 1195 2247
rect 1229 2225 1267 2247
rect 1301 2225 1339 2247
rect 1373 2225 1411 2247
rect 1445 2225 1483 2247
rect 1517 2225 1555 2247
rect 1589 2225 1627 2247
rect 1661 2225 1699 2247
rect 1733 2225 1771 2247
rect 1805 2225 1843 2247
rect 1877 2225 1915 2247
rect 1949 2225 1987 2247
rect 2021 2225 2059 2247
rect 2093 2225 2131 2247
rect 2165 2225 2203 2247
rect 2237 2225 2275 2247
rect 2309 2225 2347 2247
rect 2381 2225 2419 2247
rect 2453 2225 2491 2247
rect 2525 2225 2563 2247
rect 2597 2225 2635 2247
rect 2669 2225 2707 2247
rect 2741 2225 2779 2247
rect 2813 2225 2851 2247
rect 2885 2225 2923 2247
rect 2957 2225 2995 2247
rect 3029 2225 3067 2247
rect 105 2107 139 2225
rect 445 2157 461 2191
rect 329 2098 411 2153
rect 105 2035 139 2046
rect 105 1944 139 1978
rect 105 1595 139 1910
rect 261 2080 295 2096
rect 261 2012 295 2045
rect 261 1944 295 1973
rect 261 1894 295 1910
rect 329 2080 461 2098
rect 329 2046 417 2080
rect 451 2046 461 2080
rect 329 2012 461 2046
rect 329 1978 417 2012
rect 451 1978 461 2012
rect 329 1944 461 1978
rect 329 1910 417 1944
rect 451 1910 461 1944
rect 329 1906 461 1910
rect 184 1850 218 1866
rect 184 1782 218 1816
rect 340 1850 374 1866
rect 340 1782 374 1816
rect 218 1715 256 1749
rect 184 1714 218 1715
rect 184 1664 218 1680
rect 105 1523 139 1545
rect 105 1451 139 1477
rect 105 1393 139 1409
rect 215 1579 295 1595
rect 215 1545 261 1579
rect 215 1511 295 1545
rect 215 1477 261 1511
rect 215 1443 295 1477
rect 215 1409 261 1443
rect 215 1196 295 1409
rect 340 1296 374 1748
rect 417 1595 461 1906
rect 495 1986 529 2191
rect 563 2157 579 2191
rect 729 2147 763 2225
rect 495 1914 529 1952
rect 573 2080 607 2096
rect 573 2012 607 2046
rect 573 1944 607 1978
rect 729 2080 763 2113
rect 2616 2158 3090 2225
rect 729 2012 763 2041
rect 729 1944 763 1978
rect 2432 2060 2466 2076
rect 2432 1973 2466 2026
rect 2616 1988 2632 2158
rect 3074 1988 3090 2158
rect 3213 2174 3247 2190
rect 3213 2106 3247 2140
rect 3213 2038 3247 2072
rect 573 1902 589 1910
rect 623 1902 661 1936
rect 825 1932 841 1966
rect 875 1932 909 1966
rect 943 1932 977 1966
rect 1011 1932 1045 1966
rect 1079 1932 1113 1966
rect 1147 1932 1181 1966
rect 1215 1932 1249 1966
rect 1283 1932 1317 1966
rect 1351 1932 1385 1966
rect 1419 1932 1453 1966
rect 1487 1932 1521 1966
rect 1555 1932 1589 1966
rect 1623 1932 1657 1966
rect 1691 1932 1725 1966
rect 1759 1932 1793 1966
rect 1827 1932 1861 1966
rect 1895 1932 1929 1966
rect 1963 1932 1997 1966
rect 2031 1932 2065 1966
rect 2099 1932 2133 1966
rect 2167 1932 2183 1966
rect 573 1894 607 1902
rect 729 1894 763 1910
rect 556 1797 616 1831
rect 650 1797 684 1831
rect 718 1797 734 1831
rect 556 1764 662 1797
rect 590 1730 628 1764
rect 858 1762 891 1864
rect 1537 1762 1553 1864
rect 511 1645 527 1679
rect 561 1645 595 1679
rect 629 1645 663 1679
rect 697 1645 731 1679
rect 765 1645 781 1679
rect 417 1545 438 1595
rect 417 1523 472 1545
rect 417 1477 438 1523
rect 417 1451 472 1477
rect 417 1409 438 1451
rect 417 1393 472 1409
rect 654 1579 688 1595
rect 654 1511 688 1545
rect 654 1443 688 1477
rect 654 1381 688 1409
rect 858 1579 932 1762
rect 966 1645 982 1679
rect 1016 1645 1050 1679
rect 1084 1645 1118 1679
rect 1152 1645 1186 1679
rect 1220 1645 1236 1679
rect 858 1477 870 1579
rect 904 1477 932 1579
rect 858 1473 932 1477
rect 858 1409 870 1473
rect 904 1409 932 1473
rect 858 1393 932 1409
rect 1086 1579 1120 1595
rect 1086 1511 1120 1545
rect 1086 1443 1120 1477
rect 688 1347 726 1381
rect 1086 1371 1120 1409
rect 1270 1579 1427 1762
rect 1467 1645 1483 1679
rect 1517 1645 1551 1679
rect 1585 1645 1601 1679
rect 1641 1675 2095 1932
rect 2276 1926 2398 1942
rect 2432 1939 2444 1973
rect 2478 1939 2516 1973
rect 3213 1970 3247 2004
rect 2276 1892 2296 1926
rect 2330 1892 2364 1926
rect 2598 1895 2614 1926
rect 2276 1876 2398 1892
rect 2432 1893 2614 1895
rect 2648 1893 2682 1926
rect 2716 1893 2750 1926
rect 2784 1893 2818 1926
rect 2276 1819 2310 1876
rect 2238 1785 2276 1819
rect 2276 1766 2310 1785
rect 2276 1698 2310 1732
rect 1675 1641 1713 1675
rect 1747 1641 1785 1675
rect 1819 1641 1857 1675
rect 1891 1641 1929 1675
rect 1963 1641 2001 1675
rect 2035 1641 2073 1675
rect 2276 1630 2310 1664
rect 2094 1595 2200 1597
rect 1270 1477 1302 1579
rect 1336 1477 1427 1579
rect 1270 1473 1427 1477
rect 1270 1409 1302 1473
rect 1336 1409 1427 1473
rect 1270 1393 1427 1409
rect 1518 1579 1552 1595
rect 1518 1511 1552 1545
rect 1518 1443 1552 1477
rect 1518 1371 1552 1409
rect 1734 1523 1768 1545
rect 1734 1451 1768 1477
rect 1734 1393 1768 1409
rect 1950 1579 1984 1595
rect 1950 1511 1984 1545
rect 1950 1443 1984 1477
rect 1950 1371 1984 1409
rect 1086 1337 1098 1371
rect 1132 1337 1170 1371
rect 1518 1337 1556 1371
rect 1912 1337 1950 1371
rect 2094 1409 2166 1417
rect 340 1262 456 1296
rect 494 1262 528 1296
rect 562 1262 578 1296
rect 620 1279 636 1313
rect 670 1279 704 1313
rect 738 1296 754 1313
rect 1086 1296 1204 1337
rect 742 1279 754 1296
rect 670 1262 708 1279
rect 796 1262 812 1296
rect 846 1262 880 1296
rect 918 1262 930 1296
rect 1086 1262 1098 1296
rect 1132 1262 1170 1296
rect 1278 1269 1294 1303
rect 1328 1269 1362 1303
rect 1396 1269 1430 1303
rect 1464 1269 1498 1303
rect 1532 1269 1566 1303
rect 1600 1269 1634 1303
rect 1668 1269 1702 1303
rect 1736 1269 1770 1303
rect 1804 1269 1820 1303
rect 249 1162 295 1196
rect 215 1128 295 1162
rect 249 1094 295 1128
rect 215 1060 295 1094
rect 249 1026 295 1060
rect 215 845 295 1026
rect 438 1164 472 1180
rect 438 1096 472 1130
rect 438 1028 472 1035
rect 438 960 472 963
rect 438 925 472 926
rect 902 1175 936 1180
rect 1142 1175 1158 1224
rect 936 1141 974 1175
rect 1008 1141 1046 1175
rect 1080 1141 1118 1175
rect 1152 1141 1158 1175
rect 902 1096 936 1130
rect 1142 1122 1158 1141
rect 1804 1122 1820 1224
rect 2094 1156 2200 1409
rect 2276 1562 2310 1596
rect 2276 1494 2310 1528
rect 2276 1426 2310 1460
rect 2276 1358 2310 1392
rect 2276 1290 2310 1324
rect 2276 1240 2310 1256
rect 2432 1859 2599 1893
rect 2648 1892 2671 1893
rect 2716 1892 2743 1893
rect 2784 1892 2815 1893
rect 2852 1892 2886 1926
rect 2920 1893 2954 1926
rect 2988 1893 3022 1926
rect 3056 1893 3090 1926
rect 3124 1893 3140 1926
rect 2921 1892 2954 1893
rect 2993 1892 3022 1893
rect 3065 1892 3090 1893
rect 3137 1892 3140 1893
rect 3213 1902 3247 1936
rect 2633 1859 2671 1892
rect 2705 1859 2743 1892
rect 2777 1859 2815 1892
rect 2849 1859 2887 1892
rect 2921 1859 2959 1892
rect 2993 1859 3031 1892
rect 3065 1859 3103 1892
rect 2432 1766 2466 1859
rect 3213 1834 3247 1868
rect 2432 1698 2466 1732
rect 2432 1630 2466 1664
rect 2432 1562 2466 1596
rect 2432 1494 2466 1528
rect 2432 1426 2466 1460
rect 2432 1358 2466 1392
rect 2432 1290 2466 1324
rect 2432 1240 2466 1256
rect 2542 1766 2576 1782
rect 2542 1698 2576 1732
rect 2542 1630 2576 1664
rect 2542 1595 2576 1596
rect 2542 1523 2576 1528
rect 2542 1451 2576 1460
rect 2542 1358 2576 1392
rect 2542 1290 2576 1324
rect 2542 1156 2576 1256
rect 2698 1766 2732 1782
rect 2698 1698 2732 1732
rect 2698 1630 2732 1664
rect 2698 1562 2732 1596
rect 2698 1494 2732 1528
rect 2698 1426 2732 1460
rect 2698 1358 2732 1392
rect 2698 1290 2732 1324
rect 2698 1171 2732 1256
rect 2854 1766 2888 1782
rect 2854 1698 2888 1732
rect 2854 1630 2888 1664
rect 2854 1595 2888 1596
rect 2854 1523 2888 1528
rect 2854 1451 2888 1460
rect 2854 1358 2888 1392
rect 2854 1290 2888 1324
rect 2854 1240 2888 1256
rect 3010 1766 3044 1782
rect 3010 1698 3044 1732
rect 3010 1630 3044 1664
rect 3010 1562 3044 1596
rect 3010 1494 3044 1528
rect 3010 1426 3044 1460
rect 3010 1358 3044 1392
rect 3010 1290 3044 1324
rect 3010 1171 3044 1256
rect 3213 1766 3247 1800
rect 3213 1698 3247 1732
rect 3213 1630 3247 1664
rect 3213 1595 3247 1596
rect 3213 1523 3247 1528
rect 3213 1451 3247 1460
rect 3213 1358 3247 1392
rect 3213 1290 3247 1324
rect 3213 1240 3247 1256
rect 3369 2174 3403 2190
rect 3369 2106 3403 2140
rect 3369 2038 3403 2072
rect 3369 1970 3403 2004
rect 3369 1902 3403 1936
rect 3369 1834 3403 1868
rect 3369 1766 3403 1800
rect 3369 1698 3403 1732
rect 3369 1630 3403 1664
rect 3369 1562 3403 1596
rect 3369 1494 3403 1528
rect 3369 1426 3403 1460
rect 3369 1358 3403 1392
rect 3369 1290 3403 1324
rect 1966 1122 1982 1156
rect 2016 1122 2050 1156
rect 2084 1122 2118 1156
rect 2152 1122 2186 1156
rect 2220 1122 2254 1156
rect 2288 1122 2322 1156
rect 2356 1122 2390 1156
rect 2424 1122 2458 1156
rect 2492 1122 2526 1156
rect 2560 1122 2576 1156
rect 2697 1137 2735 1171
rect 2972 1137 3010 1171
rect 3201 1177 3217 1196
rect 3201 1162 3213 1177
rect 3251 1162 3285 1196
rect 3319 1162 3335 1196
rect 3247 1143 3285 1162
rect 902 1028 936 1062
rect 902 960 936 994
rect 902 910 936 926
rect 1012 1062 1046 1078
rect 1012 845 1046 1028
rect 1868 1069 1902 1078
rect 1868 997 1902 1028
rect 3369 941 3403 1256
rect 3525 2174 3559 2190
rect 3525 2106 3559 2140
rect 3525 2038 3559 2072
rect 3525 1970 3559 2004
rect 3525 1902 3559 1936
rect 3525 1834 3559 1868
rect 3525 1766 3559 1800
rect 3525 1698 3559 1732
rect 3525 1630 3559 1664
rect 3525 1595 3559 1596
rect 3525 1523 3559 1528
rect 3525 1451 3559 1460
rect 3525 1358 3559 1392
rect 3525 1290 3559 1324
rect 3525 1240 3559 1256
rect 3437 1162 3453 1196
rect 3487 1162 3521 1196
rect 3555 1177 3571 1196
rect 3559 1162 3571 1177
rect 3487 1143 3525 1162
rect 2985 907 3403 941
rect 3497 1062 3558 1078
rect 3497 1028 3524 1062
rect 3497 1012 3558 1028
rect 1686 868 1702 902
rect 1736 868 1770 902
rect 1804 868 1838 902
rect 1872 868 1906 902
rect 1940 868 1974 902
rect 2008 868 2042 902
rect 2076 868 2110 902
rect 2144 868 2178 902
rect 2212 868 2228 902
rect 1686 845 2228 868
rect 215 831 219 845
rect 253 811 291 845
rect 325 811 363 845
rect 1012 811 1067 845
rect 1101 811 1139 845
rect 1686 833 1687 845
rect 1721 811 1759 845
rect 1793 811 1831 845
rect 1865 811 1903 845
rect 1937 811 1975 845
rect 2009 811 2047 845
rect 2081 811 2119 845
rect 2153 811 2191 845
rect 2225 833 2228 845
rect 2719 811 2728 845
rect 2762 811 2800 845
rect 269 742 303 758
rect 269 685 303 708
rect 425 742 459 758
rect 303 651 341 685
rect 425 674 459 708
rect 581 742 615 758
rect 581 685 615 708
rect 737 742 771 758
rect 269 606 303 640
rect 269 538 303 572
rect 269 470 303 504
rect 269 402 303 436
rect 269 334 303 368
rect 269 266 303 300
rect 269 216 303 232
rect 581 674 619 685
rect 425 606 459 640
rect 425 538 459 572
rect 425 470 459 504
rect 425 402 459 436
rect 425 334 459 368
rect 425 266 459 300
rect 425 172 459 232
rect 615 651 619 674
rect 737 674 771 708
rect 893 742 927 758
rect 893 685 927 708
rect 581 606 615 640
rect 581 538 615 572
rect 581 470 615 504
rect 581 402 615 436
rect 581 334 615 368
rect 581 266 615 300
rect 581 216 615 232
rect 855 651 893 685
rect 737 606 771 640
rect 737 538 771 572
rect 737 470 771 504
rect 737 402 771 436
rect 737 334 771 368
rect 737 266 771 300
rect 737 172 771 232
rect 893 606 927 640
rect 893 538 927 572
rect 893 470 927 504
rect 893 402 927 436
rect 893 334 927 368
rect 893 266 927 300
rect 893 216 927 232
rect 1003 742 1037 758
rect 1003 674 1037 708
rect 1159 742 1193 758
rect 1159 685 1193 708
rect 1315 742 1349 758
rect 1158 674 1196 685
rect 1158 651 1159 674
rect 1003 606 1037 640
rect 1003 538 1037 551
rect 1003 470 1037 479
rect 1003 402 1037 436
rect 1003 334 1037 368
rect 1003 266 1037 300
rect 1003 216 1037 232
rect 1193 651 1196 674
rect 1315 674 1349 708
rect 1471 742 1505 758
rect 1471 685 1505 708
rect 1627 742 1661 758
rect 1159 606 1193 640
rect 1159 538 1193 572
rect 1159 470 1193 504
rect 1159 402 1193 436
rect 1159 334 1193 368
rect 1159 266 1193 300
rect 1159 172 1193 232
rect 1471 674 1509 685
rect 1315 606 1349 640
rect 1315 538 1349 551
rect 1315 470 1349 479
rect 1315 402 1349 436
rect 1315 334 1349 368
rect 1315 266 1349 300
rect 1315 216 1349 232
rect 1505 651 1509 674
rect 1627 674 1661 708
rect 1783 742 1817 758
rect 1783 685 1817 708
rect 1471 606 1505 640
rect 1471 538 1505 572
rect 1471 470 1505 504
rect 1471 402 1505 436
rect 1471 334 1505 368
rect 1471 266 1505 300
rect 1471 172 1505 232
rect 1745 651 1783 685
rect 1627 606 1661 640
rect 1627 538 1661 551
rect 1627 470 1661 479
rect 1627 402 1661 436
rect 1627 334 1661 368
rect 1627 266 1661 300
rect 1627 216 1661 232
rect 1783 606 1817 640
rect 1783 538 1817 572
rect 1783 470 1817 504
rect 1783 402 1817 436
rect 1783 334 1817 368
rect 1783 266 1817 300
rect 1783 216 1817 232
rect 1939 742 1973 758
rect 1939 674 1973 708
rect 2095 742 2129 758
rect 2095 685 2129 708
rect 2251 742 2285 758
rect 2095 674 2133 685
rect 1939 606 1973 640
rect 1939 538 1973 551
rect 1939 470 1973 479
rect 1939 402 1973 436
rect 1939 334 1973 368
rect 1939 266 1973 300
rect 1939 216 1973 232
rect 2129 651 2133 674
rect 2251 674 2285 708
rect 2095 606 2129 640
rect 2095 538 2129 572
rect 2095 470 2129 504
rect 2095 402 2129 436
rect 2095 334 2129 368
rect 2095 266 2129 300
rect 2095 216 2129 232
rect 2251 606 2285 640
rect 2251 538 2285 551
rect 2251 470 2285 479
rect 2251 402 2285 436
rect 2251 334 2285 368
rect 2251 266 2285 300
rect 2251 216 2285 232
rect 2407 742 2441 758
rect 2407 674 2441 708
rect 2563 742 2597 758
rect 2563 674 2597 708
rect 2407 636 2423 640
rect 2457 636 2495 670
rect 2407 606 2441 636
rect 2407 538 2441 572
rect 2407 470 2441 504
rect 2407 402 2441 436
rect 2407 334 2441 368
rect 2407 266 2441 300
rect 2407 216 2441 232
rect 2563 606 2597 640
rect 2563 538 2597 551
rect 2563 470 2597 479
rect 2563 402 2597 436
rect 2563 334 2597 368
rect 2563 266 2597 300
rect 2563 216 2597 232
rect 2719 742 2753 811
rect 2719 674 2753 708
rect 2719 606 2753 640
rect 2719 538 2753 572
rect 2719 470 2753 504
rect 2719 402 2753 436
rect 2719 334 2753 368
rect 2719 266 2753 300
rect 2719 216 2753 232
rect 2829 742 2863 758
rect 2829 687 2863 708
rect 2985 742 3019 907
rect 3497 857 3537 1012
rect 3297 845 3537 857
rect 3331 811 3369 845
rect 3403 811 3441 845
rect 3475 811 3537 845
rect 2863 653 2901 687
rect 2985 674 3019 708
rect 3141 742 3175 758
rect 3141 687 3175 708
rect 3297 742 3331 811
rect 3571 796 3605 812
rect 2829 606 2863 640
rect 2829 538 2863 572
rect 2829 470 2863 504
rect 2829 402 2863 436
rect 2829 334 2863 368
rect 2829 266 2863 300
rect 2829 216 2863 232
rect 3140 674 3178 687
rect 3140 653 3141 674
rect 2985 606 3019 640
rect 2985 538 3019 572
rect 2985 470 3019 504
rect 2985 402 3019 436
rect 2985 334 3019 368
rect 2985 266 3019 300
rect 2985 172 3019 232
rect 3175 653 3178 674
rect 3297 674 3331 708
rect 3453 742 3487 758
rect 3453 687 3487 708
rect 3141 606 3175 640
rect 3141 538 3175 572
rect 3141 470 3175 504
rect 3141 402 3175 436
rect 3141 334 3175 368
rect 3141 266 3175 300
rect 3141 216 3175 232
rect 3415 653 3453 687
rect 3297 606 3331 640
rect 3297 538 3331 572
rect 3297 470 3331 504
rect 3297 402 3331 436
rect 3297 334 3331 368
rect 3297 266 3331 300
rect 3297 216 3331 232
rect 3453 606 3487 640
rect 3453 538 3487 572
rect 3453 470 3487 504
rect 3453 402 3487 436
rect 3453 334 3487 368
rect 3453 266 3487 300
rect 3453 172 3487 232
rect 328 138 344 172
rect 378 138 390 172
rect 446 138 462 172
rect 514 138 534 172
rect 582 138 606 172
rect 650 138 678 172
rect 718 138 750 172
rect 786 138 820 172
rect 856 138 894 172
rect 1062 138 1078 172
rect 1119 138 1146 172
rect 1191 138 1214 172
rect 1263 138 1282 172
rect 1335 138 1350 172
rect 1407 138 1418 172
rect 1479 138 1486 172
rect 1551 138 1554 172
rect 1588 138 1604 172
rect 2279 123 2295 157
rect 2329 123 2363 157
rect 2397 123 2413 157
rect 2475 138 2491 172
rect 2525 138 2559 172
rect 2605 138 2627 172
rect 2894 138 2910 172
rect 2944 138 2978 172
rect 3012 138 3046 172
rect 3080 138 3096 172
rect 3206 138 3222 172
rect 3256 138 3290 172
rect 3324 138 3358 172
rect 3392 138 3487 172
rect 3571 728 3605 762
rect 3571 660 3605 694
rect 3571 592 3605 626
rect 3571 524 3605 551
rect 3571 456 3605 479
rect 3571 388 3605 422
rect 3571 320 3605 354
rect 3571 252 3605 286
rect 3571 184 3605 218
rect 3571 88 3605 150
rect 151 72 3605 88
rect 151 38 193 72
rect 227 38 261 72
rect 295 38 329 72
rect 363 38 397 72
rect 431 38 465 72
rect 499 38 533 72
rect 567 38 601 72
rect 635 38 669 72
rect 703 38 737 72
rect 771 38 805 72
rect 839 38 873 72
rect 907 38 941 72
rect 975 38 1009 72
rect 1043 38 1077 72
rect 1111 38 1145 72
rect 1179 38 1213 72
rect 1247 38 1281 72
rect 1315 38 1349 72
rect 1383 38 1417 72
rect 1451 38 1485 72
rect 1519 38 1553 72
rect 1587 38 1621 72
rect 1655 38 1689 72
rect 1723 38 1757 72
rect 1791 38 1825 72
rect 1859 38 1893 72
rect 1927 38 1961 72
rect 1995 38 2029 72
rect 2063 38 2097 72
rect 2131 38 2165 72
rect 2199 38 2233 72
rect 2267 38 2301 72
rect 2335 38 2369 72
rect 2403 38 2437 72
rect 2471 38 2505 72
rect 2539 38 2573 72
rect 2607 38 2641 72
rect 2675 38 2709 72
rect 2743 38 2777 72
rect 2811 38 2845 72
rect 2879 38 2913 72
rect 2947 38 2981 72
rect 3015 38 3049 72
rect 3083 38 3117 72
rect 3151 38 3185 72
rect 3219 38 3253 72
rect 3287 38 3321 72
rect 3355 38 3389 72
rect 3423 38 3457 72
rect 3491 38 3525 72
rect 3559 38 3605 72
<< viali >>
rect 115 2247 116 2259
rect 116 2247 149 2259
rect 187 2247 218 2259
rect 218 2247 221 2259
rect 259 2247 286 2259
rect 286 2247 293 2259
rect 115 2225 149 2247
rect 187 2225 221 2247
rect 259 2225 293 2247
rect 305 2247 320 2259
rect 320 2247 354 2259
rect 354 2247 388 2259
rect 388 2247 422 2259
rect 422 2247 437 2259
rect 475 2247 490 2259
rect 490 2247 509 2259
rect 547 2247 558 2259
rect 558 2247 581 2259
rect 619 2247 626 2259
rect 626 2247 653 2259
rect 691 2247 694 2259
rect 694 2247 725 2259
rect 763 2247 796 2259
rect 796 2247 797 2259
rect 835 2247 864 2259
rect 864 2247 869 2259
rect 907 2247 932 2259
rect 932 2247 941 2259
rect 979 2247 1000 2259
rect 1000 2247 1013 2259
rect 1051 2247 1068 2259
rect 1068 2247 1085 2259
rect 1123 2247 1136 2259
rect 1136 2247 1157 2259
rect 1195 2247 1204 2259
rect 1204 2247 1229 2259
rect 1267 2247 1272 2259
rect 1272 2247 1301 2259
rect 1339 2247 1340 2259
rect 1340 2247 1373 2259
rect 1411 2247 1442 2259
rect 1442 2247 1445 2259
rect 1483 2247 1510 2259
rect 1510 2247 1517 2259
rect 1555 2247 1578 2259
rect 1578 2247 1589 2259
rect 1627 2247 1646 2259
rect 1646 2247 1661 2259
rect 1699 2247 1714 2259
rect 1714 2247 1733 2259
rect 1771 2247 1782 2259
rect 1782 2247 1805 2259
rect 1843 2247 1850 2259
rect 1850 2247 1877 2259
rect 1915 2247 1918 2259
rect 1918 2247 1949 2259
rect 1987 2247 2020 2259
rect 2020 2247 2021 2259
rect 2059 2247 2088 2259
rect 2088 2247 2093 2259
rect 2131 2247 2156 2259
rect 2156 2247 2165 2259
rect 2203 2247 2224 2259
rect 2224 2247 2237 2259
rect 2275 2247 2292 2259
rect 2292 2247 2309 2259
rect 2347 2247 2360 2259
rect 2360 2247 2381 2259
rect 2419 2247 2428 2259
rect 2428 2247 2453 2259
rect 2491 2247 2496 2259
rect 2496 2247 2525 2259
rect 2563 2247 2564 2259
rect 2564 2247 2597 2259
rect 2635 2247 2666 2259
rect 2666 2247 2669 2259
rect 2707 2247 2734 2259
rect 2734 2247 2741 2259
rect 2779 2247 2802 2259
rect 2802 2247 2813 2259
rect 2851 2247 2870 2259
rect 2870 2247 2885 2259
rect 2923 2247 2938 2259
rect 2938 2247 2957 2259
rect 2995 2247 3006 2259
rect 3006 2247 3029 2259
rect 3067 2247 3074 2259
rect 3074 2247 3101 2259
rect 305 2225 437 2247
rect 475 2225 509 2247
rect 547 2225 581 2247
rect 619 2225 653 2247
rect 691 2225 725 2247
rect 763 2225 797 2247
rect 835 2225 869 2247
rect 907 2225 941 2247
rect 979 2225 1013 2247
rect 1051 2225 1085 2247
rect 1123 2225 1157 2247
rect 1195 2225 1229 2247
rect 1267 2225 1301 2247
rect 1339 2225 1373 2247
rect 1411 2225 1445 2247
rect 1483 2225 1517 2247
rect 1555 2225 1589 2247
rect 1627 2225 1661 2247
rect 1699 2225 1733 2247
rect 1771 2225 1805 2247
rect 1843 2225 1877 2247
rect 1915 2225 1949 2247
rect 1987 2225 2021 2247
rect 2059 2225 2093 2247
rect 2131 2225 2165 2247
rect 2203 2225 2237 2247
rect 2275 2225 2309 2247
rect 2347 2225 2381 2247
rect 2419 2225 2453 2247
rect 2491 2225 2525 2247
rect 2563 2225 2597 2247
rect 2635 2225 2669 2247
rect 2707 2225 2741 2247
rect 2779 2225 2813 2247
rect 2851 2225 2885 2247
rect 2923 2225 2957 2247
rect 2995 2225 3029 2247
rect 3067 2225 3101 2247
rect 305 2153 411 2225
rect 105 2080 139 2107
rect 105 2073 139 2080
rect 105 2012 139 2035
rect 105 2001 139 2012
rect 261 2046 295 2079
rect 261 2045 295 2046
rect 261 1978 295 2007
rect 261 1973 295 1978
rect 184 1748 218 1749
rect 184 1715 218 1748
rect 256 1715 290 1749
rect 105 1579 139 1595
rect 105 1561 139 1579
rect 105 1511 139 1523
rect 105 1489 139 1511
rect 105 1443 139 1451
rect 105 1417 139 1443
rect 729 2113 763 2147
rect 495 1952 529 1986
rect 495 1880 529 1914
rect 729 2046 763 2075
rect 729 2041 763 2046
rect 589 1910 607 1936
rect 607 1910 623 1936
rect 589 1902 623 1910
rect 661 1902 695 1936
rect 556 1730 590 1764
rect 628 1730 662 1764
rect 438 1579 472 1595
rect 438 1561 472 1579
rect 438 1511 472 1523
rect 438 1489 472 1511
rect 438 1443 472 1451
rect 438 1417 472 1443
rect 870 1511 904 1545
rect 870 1443 904 1473
rect 870 1439 904 1443
rect 654 1347 688 1381
rect 726 1347 760 1381
rect 2444 1939 2478 1973
rect 2516 1939 2550 1973
rect 2204 1785 2238 1819
rect 2276 1785 2310 1819
rect 1641 1641 1675 1675
rect 1713 1641 1747 1675
rect 1785 1641 1819 1675
rect 1857 1641 1891 1675
rect 1929 1641 1963 1675
rect 2001 1641 2035 1675
rect 2073 1641 2107 1675
rect 1302 1511 1336 1545
rect 1302 1443 1336 1473
rect 1302 1439 1336 1443
rect 1734 1579 1768 1595
rect 1734 1561 1768 1579
rect 1734 1511 1768 1523
rect 1734 1489 1768 1511
rect 1734 1443 1768 1451
rect 1734 1417 1768 1443
rect 1098 1337 1132 1371
rect 1170 1337 1204 1371
rect 1484 1337 1518 1371
rect 1556 1337 1590 1371
rect 1878 1337 1912 1371
rect 1950 1337 1984 1371
rect 2094 1579 2200 1595
rect 2094 1545 2166 1579
rect 2166 1545 2200 1579
rect 2094 1511 2200 1545
rect 2094 1477 2166 1511
rect 2166 1477 2200 1511
rect 2094 1443 2200 1477
rect 2094 1417 2166 1443
rect 2166 1417 2200 1443
rect 456 1262 460 1296
rect 460 1262 490 1296
rect 528 1262 562 1296
rect 636 1279 670 1296
rect 708 1279 738 1296
rect 738 1279 742 1296
rect 636 1262 670 1279
rect 708 1262 742 1279
rect 812 1262 846 1296
rect 884 1262 914 1296
rect 914 1262 918 1296
rect 1098 1262 1132 1296
rect 1170 1262 1204 1296
rect 438 1062 472 1069
rect 438 1035 472 1062
rect 438 994 472 997
rect 438 963 472 994
rect 438 891 472 925
rect 902 1164 936 1175
rect 902 1141 936 1164
rect 974 1141 1008 1175
rect 1046 1141 1080 1175
rect 1118 1141 1152 1175
rect 1190 1141 1224 1175
rect 1262 1141 1296 1175
rect 1334 1141 1368 1175
rect 1406 1141 1440 1175
rect 1478 1141 1512 1175
rect 1550 1141 1584 1175
rect 1622 1141 1656 1175
rect 1694 1141 1728 1175
rect 1766 1141 1800 1175
rect 2599 1892 2614 1893
rect 2614 1892 2633 1893
rect 2671 1892 2682 1893
rect 2682 1892 2705 1893
rect 2743 1892 2750 1893
rect 2750 1892 2777 1893
rect 2815 1892 2818 1893
rect 2818 1892 2849 1893
rect 2887 1892 2920 1893
rect 2920 1892 2921 1893
rect 2959 1892 2988 1893
rect 2988 1892 2993 1893
rect 3031 1892 3056 1893
rect 3056 1892 3065 1893
rect 3103 1892 3124 1893
rect 3124 1892 3137 1893
rect 2599 1859 2633 1892
rect 2671 1859 2705 1892
rect 2743 1859 2777 1892
rect 2815 1859 2849 1892
rect 2887 1859 2921 1892
rect 2959 1859 2993 1892
rect 3031 1859 3065 1892
rect 3103 1859 3137 1892
rect 2542 1562 2576 1595
rect 2542 1561 2576 1562
rect 2542 1494 2576 1523
rect 2542 1489 2576 1494
rect 2542 1426 2576 1451
rect 2542 1417 2576 1426
rect 2854 1562 2888 1595
rect 2854 1561 2888 1562
rect 2854 1494 2888 1523
rect 2854 1489 2888 1494
rect 2854 1426 2888 1451
rect 2854 1417 2888 1426
rect 3213 1562 3247 1595
rect 3213 1561 3247 1562
rect 3213 1494 3247 1523
rect 3213 1489 3247 1494
rect 3213 1426 3247 1451
rect 3213 1417 3247 1426
rect 2663 1137 2697 1171
rect 2735 1137 2769 1171
rect 2938 1137 2972 1171
rect 3010 1137 3044 1171
rect 3213 1162 3217 1177
rect 3217 1162 3247 1177
rect 3285 1162 3319 1177
rect 3213 1143 3247 1162
rect 3285 1143 3319 1162
rect 1868 1062 1902 1069
rect 1868 1035 1902 1062
rect 1868 963 1902 997
rect 3525 1562 3559 1595
rect 3525 1561 3559 1562
rect 3525 1494 3559 1523
rect 3525 1489 3559 1494
rect 3525 1426 3559 1451
rect 3525 1417 3559 1426
rect 3453 1162 3487 1177
rect 3525 1162 3555 1177
rect 3555 1162 3559 1177
rect 3453 1143 3487 1162
rect 3525 1143 3559 1162
rect 219 811 253 845
rect 291 811 325 845
rect 363 811 397 845
rect 1067 811 1101 845
rect 1139 811 1173 845
rect 1687 811 1721 845
rect 1759 811 1793 845
rect 1831 811 1865 845
rect 1903 811 1937 845
rect 1975 811 2009 845
rect 2047 811 2081 845
rect 2119 811 2153 845
rect 2191 811 2225 845
rect 2728 811 2762 845
rect 2800 811 2834 845
rect 269 674 303 685
rect 269 651 303 674
rect 341 651 375 685
rect 547 651 581 685
rect 619 651 653 685
rect 821 651 855 685
rect 893 674 927 685
rect 893 651 927 674
rect 1124 651 1158 685
rect 1003 572 1037 585
rect 1003 551 1037 572
rect 1003 504 1037 513
rect 1003 479 1037 504
rect 1196 651 1230 685
rect 1437 651 1471 685
rect 1315 572 1349 585
rect 1315 551 1349 572
rect 1315 504 1349 513
rect 1315 479 1349 504
rect 1509 651 1543 685
rect 1711 651 1745 685
rect 1783 674 1817 685
rect 1783 651 1817 674
rect 1627 572 1661 585
rect 1627 551 1661 572
rect 1627 504 1661 513
rect 1627 479 1661 504
rect 2061 651 2095 685
rect 1939 572 1973 585
rect 1939 551 1973 572
rect 1939 504 1973 513
rect 1939 479 1973 504
rect 2133 651 2167 685
rect 2251 572 2285 585
rect 2251 551 2285 572
rect 2251 504 2285 513
rect 2251 479 2285 504
rect 2423 640 2441 670
rect 2441 640 2457 670
rect 2423 636 2457 640
rect 2495 636 2529 670
rect 2563 572 2597 585
rect 2563 551 2597 572
rect 2563 504 2597 513
rect 2563 479 2597 504
rect 3297 811 3331 845
rect 3369 811 3403 845
rect 3441 811 3475 845
rect 2829 674 2863 687
rect 2829 653 2863 674
rect 2901 653 2935 687
rect 3106 653 3140 687
rect 3178 653 3212 687
rect 3381 653 3415 687
rect 3453 674 3487 687
rect 3453 653 3487 674
rect 390 138 412 172
rect 412 138 424 172
rect 462 138 480 172
rect 480 138 496 172
rect 534 138 548 172
rect 548 138 568 172
rect 606 138 616 172
rect 616 138 640 172
rect 678 138 684 172
rect 684 138 712 172
rect 750 138 752 172
rect 752 138 784 172
rect 822 138 854 172
rect 854 138 856 172
rect 894 138 928 172
rect 1085 138 1112 172
rect 1112 138 1119 172
rect 1157 138 1180 172
rect 1180 138 1191 172
rect 1229 138 1248 172
rect 1248 138 1263 172
rect 1301 138 1316 172
rect 1316 138 1335 172
rect 1373 138 1384 172
rect 1384 138 1407 172
rect 1445 138 1452 172
rect 1452 138 1479 172
rect 1517 138 1520 172
rect 1520 138 1551 172
rect 2571 138 2593 172
rect 2593 138 2605 172
rect 2643 138 2661 172
rect 2661 138 2677 172
rect 3571 558 3605 585
rect 3571 551 3605 558
rect 3571 490 3605 513
rect 3571 479 3605 490
<< metal1 >>
rect 0 2259 3633 2265
rect 0 2225 115 2259
rect 149 2225 187 2259
rect 221 2225 259 2259
rect 293 2225 305 2259
rect 437 2225 475 2259
rect 509 2225 547 2259
rect 581 2225 619 2259
rect 653 2225 691 2259
rect 725 2225 763 2259
rect 797 2225 835 2259
rect 869 2225 907 2259
rect 941 2225 979 2259
rect 1013 2225 1051 2259
rect 1085 2225 1123 2259
rect 1157 2225 1195 2259
rect 1229 2225 1267 2259
rect 1301 2225 1339 2259
rect 1373 2225 1411 2259
rect 1445 2225 1483 2259
rect 1517 2225 1555 2259
rect 1589 2225 1627 2259
rect 1661 2225 1699 2259
rect 1733 2225 1771 2259
rect 1805 2225 1843 2259
rect 1877 2225 1915 2259
rect 1949 2225 1987 2259
rect 2021 2225 2059 2259
rect 2093 2225 2131 2259
rect 2165 2225 2203 2259
rect 2237 2225 2275 2259
rect 2309 2225 2347 2259
rect 2381 2225 2419 2259
rect 2453 2225 2491 2259
rect 2525 2225 2563 2259
rect 2597 2225 2635 2259
rect 2669 2225 2707 2259
rect 2741 2225 2779 2259
rect 2813 2225 2851 2259
rect 2885 2225 2923 2259
rect 2957 2225 2995 2259
rect 3029 2225 3067 2259
rect 3101 2225 3633 2259
rect 0 2153 305 2225
rect 411 2153 3633 2225
rect 0 2147 3633 2153
rect 0 2119 729 2147
tri 74 2094 99 2119 ne
rect 99 2107 145 2119
rect 99 2073 105 2107
rect 139 2073 145 2107
tri 145 2094 170 2119 nw
tri 698 2094 723 2119 ne
rect 723 2113 729 2119
rect 763 2119 3633 2147
rect 763 2113 769 2119
rect 99 2035 145 2073
rect 99 2001 105 2035
rect 139 2001 145 2035
rect 99 1989 145 2001
rect 255 2079 505 2091
rect 255 2045 261 2079
rect 295 2045 505 2079
rect 255 2039 505 2045
rect 557 2039 569 2091
rect 621 2039 627 2091
rect 723 2075 769 2113
tri 769 2094 794 2119 nw
rect 723 2041 729 2075
rect 763 2041 769 2075
rect 255 2007 301 2039
tri 301 2009 331 2039 nw
rect 723 2029 769 2041
rect 829 2039 835 2091
rect 887 2039 899 2091
rect 951 2063 3633 2091
rect 951 2039 957 2063
tri 957 2039 981 2063 nw
rect 255 1973 261 2007
rect 295 1973 301 2007
tri 2365 1998 2402 2035 se
rect 2402 2007 3633 2035
rect 2402 1998 2410 2007
tri 2410 1998 2419 2007 nw
rect 255 1961 301 1973
rect 489 1986 2382 1998
rect 489 1952 495 1986
rect 529 1970 2382 1986
tri 2382 1970 2410 1998 nw
rect 2432 1973 2595 1979
rect 2597 1978 2633 1979
rect 529 1952 535 1970
rect 489 1914 535 1952
tri 535 1940 565 1970 nw
rect 489 1880 495 1914
rect 529 1880 535 1914
rect 577 1936 2239 1942
rect 577 1902 589 1936
rect 623 1902 661 1936
rect 695 1902 2239 1936
rect 577 1899 2239 1902
tri 2239 1899 2282 1942 sw
rect 2432 1939 2444 1973
rect 2478 1939 2516 1973
rect 2550 1939 2595 1973
rect 2432 1927 2595 1939
rect 2596 1928 2634 1978
rect 2597 1927 2633 1928
rect 2635 1927 2658 1979
rect 2710 1927 2722 1979
rect 2774 1927 2780 1979
rect 577 1896 3149 1899
rect 489 1868 535 1880
tri 2219 1853 2262 1896 ne
rect 2262 1893 3149 1896
rect 2262 1859 2599 1893
rect 2633 1859 2671 1893
rect 2705 1859 2743 1893
rect 2777 1859 2815 1893
rect 2849 1859 2887 1893
rect 2921 1859 2959 1893
rect 2993 1859 3031 1893
rect 3065 1859 3103 1893
rect 3137 1859 3149 1893
rect 2262 1853 3149 1859
rect 622 1846 674 1852
tri 597 1770 622 1795 se
rect 622 1782 674 1794
tri 424 1755 439 1770 se
rect 439 1764 622 1770
rect 439 1755 556 1764
rect 172 1749 556 1755
rect 172 1715 184 1749
rect 218 1715 256 1749
rect 290 1730 556 1749
rect 590 1730 622 1764
rect 290 1724 674 1730
rect 702 1800 708 1852
rect 760 1800 772 1852
rect 824 1825 947 1852
tri 947 1825 974 1852 sw
tri 2817 1833 2837 1853 ne
rect 2837 1833 2889 1853
tri 2889 1833 2909 1853 nw
rect 2838 1831 2888 1832
rect 824 1819 2486 1825
rect 824 1800 2204 1819
rect 702 1753 748 1800
tri 748 1775 773 1800 nw
tri 925 1773 952 1800 ne
rect 952 1785 2204 1800
rect 2238 1785 2276 1819
rect 2310 1785 2486 1819
rect 952 1773 2486 1785
tri 2486 1773 2538 1825 sw
rect 2838 1794 2888 1795
tri 2817 1773 2837 1793 se
rect 2837 1773 2889 1793
tri 2889 1773 2909 1793 sw
rect 703 1751 747 1752
rect 290 1715 444 1724
rect 172 1709 444 1715
tri 444 1709 459 1724 nw
rect 702 1715 748 1751
tri 2464 1721 2516 1773 ne
rect 2516 1721 3133 1773
rect 703 1714 747 1715
rect 702 1681 748 1713
tri 748 1681 773 1706 sw
rect 702 1675 3633 1681
rect 702 1641 1641 1675
rect 1675 1641 1713 1675
rect 1747 1641 1785 1675
rect 1819 1641 1857 1675
rect 1891 1641 1929 1675
rect 1963 1641 2001 1675
rect 2035 1641 2073 1675
rect 2107 1641 3633 1675
rect 702 1635 3633 1641
rect 0 1595 3633 1607
rect 0 1561 105 1595
rect 139 1561 438 1595
rect 472 1561 1734 1595
rect 1768 1561 2094 1595
rect 0 1545 2094 1561
rect 0 1523 870 1545
rect 0 1489 105 1523
rect 139 1489 438 1523
rect 472 1511 870 1523
rect 904 1511 1302 1545
rect 1336 1523 2094 1545
rect 1336 1511 1734 1523
rect 472 1489 1734 1511
rect 1768 1489 2094 1523
rect 0 1473 2094 1489
rect 0 1451 870 1473
rect 0 1417 105 1451
rect 139 1417 438 1451
rect 472 1441 870 1451
rect 472 1417 614 1441
rect 0 1405 614 1417
tri 614 1405 650 1441 nw
tri 764 1405 800 1441 ne
rect 800 1439 870 1441
rect 904 1439 1302 1473
rect 1336 1451 2094 1473
rect 1336 1439 1734 1451
rect 800 1417 1734 1439
rect 1768 1417 2094 1451
rect 2200 1561 2542 1595
rect 2576 1561 2854 1595
rect 2888 1561 3213 1595
rect 3247 1561 3525 1595
rect 3559 1561 3633 1595
rect 2200 1523 3633 1561
rect 2200 1489 2542 1523
rect 2576 1489 2854 1523
rect 2888 1489 3213 1523
rect 3247 1489 3525 1523
rect 3559 1489 3633 1523
rect 2200 1451 3633 1489
rect 2200 1417 2542 1451
rect 2576 1417 2854 1451
rect 2888 1417 3213 1451
rect 3247 1417 3525 1451
rect 3559 1417 3633 1451
rect 800 1405 3633 1417
rect 642 1381 772 1387
rect 642 1347 654 1381
rect 688 1347 726 1381
rect 760 1377 772 1381
tri 772 1377 782 1387 sw
rect 760 1371 1408 1377
rect 1410 1376 1446 1377
rect 760 1347 1098 1371
rect 642 1341 1098 1347
tri 752 1331 762 1341 ne
rect 762 1337 1098 1341
rect 1132 1337 1170 1371
rect 1204 1337 1408 1371
rect 762 1331 1408 1337
rect 1409 1332 1447 1376
rect 1448 1371 1996 1377
rect 1448 1337 1484 1371
rect 1518 1337 1556 1371
rect 1590 1337 1878 1371
rect 1912 1337 1950 1371
rect 1984 1337 1996 1371
rect 1410 1331 1446 1332
rect 1448 1331 1996 1337
rect 444 1296 574 1303
rect 444 1262 456 1296
rect 490 1262 528 1296
rect 562 1262 574 1296
rect 444 1251 574 1262
rect 575 1252 576 1302
rect 612 1252 613 1302
rect 614 1251 632 1303
rect 684 1251 696 1303
rect 748 1251 754 1303
rect 800 1251 810 1303
rect 862 1251 874 1303
rect 926 1251 932 1303
rect 960 1251 966 1303
rect 1018 1251 1030 1303
rect 1082 1296 2483 1303
rect 1082 1262 1098 1296
rect 1132 1262 1170 1296
rect 1204 1262 2483 1296
rect 1082 1251 2483 1262
rect 2535 1251 2547 1303
rect 2599 1251 3633 1303
rect 651 1131 657 1183
rect 709 1131 721 1183
rect 773 1175 2658 1183
rect 773 1141 902 1175
rect 936 1141 974 1175
rect 1008 1141 1046 1175
rect 1080 1141 1118 1175
rect 1152 1141 1190 1175
rect 1224 1141 1262 1175
rect 1296 1141 1334 1175
rect 1368 1141 1406 1175
rect 1440 1141 1478 1175
rect 1512 1141 1550 1175
rect 1584 1141 1622 1175
rect 1656 1141 1694 1175
rect 1728 1141 1766 1175
rect 1800 1141 2658 1175
rect 773 1131 2658 1141
rect 2710 1131 2722 1183
rect 2774 1177 3571 1183
rect 2774 1171 3213 1177
rect 2774 1137 2938 1171
rect 2972 1137 3010 1171
rect 3044 1143 3213 1171
rect 3247 1143 3285 1177
rect 3319 1143 3453 1177
rect 3487 1143 3525 1177
rect 3559 1143 3571 1177
rect 3044 1137 3571 1143
rect 2774 1131 3571 1137
rect 0 1071 3633 1081
rect 0 1069 2713 1071
rect 0 1035 438 1069
rect 472 1035 1868 1069
rect 1902 1035 2713 1069
rect 0 1019 2713 1035
rect 2765 1019 3633 1071
rect 0 1007 3633 1019
rect 0 997 2713 1007
rect 0 963 438 997
rect 472 963 1868 997
rect 1902 963 2713 997
rect 0 955 2713 963
rect 2765 955 3633 1007
rect 0 943 3633 955
rect 0 925 2713 943
rect 0 891 438 925
rect 472 891 2713 925
rect 2765 891 3633 943
rect 0 879 3633 891
rect 207 845 538 851
rect 207 811 219 845
rect 253 811 291 845
rect 325 811 363 845
rect 397 811 538 845
rect 207 799 538 811
tri 538 799 590 851 sw
rect 884 799 890 851
rect 942 799 954 851
rect 1006 799 1013 851
rect 1015 850 1051 851
rect 1014 800 1052 850
rect 1053 845 1189 851
rect 1053 811 1067 845
rect 1101 811 1139 845
rect 1173 811 1189 845
rect 1015 799 1051 800
rect 1053 799 1189 811
rect 1675 845 3487 851
rect 1675 811 1687 845
rect 1721 811 1759 845
rect 1793 811 1831 845
rect 1865 811 1903 845
rect 1937 811 1975 845
rect 2009 811 2047 845
rect 2081 811 2119 845
rect 2153 811 2191 845
rect 2225 811 2728 845
rect 2762 811 2800 845
rect 2834 811 3297 845
rect 3331 811 3369 845
rect 3403 811 3441 845
rect 3475 811 3487 845
rect 1675 805 3487 811
tri 516 771 544 799 ne
rect 544 771 590 799
tri 590 771 618 799 sw
tri 544 719 596 771 ne
rect 596 765 2685 771
rect 596 719 2633 765
tri 2608 694 2633 719 ne
rect 2633 701 2685 713
rect 257 685 1607 691
rect 1609 690 1645 691
rect 257 651 269 685
rect 303 651 341 685
rect 375 651 547 685
rect 581 651 619 685
rect 653 651 821 685
rect 855 651 893 685
rect 927 651 1124 685
rect 1158 651 1196 685
rect 1230 651 1437 685
rect 1471 651 1509 685
rect 1543 651 1607 685
rect 257 645 1607 651
rect 1608 646 1646 690
rect 1647 685 2179 691
rect 1647 651 1711 685
rect 1745 651 1783 685
rect 1817 651 2061 685
rect 2095 651 2133 685
rect 2167 651 2179 685
rect 1609 645 1645 646
rect 1647 645 2179 651
rect 2411 670 2483 682
rect 2411 636 2423 670
rect 2457 636 2483 670
rect 2411 630 2483 636
rect 2535 630 2547 682
rect 2599 630 2605 682
rect 2633 643 2685 649
rect 2817 687 3499 693
rect 2817 653 2829 687
rect 2863 653 2901 687
rect 2935 653 3106 687
rect 3140 653 3178 687
rect 3212 653 3381 687
rect 3415 653 3453 687
rect 3487 653 3499 687
rect 2817 647 3499 653
rect 0 591 3633 597
rect 0 585 2713 591
rect 0 551 1003 585
rect 1037 551 1315 585
rect 1349 551 1627 585
rect 1661 551 1939 585
rect 1973 551 2251 585
rect 2285 551 2563 585
rect 2597 551 2713 585
rect 0 539 2713 551
rect 2765 585 3633 591
rect 2765 551 3571 585
rect 3605 551 3633 585
rect 2765 539 3633 551
rect 0 527 3633 539
rect 0 513 2713 527
rect 0 479 1003 513
rect 1037 479 1315 513
rect 1349 479 1627 513
rect 1661 479 1939 513
rect 1973 479 2251 513
rect 2285 479 2563 513
rect 2597 479 2713 513
rect 0 475 2713 479
rect 2765 513 3633 527
rect 2765 479 3571 513
rect 3605 479 3633 513
rect 2765 475 3633 479
rect 0 467 3633 475
rect 378 172 890 178
rect 378 138 390 172
rect 424 138 462 172
rect 496 138 534 172
rect 568 138 606 172
rect 640 138 678 172
rect 712 138 750 172
rect 784 138 822 172
rect 856 138 890 172
rect 378 126 890 138
rect 942 126 954 178
rect 1006 126 1013 178
rect 1014 127 1015 177
rect 1046 177 1051 178
rect 1046 127 1052 177
rect 1053 172 1604 178
rect 1053 138 1085 172
rect 1119 138 1157 172
rect 1191 138 1229 172
rect 1263 138 1301 172
rect 1335 138 1373 172
rect 1407 138 1445 172
rect 1479 138 1517 172
rect 1551 138 1604 172
rect 1046 126 1051 127
rect 1053 126 1604 138
rect 2559 172 2639 186
rect 2559 138 2571 172
rect 2605 138 2639 172
rect 2559 134 2639 138
rect 2691 134 2703 186
rect 2755 134 2763 186
rect 2559 132 2763 134
<< rmetal1 >>
rect 2595 1978 2597 1979
rect 2633 1978 2635 1979
rect 2595 1928 2596 1978
rect 2634 1928 2635 1978
rect 2595 1927 2597 1928
rect 2633 1927 2635 1928
rect 2837 1832 2889 1833
rect 2837 1831 2838 1832
rect 2888 1831 2889 1832
rect 2837 1794 2838 1795
rect 2888 1794 2889 1795
rect 2837 1793 2889 1794
rect 702 1752 748 1753
rect 702 1751 703 1752
rect 747 1751 748 1752
rect 702 1714 703 1715
rect 747 1714 748 1715
rect 702 1713 748 1714
rect 1408 1376 1410 1377
rect 1446 1376 1448 1377
rect 1408 1332 1409 1376
rect 1447 1332 1448 1376
rect 1408 1331 1410 1332
rect 1446 1331 1448 1332
rect 574 1302 576 1303
rect 574 1252 575 1302
rect 574 1251 576 1252
rect 612 1302 614 1303
rect 613 1252 614 1302
rect 612 1251 614 1252
rect 1013 850 1015 851
rect 1051 850 1053 851
rect 1013 800 1014 850
rect 1052 800 1053 850
rect 1013 799 1015 800
rect 1051 799 1053 800
rect 1607 690 1609 691
rect 1645 690 1647 691
rect 1607 646 1608 690
rect 1646 646 1647 690
rect 1607 645 1609 646
rect 1645 645 1647 646
rect 1013 177 1015 178
rect 1013 127 1014 177
rect 1013 126 1015 127
rect 1051 177 1053 178
rect 1052 127 1053 177
rect 1051 126 1053 127
<< via1 >>
rect 505 2039 557 2091
rect 569 2039 621 2091
rect 835 2039 887 2091
rect 899 2039 951 2091
rect 2658 1927 2710 1979
rect 2722 1927 2774 1979
rect 622 1794 674 1846
rect 622 1764 674 1782
rect 622 1730 628 1764
rect 628 1730 662 1764
rect 662 1730 674 1764
rect 708 1800 760 1852
rect 772 1800 824 1852
rect 632 1296 684 1303
rect 632 1262 636 1296
rect 636 1262 670 1296
rect 670 1262 684 1296
rect 632 1251 684 1262
rect 696 1296 748 1303
rect 696 1262 708 1296
rect 708 1262 742 1296
rect 742 1262 748 1296
rect 696 1251 748 1262
rect 810 1296 862 1303
rect 810 1262 812 1296
rect 812 1262 846 1296
rect 846 1262 862 1296
rect 810 1251 862 1262
rect 874 1296 926 1303
rect 874 1262 884 1296
rect 884 1262 918 1296
rect 918 1262 926 1296
rect 874 1251 926 1262
rect 966 1251 1018 1303
rect 1030 1251 1082 1303
rect 2483 1251 2535 1303
rect 2547 1251 2599 1303
rect 657 1131 709 1183
rect 721 1131 773 1183
rect 2658 1171 2710 1183
rect 2658 1137 2663 1171
rect 2663 1137 2697 1171
rect 2697 1137 2710 1171
rect 2658 1131 2710 1137
rect 2722 1171 2774 1183
rect 2722 1137 2735 1171
rect 2735 1137 2769 1171
rect 2769 1137 2774 1171
rect 2722 1131 2774 1137
rect 2713 1019 2765 1071
rect 2713 955 2765 1007
rect 2713 891 2765 943
rect 890 799 942 851
rect 954 799 1006 851
rect 2633 713 2685 765
rect 2483 670 2535 682
rect 2483 636 2495 670
rect 2495 636 2529 670
rect 2529 636 2535 670
rect 2483 630 2535 636
rect 2547 630 2599 682
rect 2633 649 2685 701
rect 2713 539 2765 591
rect 2713 475 2765 527
rect 890 172 942 178
rect 890 138 894 172
rect 894 138 928 172
rect 928 138 942 172
rect 890 126 942 138
rect 954 126 1006 178
rect 2639 172 2691 186
rect 2639 138 2643 172
rect 2643 138 2677 172
rect 2677 138 2691 172
rect 2639 134 2691 138
rect 2703 134 2755 186
<< metal2 >>
rect 499 2039 505 2091
rect 557 2039 569 2091
rect 621 2039 627 2091
rect 829 2039 835 2091
rect 887 2039 899 2091
rect 951 2039 957 2091
rect 499 1251 563 2039
tri 563 2014 588 2039 nw
tri 855 2014 880 2039 ne
tri 855 1941 880 1966 se
rect 880 1941 932 2039
tri 932 2014 957 2039 nw
rect 622 1889 932 1941
rect 622 1846 674 1889
tri 674 1864 699 1889 nw
tri 855 1864 880 1889 ne
rect 622 1782 674 1794
rect 622 1724 674 1730
rect 702 1800 708 1852
rect 760 1800 772 1852
rect 824 1800 830 1852
tri 677 1303 702 1328 se
rect 702 1303 754 1800
tri 754 1775 779 1800 nw
tri 855 1303 880 1328 se
rect 880 1303 932 1889
rect 2652 1927 2658 1979
rect 2710 1927 2722 1979
rect 2774 1927 2780 1979
tri 563 1251 584 1272 sw
rect 626 1251 632 1303
rect 684 1251 696 1303
rect 748 1251 754 1303
rect 804 1251 810 1303
rect 862 1251 874 1303
rect 926 1251 932 1303
rect 960 1251 966 1303
rect 1018 1251 1030 1303
rect 1082 1251 1088 1303
rect 2477 1251 2483 1303
rect 2535 1251 2547 1303
rect 2599 1251 2605 1303
rect 499 1246 584 1251
tri 499 1182 563 1246 ne
rect 563 1183 584 1246
tri 584 1183 652 1251 sw
rect 563 1182 657 1183
tri 563 1131 614 1182 ne
rect 614 1131 657 1182
rect 709 1131 721 1183
rect 773 1131 779 1183
tri 935 851 960 876 se
rect 960 851 1012 1251
tri 1012 1226 1037 1251 nw
tri 2528 1226 2553 1251 ne
rect 884 799 890 851
rect 942 799 954 851
rect 1006 799 1012 851
tri 935 774 960 799 ne
tri 935 178 960 203 se
rect 960 178 1012 799
tri 2528 682 2553 707 se
rect 2553 682 2605 1251
rect 2652 1183 2704 1927
tri 2704 1902 2729 1927 nw
tri 2704 1183 2729 1208 sw
rect 2652 1131 2658 1183
rect 2710 1131 2722 1183
rect 2774 1131 2780 1183
rect 2713 1071 2765 1081
rect 2713 1007 2765 1019
rect 2713 943 2765 955
rect 2477 630 2483 682
rect 2535 630 2547 682
rect 2599 630 2605 682
rect 2633 765 2685 771
rect 2633 701 2685 713
rect 884 126 890 178
rect 942 126 954 178
rect 1006 126 1012 178
rect 2633 186 2685 649
rect 2713 591 2765 891
rect 2713 527 2765 539
rect 2713 469 2765 475
tri 2685 186 2710 211 sw
rect 2633 134 2639 186
rect 2691 134 2703 186
rect 2755 134 2761 186
use sky130_fd_io__tk_em1o_cdns_5595914180880  sky130_fd_io__tk_em1o_cdns_5595914180880_0
timestamp 1676037725
transform 1 0 522 0 1 1251
box 0 0 1 1
use sky130_fd_io__tk_em1o_cdns_5595914180880  sky130_fd_io__tk_em1o_cdns_5595914180880_1
timestamp 1676037725
transform -1 0 1105 0 1 126
box 0 0 1 1
use sky130_fd_io__tk_em1o_cdns_55959141808302  sky130_fd_io__tk_em1o_cdns_55959141808302_0
timestamp 1676037725
transform 0 -1 2889 1 0 1741
box 0 0 1 1
use sky130_fd_io__tk_em1s_cdns_5595914180881  sky130_fd_io__tk_em1s_cdns_5595914180881_0
timestamp 1676037725
transform 1 0 1555 0 1 645
box 0 0 1 1
use sky130_fd_io__tk_em1s_cdns_5595914180881  sky130_fd_io__tk_em1s_cdns_5595914180881_1
timestamp 1676037725
transform 1 0 1356 0 1 1331
box 0 0 1 1
use sky130_fd_io__tk_em1s_cdns_5595914180882  sky130_fd_io__tk_em1s_cdns_5595914180882_0
timestamp 1676037725
transform -1 0 1105 0 1 799
box 0 0 1 1
use sky130_fd_io__tk_em1s_cdns_5595914180882  sky130_fd_io__tk_em1s_cdns_5595914180882_1
timestamp 1676037725
transform -1 0 2687 0 1 1927
box 0 0 1 1
use sky130_fd_io__tk_em1s_cdns_55959141808301  sky130_fd_io__tk_em1s_cdns_55959141808301_0
timestamp 1676037725
transform 0 -1 748 -1 0 1805
box 0 0 1 1
use sky130_fd_pr__nfet_01v8__example_55959141808281  sky130_fd_pr__nfet_01v8__example_55959141808281_0
timestamp 1676037725
transform -1 0 1857 0 -1 1074
box -1 0 801 1
use sky130_fd_pr__nfet_01v8__example_55959141808282  sky130_fd_pr__nfet_01v8__example_55959141808282_0
timestamp 1676037725
transform 1 0 483 0 1 914
box -1 0 0 1
use sky130_fd_pr__nfet_01v8__example_55959141808303  sky130_fd_pr__nfet_01v8__example_55959141808303_0
timestamp 1676037725
transform 1 0 1913 0 -1 1074
box -1 0 1601 1
use sky130_fd_pr__nfet_01v8__example_55959141808304  sky130_fd_pr__nfet_01v8__example_55959141808304_0
timestamp 1676037725
transform 1 0 2452 0 1 220
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808304  sky130_fd_pr__nfet_01v8__example_55959141808304_1
timestamp 1676037725
transform -1 0 2396 0 1 220
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808304  sky130_fd_pr__nfet_01v8__example_55959141808304_2
timestamp 1676037725
transform 1 0 2608 0 1 220
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808305  sky130_fd_pr__nfet_01v8__example_55959141808305_0
timestamp 1676037725
transform -1 0 3442 0 1 220
box -1 0 257 1
use sky130_fd_pr__nfet_01v8__example_55959141808307  sky130_fd_pr__nfet_01v8__example_55959141808307_0
timestamp 1676037725
transform -1 0 882 0 1 220
box -1 0 569 1
use sky130_fd_pr__nfet_01v8__example_55959141808307  sky130_fd_pr__nfet_01v8__example_55959141808307_1
timestamp 1676037725
transform -1 0 2240 0 1 220
box -1 0 569 1
use sky130_fd_pr__nfet_01v8__example_55959141808307  sky130_fd_pr__nfet_01v8__example_55959141808307_2
timestamp 1676037725
transform -1 0 1616 0 1 220
box -1 0 569 1
use sky130_fd_pr__nfet_01v8__example_55959141808308  sky130_fd_pr__nfet_01v8__example_55959141808308_0
timestamp 1676037725
transform 1 0 637 0 1 914
box 0 0 1 1
use sky130_fd_pr__nfet_01v8__example_55959141808309  sky130_fd_pr__nfet_01v8__example_55959141808309_0
timestamp 1676037725
transform 1 0 791 0 1 914
box 100 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808310  sky130_fd_pr__nfet_01v8__example_55959141808310_0
timestamp 1676037725
transform 1 0 2874 0 1 220
box -1 0 257 1
use sky130_fd_pr__nfet_01v8__example_55959141808311  sky130_fd_pr__nfet_01v8__example_55959141808311_0
timestamp 1676037725
transform -1 0 380 0 1 1014
box 120 0 121 1
use sky130_fd_pr__pfet_01v8__example_55959141808312  sky130_fd_pr__pfet_01v8__example_55959141808312_0
timestamp 1676037725
transform 1 0 3258 0 1 1244
box -1 0 257 1
use sky130_fd_pr__pfet_01v8__example_55959141808313  sky130_fd_pr__pfet_01v8__example_55959141808313_0
timestamp 1676037725
transform 1 0 462 0 1 1898
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808313  sky130_fd_pr__pfet_01v8__example_55959141808313_1
timestamp 1676037725
transform -1 0 718 0 1 1898
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808313  sky130_fd_pr__pfet_01v8__example_55959141808313_2
timestamp 1676037725
transform 1 0 150 0 1 1898
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808313  sky130_fd_pr__pfet_01v8__example_55959141808313_3
timestamp 1676037725
transform -1 0 406 0 1 1898
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808314  sky130_fd_pr__pfet_01v8__example_55959141808314_0
timestamp 1676037725
transform -1 0 2421 0 1 1244
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808315  sky130_fd_pr__pfet_01v8__example_55959141808315_0
timestamp 1676037725
transform 1 0 1347 0 1 1397
box -1 0 809 1
use sky130_fd_pr__pfet_01v8__example_55959141808315  sky130_fd_pr__pfet_01v8__example_55959141808315_1
timestamp 1676037725
transform 1 0 483 0 1 1397
box -1 0 809 1
use sky130_fd_pr__pfet_01v8__example_55959141808317  sky130_fd_pr__pfet_01v8__example_55959141808317_0
timestamp 1676037725
transform 1 0 2587 0 1 1244
box -1 0 413 1
use sky130_fd_pr__pfet_01v8__example_55959141808318  sky130_fd_pr__pfet_01v8__example_55959141808318_0
timestamp 1676037725
transform 1 0 150 0 1 1397
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808319  sky130_fd_pr__pfet_01v8__example_55959141808319_0
timestamp 1676037725
transform 1 0 821 0 1 2014
box 1600 0 1601 1
use sky130_fd_pr__tpl1__example_55959141808299  sky130_fd_pr__tpl1__example_55959141808299_0
timestamp 1676037725
transform 0 1 867 -1 0 1888
box 0 0 1 1
use sky130_fd_pr__tpl1__example_55959141808300  sky130_fd_pr__tpl1__example_55959141808300_0
timestamp 1676037725
transform 0 1 2608 -1 0 2182
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_0
timestamp 1676037725
transform 0 1 3571 1 0 479
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_1
timestamp 1676037725
transform 0 -1 529 -1 0 1986
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_2
timestamp 1676037725
transform 1 0 556 0 1 1730
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_3
timestamp 1676037725
transform 1 0 184 0 1 1715
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_4
timestamp 1676037725
transform 1 0 2571 0 1 138
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_5
timestamp 1676037725
transform 1 0 654 0 -1 1381
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_6
timestamp 1676037725
transform 1 0 2728 0 -1 845
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_7
timestamp 1676037725
transform 1 0 547 0 -1 685
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_8
timestamp 1676037725
transform -1 0 2529 0 -1 670
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_9
timestamp 1676037725
transform 1 0 1098 0 -1 1296
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_10
timestamp 1676037725
transform -1 0 1590 0 1 1337
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_11
timestamp 1676037725
transform 1 0 1098 0 -1 1371
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_12
timestamp 1676037725
transform 0 -1 295 1 0 1973
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_13
timestamp 1676037725
transform 1 0 3106 0 -1 687
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_14
timestamp 1676037725
transform -1 0 2769 0 1 1137
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_15
timestamp 1676037725
transform -1 0 3044 0 1 1137
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_16
timestamp 1676037725
transform 1 0 3453 0 -1 1177
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_17
timestamp 1676037725
transform -1 0 2550 0 -1 1973
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_18
timestamp 1676037725
transform 1 0 589 0 1 1902
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_19
timestamp 1676037725
transform -1 0 2310 0 1 1785
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_20
timestamp 1676037725
transform 1 0 636 0 1 1262
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_21
timestamp 1676037725
transform -1 0 562 0 1 1262
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_22
timestamp 1676037725
transform 0 -1 1902 -1 0 1069
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_23
timestamp 1676037725
transform 0 -1 1336 1 0 1439
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_24
timestamp 1676037725
transform 1 0 812 0 1 1262
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_25
timestamp 1676037725
transform 1 0 821 0 -1 685
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_26
timestamp 1676037725
transform 1 0 269 0 -1 685
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_27
timestamp 1676037725
transform 0 1 1003 1 0 479
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_28
timestamp 1676037725
transform 0 1 2251 1 0 479
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_29
timestamp 1676037725
transform 0 1 1627 1 0 479
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_30
timestamp 1676037725
transform 0 1 1939 1 0 479
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_31
timestamp 1676037725
transform 0 1 1315 1 0 479
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_32
timestamp 1676037725
transform 0 1 2563 1 0 479
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_33
timestamp 1676037725
transform 1 0 3381 0 -1 687
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_34
timestamp 1676037725
transform 1 0 2829 0 -1 687
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_35
timestamp 1676037725
transform 1 0 1711 0 -1 685
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_36
timestamp 1676037725
transform 0 -1 904 1 0 1439
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_37
timestamp 1676037725
transform 1 0 3213 0 -1 1177
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_38
timestamp 1676037725
transform 1 0 1067 0 -1 845
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_39
timestamp 1676037725
transform 0 1 105 -1 0 2107
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_40
timestamp 1676037725
transform 0 1 729 -1 0 2147
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_41
timestamp 1676037725
transform 1 0 1437 0 -1 685
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_42
timestamp 1676037725
transform 1 0 1124 0 -1 685
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_43
timestamp 1676037725
transform -1 0 1984 0 1 1337
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_44
timestamp 1676037725
transform 1 0 2061 0 -1 685
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_45
timestamp 1676037725
transform 1 0 305 0 1 2153
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180857  sky130_fd_pr__via_l1m1__example_5595914180857_0
timestamp 1676037725
transform 0 1 2094 -1 0 1595
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_0
timestamp 1676037725
transform -1 0 397 0 1 811
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_1
timestamp 1676037725
transform -1 0 3475 0 -1 845
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_2
timestamp 1676037725
transform 0 -1 3559 -1 0 1595
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_3
timestamp 1676037725
transform 0 -1 3247 -1 0 1595
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_4
timestamp 1676037725
transform 0 -1 2888 -1 0 1595
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_5
timestamp 1676037725
transform 0 -1 2576 -1 0 1595
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_6
timestamp 1676037725
transform 0 -1 472 -1 0 1069
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_7
timestamp 1676037725
transform 0 -1 472 1 0 1417
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_8
timestamp 1676037725
transform 0 -1 139 1 0 1417
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_9
timestamp 1676037725
transform 0 -1 1768 -1 0 1595
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808290  sky130_fd_pr__via_l1m1__example_55959141808290_0
timestamp 1676037725
transform 1 0 1687 0 -1 845
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808290  sky130_fd_pr__via_l1m1__example_55959141808290_1
timestamp 1676037725
transform -1 0 928 0 -1 172
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808290  sky130_fd_pr__via_l1m1__example_55959141808290_2
timestamp 1676037725
transform -1 0 3137 0 1 1859
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808291  sky130_fd_pr__via_l1m1__example_55959141808291_0
timestamp 1676037725
transform 1 0 1085 0 -1 172
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808291  sky130_fd_pr__via_l1m1__example_55959141808291_1
timestamp 1676037725
transform -1 0 2107 0 1 1641
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808292  sky130_fd_pr__via_l1m1__example_55959141808292_0
timestamp 1676037725
transform -1 0 1800 0 -1 1175
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808293  sky130_fd_pr__via_l1m1__example_55959141808293_0
timestamp 1676037725
transform -1 0 3101 0 1 2225
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_0
timestamp 1676037725
transform -1 0 957 0 1 2039
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_1
timestamp 1676037725
transform 0 -1 2685 -1 0 771
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_2
timestamp 1676037725
transform 1 0 2633 0 -1 186
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_3
timestamp 1676037725
transform 0 -1 2765 1 0 469
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_4
timestamp 1676037725
transform 1 0 2652 0 1 1131
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_5
timestamp 1676037725
transform 1 0 2477 0 1 1251
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_6
timestamp 1676037725
transform -1 0 1012 0 1 799
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_7
timestamp 1676037725
transform 1 0 884 0 -1 178
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_8
timestamp 1676037725
transform -1 0 1088 0 1 1251
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_9
timestamp 1676037725
transform 1 0 499 0 -1 2091
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_10
timestamp 1676037725
transform 1 0 651 0 1 1131
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_11
timestamp 1676037725
transform -1 0 2780 0 1 1927
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_12
timestamp 1676037725
transform 1 0 702 0 -1 1852
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_13
timestamp 1676037725
transform -1 0 754 0 1 1251
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_14
timestamp 1676037725
transform 1 0 804 0 -1 1303
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_15
timestamp 1676037725
transform 0 1 622 1 0 1724
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_16
timestamp 1676037725
transform -1 0 2605 0 1 630
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808261  sky130_fd_pr__via_m1m2__example_55959141808261_0
timestamp 1676037725
transform 0 -1 2765 -1 0 1077
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_0
timestamp 1676037725
transform 1 0 2280 0 1 1876
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_0
timestamp 1676037725
transform 0 -1 1601 1 0 1629
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_1
timestamp 1676037725
transform 0 1 3201 1 0 1146
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_2
timestamp 1676037725
transform 0 1 445 1 0 2141
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_3
timestamp 1676037725
transform 1 0 324 0 1 1732
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_4
timestamp 1676037725
transform 0 1 600 -1 0 1847
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_5
timestamp 1676037725
transform 0 1 620 -1 0 1329
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_6
timestamp 1676037725
transform 0 1 2279 1 0 107
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_7
timestamp 1676037725
transform 0 1 3437 1 0 1146
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_8
timestamp 1676037725
transform 0 -1 578 -1 0 1312
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_9
timestamp 1676037725
transform 0 1 796 -1 0 1312
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808274  sky130_fd_pr__via_pol1__example_55959141808274_0
timestamp 1676037725
transform 0 1 3206 1 0 122
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808274  sky130_fd_pr__via_pol1__example_55959141808274_1
timestamp 1676037725
transform 0 1 2894 1 0 122
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808274  sky130_fd_pr__via_pol1__example_55959141808274_2
timestamp 1676037725
transform 0 -1 2677 1 0 122
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808274  sky130_fd_pr__via_pol1__example_55959141808274_3
timestamp 1676037725
transform 1 0 168 0 -1 1866
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808294  sky130_fd_pr__via_pol1__example_55959141808294_0
timestamp 1676037725
transform 0 1 328 -1 0 188
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808294  sky130_fd_pr__via_pol1__example_55959141808294_1
timestamp 1676037725
transform 0 1 1062 -1 0 188
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808294  sky130_fd_pr__via_pol1__example_55959141808294_2
timestamp 1676037725
transform 0 1 1686 -1 0 918
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808294  sky130_fd_pr__via_pol1__example_55959141808294_3
timestamp 1676037725
transform 0 1 2598 1 0 1876
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808294  sky130_fd_pr__via_pol1__example_55959141808294_4
timestamp 1676037725
transform 0 -1 1820 1 0 1253
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808295  sky130_fd_pr__via_pol1__example_55959141808295_0
timestamp 1676037725
transform 0 1 1966 -1 0 1172
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808296  sky130_fd_pr__via_pol1__example_55959141808296_0
timestamp 1676037725
transform 0 1 825 1 0 1916
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808297  sky130_fd_pr__via_pol1__example_55959141808297_0
timestamp 1676037725
transform 0 -1 1820 1 0 1106
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808298  sky130_fd_pr__via_pol1__example_55959141808298_0
timestamp 1676037725
transform 0 -1 1236 1 0 1629
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808298  sky130_fd_pr__via_pol1__example_55959141808298_1
timestamp 1676037725
transform 0 1 511 1 0 1629
box 0 0 1 1
<< labels >>
flabel locali s 2363 123 2413 157 0 FreeSans 300 0 0 0 EN_H_N
port 2 nsew
flabel locali s 340 1795 374 1866 8 FreeSans 300 0 0 0 EN_H
port 1 nsew
flabel metal1 s 3591 467 3633 597 7 FreeSans 300 180 0 0 VGND_IO
port 3 nsew
flabel metal1 s 3593 1251 3633 1303 7 FreeSans 300 180 0 0 NBIAS
port 5 nsew
flabel metal1 s 3593 2063 3633 2091 7 FreeSans 300 180 0 0 DRVHI_H
port 4 nsew
flabel metal1 s 3593 2007 3633 2035 7 FreeSans 300 180 0 0 PUEN_H
port 6 nsew
flabel metal1 s 3591 879 3633 1081 7 FreeSans 300 180 0 0 VGND_IO
port 3 nsew
flabel metal1 s 3593 1405 3633 1607 7 FreeSans 300 180 0 0 VCC_IO
port 7 nsew
flabel metal1 s 3593 1635 3633 1681 7 FreeSans 300 180 0 0 PU_H_N
port 8 nsew
flabel metal1 s 0 467 42 597 7 FreeSans 300 0 0 0 VGND_IO
port 3 nsew
flabel metal1 s 0 879 42 1081 7 FreeSans 300 0 0 0 VGND_IO
port 3 nsew
flabel metal1 s 0 1405 42 1607 6 FreeSans 300 0 0 0 VCC_IO
port 7 nsew
flabel metal1 s 702 1635 744 1681 7 FreeSans 300 180 0 0 PU_H_N
port 8 nsew
flabel metal1 s 0 2119 37 2265 6 FreeSans 300 0 0 0 VCC_IO
port 7 nsew
flabel metal1 s 3593 2119 3633 2265 7 FreeSans 300 180 0 0 VCC_IO
port 7 nsew
flabel comment s 1970 676 1970 676 0 FreeSans 300 0 0 0 M1 OPT N<6>
flabel comment s 941 668 941 668 0 FreeSans 300 0 0 0 N<6>
flabel comment s 2579 791 2579 791 0 FreeSans 300 90 0 0 NBIAS
flabel comment s 3136 843 3136 843 0 FreeSans 300 0 0 0 VCCIO_2VTN
flabel comment s 361 1870 361 1870 0 FreeSans 300 180 0 0 EN_H
flabel comment s 888 1310 888 1310 0 FreeSans 300 0 0 0 DRVHI_H
flabel comment s 671 1239 671 1239 0 FreeSans 300 0 0 0 M1 OPT EN_H
flabel comment s 508 1310 508 1310 0 FreeSans 300 0 0 0 EN_H
flabel comment s 2891 1884 2891 1884 0 FreeSans 300 0 0 0 N<1>
flabel comment s 2353 1940 2353 1940 0 FreeSans 300 0 0 0 N<2>
flabel comment s 3336 1210 3336 1210 0 FreeSans 300 0 0 0 BIAS_G
flabel comment s 1283 1629 1283 1629 0 FreeSans 300 0 0 0 BIAS_G
flabel comment s 2879 1108 2879 1108 0 FreeSans 300 0 0 0 VCCIO
flabel comment s 1423 1201 1423 1201 0 FreeSans 300 0 0 0 BIAS_G
flabel comment s 1881 1032 1881 1032 0 FreeSans 300 270 0 0 VGND_IO
flabel comment s 3082 677 3082 677 0 FreeSans 300 0 0 0 N<8>
flabel comment s 1883 525 1883 525 0 FreeSans 300 0 0 0 VGND_IO
flabel comment s 2755 737 2755 737 0 FreeSans 300 90 0 0 VCCIO_2VTN
flabel comment s 1891 857 1891 857 0 FreeSans 300 0 0 0 VCCIO_2VTN
flabel comment s 2587 192 2587 192 0 FreeSans 300 0 0 0 DRVHI_H_N
flabel comment s 2341 192 2341 192 0 FreeSans 300 0 0 0 EN_H_N
flabel comment s 1267 190 1267 190 0 FreeSans 300 0 0 0 N<6>
flabel comment s 533 190 533 190 0 FreeSans 300 0 0 0 NBIAS
flabel comment s 1967 1990 1967 1990 0 FreeSans 300 180 0 0 PU_H_N
flabel comment s 2238 1522 2238 1522 0 FreeSans 300 0 0 0 VCCIO
flabel comment s 429 2046 429 2046 0 FreeSans 300 0 0 0 VCCIO
flabel comment s 203 1352 203 1352 0 FreeSans 300 0 0 0 DRVHI_H_N
flabel comment s 611 1709 611 1709 0 FreeSans 300 90 0 0 N<2>
flabel comment s 2853 920 2853 920 0 FreeSans 300 0 0 0 VGND_IO
flabel comment s 1305 1800 1305 1800 0 FreeSans 300 180 0 0 N<2>
flabel comment s 1307 1934 1307 1934 0 FreeSans 300 0 0 0 N<1>
flabel comment s 620 1151 620 1151 0 FreeSans 300 270 0 0 N<4>
flabel comment s 776 1151 776 1151 0 FreeSans 300 270 0 0 N<3>
flabel comment s 887 1361 887 1361 0 FreeSans 300 0 0 0 NBIAS
flabel comment s 2043 1291 2043 1291 0 FreeSans 300 0 0 0 NBIAS
flabel comment s 2215 1686 2215 1686 0 FreeSans 300 180 0 0 PU_H_N
flabel comment s 3307 179 3307 179 0 FreeSans 300 0 0 0 N<8>
flabel comment s 2992 179 2992 179 0 FreeSans 300 0 0 0 N<7>
<< properties >>
string GDS_END 48824286
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 48791154
<< end >>
