VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wb_buttons_leds
  CLASS BLOCK ;
  FOREIGN wb_buttons_leds ;
  ORIGIN 0.000 0.000 ;
  SIZE 550.000 BY 550.000 ;
  PIN buttons
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.270 0.000 15.550 4.000 ;
    END
  END buttons
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.250 546.000 412.530 550.000 ;
    END
  END clk
  PIN i_wb_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 16.360 4.000 16.960 ;
    END
  END i_wb_addr[0]
  PIN i_wb_addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.760 4.000 71.360 ;
    END
  END i_wb_addr[10]
  PIN i_wb_addr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.200 4.000 76.800 ;
    END
  END i_wb_addr[11]
  PIN i_wb_addr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END i_wb_addr[12]
  PIN i_wb_addr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.080 4.000 87.680 ;
    END
  END i_wb_addr[13]
  PIN i_wb_addr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 92.520 4.000 93.120 ;
    END
  END i_wb_addr[14]
  PIN i_wb_addr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.960 4.000 98.560 ;
    END
  END i_wb_addr[15]
  PIN i_wb_addr[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 103.400 4.000 104.000 ;
    END
  END i_wb_addr[16]
  PIN i_wb_addr[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END i_wb_addr[17]
  PIN i_wb_addr[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 114.280 4.000 114.880 ;
    END
  END i_wb_addr[18]
  PIN i_wb_addr[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.720 4.000 120.320 ;
    END
  END i_wb_addr[19]
  PIN i_wb_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.800 4.000 22.400 ;
    END
  END i_wb_addr[1]
  PIN i_wb_addr[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.160 4.000 125.760 ;
    END
  END i_wb_addr[20]
  PIN i_wb_addr[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 130.600 4.000 131.200 ;
    END
  END i_wb_addr[21]
  PIN i_wb_addr[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 4.000 136.640 ;
    END
  END i_wb_addr[22]
  PIN i_wb_addr[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 141.480 4.000 142.080 ;
    END
  END i_wb_addr[23]
  PIN i_wb_addr[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.920 4.000 147.520 ;
    END
  END i_wb_addr[24]
  PIN i_wb_addr[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 152.360 4.000 152.960 ;
    END
  END i_wb_addr[25]
  PIN i_wb_addr[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 157.800 4.000 158.400 ;
    END
  END i_wb_addr[26]
  PIN i_wb_addr[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 4.000 163.840 ;
    END
  END i_wb_addr[27]
  PIN i_wb_addr[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.680 4.000 169.280 ;
    END
  END i_wb_addr[28]
  PIN i_wb_addr[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.120 4.000 174.720 ;
    END
  END i_wb_addr[29]
  PIN i_wb_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END i_wb_addr[2]
  PIN i_wb_addr[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 179.560 4.000 180.160 ;
    END
  END i_wb_addr[30]
  PIN i_wb_addr[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 185.000 4.000 185.600 ;
    END
  END i_wb_addr[31]
  PIN i_wb_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.680 4.000 33.280 ;
    END
  END i_wb_addr[3]
  PIN i_wb_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.120 4.000 38.720 ;
    END
  END i_wb_addr[4]
  PIN i_wb_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.560 4.000 44.160 ;
    END
  END i_wb_addr[5]
  PIN i_wb_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.000 4.000 49.600 ;
    END
  END i_wb_addr[6]
  PIN i_wb_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END i_wb_addr[7]
  PIN i_wb_addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.880 4.000 60.480 ;
    END
  END i_wb_addr[8]
  PIN i_wb_addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 65.320 4.000 65.920 ;
    END
  END i_wb_addr[9]
  PIN i_wb_cyc
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 55.800 550.000 56.400 ;
    END
  END i_wb_cyc
  PIN i_wb_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 190.440 4.000 191.040 ;
    END
  END i_wb_data[0]
  PIN i_wb_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.840 4.000 245.440 ;
    END
  END i_wb_data[10]
  PIN i_wb_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 250.280 4.000 250.880 ;
    END
  END i_wb_data[11]
  PIN i_wb_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.720 4.000 256.320 ;
    END
  END i_wb_data[12]
  PIN i_wb_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 261.160 4.000 261.760 ;
    END
  END i_wb_data[13]
  PIN i_wb_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 266.600 4.000 267.200 ;
    END
  END i_wb_data[14]
  PIN i_wb_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.040 4.000 272.640 ;
    END
  END i_wb_data[15]
  PIN i_wb_data[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 277.480 4.000 278.080 ;
    END
  END i_wb_data[16]
  PIN i_wb_data[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.920 4.000 283.520 ;
    END
  END i_wb_data[17]
  PIN i_wb_data[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 288.360 4.000 288.960 ;
    END
  END i_wb_data[18]
  PIN i_wb_data[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 293.800 4.000 294.400 ;
    END
  END i_wb_data[19]
  PIN i_wb_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 195.880 4.000 196.480 ;
    END
  END i_wb_data[1]
  PIN i_wb_data[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.240 4.000 299.840 ;
    END
  END i_wb_data[20]
  PIN i_wb_data[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 304.680 4.000 305.280 ;
    END
  END i_wb_data[21]
  PIN i_wb_data[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 310.120 4.000 310.720 ;
    END
  END i_wb_data[22]
  PIN i_wb_data[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 315.560 4.000 316.160 ;
    END
  END i_wb_data[23]
  PIN i_wb_data[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 321.000 4.000 321.600 ;
    END
  END i_wb_data[24]
  PIN i_wb_data[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 326.440 4.000 327.040 ;
    END
  END i_wb_data[25]
  PIN i_wb_data[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 331.880 4.000 332.480 ;
    END
  END i_wb_data[26]
  PIN i_wb_data[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 337.320 4.000 337.920 ;
    END
  END i_wb_data[27]
  PIN i_wb_data[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 342.760 4.000 343.360 ;
    END
  END i_wb_data[28]
  PIN i_wb_data[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 348.200 4.000 348.800 ;
    END
  END i_wb_data[29]
  PIN i_wb_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 201.320 4.000 201.920 ;
    END
  END i_wb_data[2]
  PIN i_wb_data[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 353.640 4.000 354.240 ;
    END
  END i_wb_data[30]
  PIN i_wb_data[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 359.080 4.000 359.680 ;
    END
  END i_wb_data[31]
  PIN i_wb_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 206.760 4.000 207.360 ;
    END
  END i_wb_data[3]
  PIN i_wb_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 212.200 4.000 212.800 ;
    END
  END i_wb_data[4]
  PIN i_wb_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 217.640 4.000 218.240 ;
    END
  END i_wb_data[5]
  PIN i_wb_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 223.080 4.000 223.680 ;
    END
  END i_wb_data[6]
  PIN i_wb_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 228.520 4.000 229.120 ;
    END
  END i_wb_data[7]
  PIN i_wb_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 233.960 4.000 234.560 ;
    END
  END i_wb_data[8]
  PIN i_wb_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 239.400 4.000 240.000 ;
    END
  END i_wb_data[9]
  PIN i_wb_stb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 165.280 550.000 165.880 ;
    END
  END i_wb_stb
  PIN i_wb_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 274.760 550.000 275.360 ;
    END
  END i_wb_we
  PIN led_enb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.890 0.000 37.170 4.000 ;
    END
  END led_enb[0]
  PIN led_enb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.090 0.000 253.370 4.000 ;
    END
  END led_enb[10]
  PIN led_enb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.710 0.000 274.990 4.000 ;
    END
  END led_enb[11]
  PIN led_enb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.510 0.000 58.790 4.000 ;
    END
  END led_enb[1]
  PIN led_enb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.130 0.000 80.410 4.000 ;
    END
  END led_enb[2]
  PIN led_enb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.750 0.000 102.030 4.000 ;
    END
  END led_enb[3]
  PIN led_enb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.370 0.000 123.650 4.000 ;
    END
  END led_enb[4]
  PIN led_enb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 0.000 145.270 4.000 ;
    END
  END led_enb[5]
  PIN led_enb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.610 0.000 166.890 4.000 ;
    END
  END led_enb[6]
  PIN led_enb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.230 0.000 188.510 4.000 ;
    END
  END led_enb[7]
  PIN led_enb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.850 0.000 210.130 4.000 ;
    END
  END led_enb[8]
  PIN led_enb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.470 0.000 231.750 4.000 ;
    END
  END led_enb[9]
  PIN leds[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.330 0.000 296.610 4.000 ;
    END
  END leds[0]
  PIN leds[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.530 0.000 512.810 4.000 ;
    END
  END leds[10]
  PIN leds[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.150 0.000 534.430 4.000 ;
    END
  END leds[11]
  PIN leds[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.950 0.000 318.230 4.000 ;
    END
  END leds[1]
  PIN leds[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.570 0.000 339.850 4.000 ;
    END
  END leds[2]
  PIN leds[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.190 0.000 361.470 4.000 ;
    END
  END leds[3]
  PIN leds[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 382.810 0.000 383.090 4.000 ;
    END
  END leds[4]
  PIN leds[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.430 0.000 404.710 4.000 ;
    END
  END leds[5]
  PIN leds[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.050 0.000 426.330 4.000 ;
    END
  END leds[6]
  PIN leds[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.670 0.000 447.950 4.000 ;
    END
  END leds[7]
  PIN leds[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.290 0.000 469.570 4.000 ;
    END
  END leds[8]
  PIN leds[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 490.910 0.000 491.190 4.000 ;
    END
  END leds[9]
  PIN o_wb_ack
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 384.240 550.000 384.840 ;
    END
  END o_wb_ack
  PIN o_wb_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 364.520 4.000 365.120 ;
    END
  END o_wb_data[0]
  PIN o_wb_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 418.920 4.000 419.520 ;
    END
  END o_wb_data[10]
  PIN o_wb_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 424.360 4.000 424.960 ;
    END
  END o_wb_data[11]
  PIN o_wb_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 429.800 4.000 430.400 ;
    END
  END o_wb_data[12]
  PIN o_wb_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 435.240 4.000 435.840 ;
    END
  END o_wb_data[13]
  PIN o_wb_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 440.680 4.000 441.280 ;
    END
  END o_wb_data[14]
  PIN o_wb_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 446.120 4.000 446.720 ;
    END
  END o_wb_data[15]
  PIN o_wb_data[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 451.560 4.000 452.160 ;
    END
  END o_wb_data[16]
  PIN o_wb_data[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 457.000 4.000 457.600 ;
    END
  END o_wb_data[17]
  PIN o_wb_data[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 462.440 4.000 463.040 ;
    END
  END o_wb_data[18]
  PIN o_wb_data[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 467.880 4.000 468.480 ;
    END
  END o_wb_data[19]
  PIN o_wb_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 369.960 4.000 370.560 ;
    END
  END o_wb_data[1]
  PIN o_wb_data[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 473.320 4.000 473.920 ;
    END
  END o_wb_data[20]
  PIN o_wb_data[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 478.760 4.000 479.360 ;
    END
  END o_wb_data[21]
  PIN o_wb_data[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 484.200 4.000 484.800 ;
    END
  END o_wb_data[22]
  PIN o_wb_data[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 489.640 4.000 490.240 ;
    END
  END o_wb_data[23]
  PIN o_wb_data[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 495.080 4.000 495.680 ;
    END
  END o_wb_data[24]
  PIN o_wb_data[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 500.520 4.000 501.120 ;
    END
  END o_wb_data[25]
  PIN o_wb_data[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 505.960 4.000 506.560 ;
    END
  END o_wb_data[26]
  PIN o_wb_data[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 511.400 4.000 512.000 ;
    END
  END o_wb_data[27]
  PIN o_wb_data[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 516.840 4.000 517.440 ;
    END
  END o_wb_data[28]
  PIN o_wb_data[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 522.280 4.000 522.880 ;
    END
  END o_wb_data[29]
  PIN o_wb_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 375.400 4.000 376.000 ;
    END
  END o_wb_data[2]
  PIN o_wb_data[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 527.720 4.000 528.320 ;
    END
  END o_wb_data[30]
  PIN o_wb_data[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 533.160 4.000 533.760 ;
    END
  END o_wb_data[31]
  PIN o_wb_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 380.840 4.000 381.440 ;
    END
  END o_wb_data[3]
  PIN o_wb_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 386.280 4.000 386.880 ;
    END
  END o_wb_data[4]
  PIN o_wb_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 391.720 4.000 392.320 ;
    END
  END o_wb_data[5]
  PIN o_wb_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 397.160 4.000 397.760 ;
    END
  END o_wb_data[6]
  PIN o_wb_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 402.600 4.000 403.200 ;
    END
  END o_wb_data[7]
  PIN o_wb_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 408.040 4.000 408.640 ;
    END
  END o_wb_data[8]
  PIN o_wb_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 413.480 4.000 414.080 ;
    END
  END o_wb_data[9]
  PIN o_wb_stall
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 493.720 550.000 494.320 ;
    END
  END o_wb_stall
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.170 546.000 137.450 550.000 ;
    END
  END reset
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 538.800 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 538.800 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 544.180 538.645 ;
      LAYER met1 ;
        RECT 0.530 4.460 545.490 538.800 ;
      LAYER met2 ;
        RECT 0.550 545.720 136.890 546.000 ;
        RECT 137.730 545.720 411.970 546.000 ;
        RECT 412.810 545.720 545.470 546.000 ;
        RECT 0.550 4.280 545.470 545.720 ;
        RECT 0.550 4.000 14.990 4.280 ;
        RECT 15.830 4.000 36.610 4.280 ;
        RECT 37.450 4.000 58.230 4.280 ;
        RECT 59.070 4.000 79.850 4.280 ;
        RECT 80.690 4.000 101.470 4.280 ;
        RECT 102.310 4.000 123.090 4.280 ;
        RECT 123.930 4.000 144.710 4.280 ;
        RECT 145.550 4.000 166.330 4.280 ;
        RECT 167.170 4.000 187.950 4.280 ;
        RECT 188.790 4.000 209.570 4.280 ;
        RECT 210.410 4.000 231.190 4.280 ;
        RECT 232.030 4.000 252.810 4.280 ;
        RECT 253.650 4.000 274.430 4.280 ;
        RECT 275.270 4.000 296.050 4.280 ;
        RECT 296.890 4.000 317.670 4.280 ;
        RECT 318.510 4.000 339.290 4.280 ;
        RECT 340.130 4.000 360.910 4.280 ;
        RECT 361.750 4.000 382.530 4.280 ;
        RECT 383.370 4.000 404.150 4.280 ;
        RECT 404.990 4.000 425.770 4.280 ;
        RECT 426.610 4.000 447.390 4.280 ;
        RECT 448.230 4.000 469.010 4.280 ;
        RECT 469.850 4.000 490.630 4.280 ;
        RECT 491.470 4.000 512.250 4.280 ;
        RECT 513.090 4.000 533.870 4.280 ;
        RECT 534.710 4.000 545.470 4.280 ;
      LAYER met3 ;
        RECT 0.525 534.160 546.000 538.725 ;
        RECT 4.400 532.760 546.000 534.160 ;
        RECT 0.525 528.720 546.000 532.760 ;
        RECT 4.400 527.320 546.000 528.720 ;
        RECT 0.525 523.280 546.000 527.320 ;
        RECT 4.400 521.880 546.000 523.280 ;
        RECT 0.525 517.840 546.000 521.880 ;
        RECT 4.400 516.440 546.000 517.840 ;
        RECT 0.525 512.400 546.000 516.440 ;
        RECT 4.400 511.000 546.000 512.400 ;
        RECT 0.525 506.960 546.000 511.000 ;
        RECT 4.400 505.560 546.000 506.960 ;
        RECT 0.525 501.520 546.000 505.560 ;
        RECT 4.400 500.120 546.000 501.520 ;
        RECT 0.525 496.080 546.000 500.120 ;
        RECT 4.400 494.720 546.000 496.080 ;
        RECT 4.400 494.680 545.600 494.720 ;
        RECT 0.525 493.320 545.600 494.680 ;
        RECT 0.525 490.640 546.000 493.320 ;
        RECT 4.400 489.240 546.000 490.640 ;
        RECT 0.525 485.200 546.000 489.240 ;
        RECT 4.400 483.800 546.000 485.200 ;
        RECT 0.525 479.760 546.000 483.800 ;
        RECT 4.400 478.360 546.000 479.760 ;
        RECT 0.525 474.320 546.000 478.360 ;
        RECT 4.400 472.920 546.000 474.320 ;
        RECT 0.525 468.880 546.000 472.920 ;
        RECT 4.400 467.480 546.000 468.880 ;
        RECT 0.525 463.440 546.000 467.480 ;
        RECT 4.400 462.040 546.000 463.440 ;
        RECT 0.525 458.000 546.000 462.040 ;
        RECT 4.400 456.600 546.000 458.000 ;
        RECT 0.525 452.560 546.000 456.600 ;
        RECT 4.400 451.160 546.000 452.560 ;
        RECT 0.525 447.120 546.000 451.160 ;
        RECT 4.400 445.720 546.000 447.120 ;
        RECT 0.525 441.680 546.000 445.720 ;
        RECT 4.400 440.280 546.000 441.680 ;
        RECT 0.525 436.240 546.000 440.280 ;
        RECT 4.400 434.840 546.000 436.240 ;
        RECT 0.525 430.800 546.000 434.840 ;
        RECT 4.400 429.400 546.000 430.800 ;
        RECT 0.525 425.360 546.000 429.400 ;
        RECT 4.400 423.960 546.000 425.360 ;
        RECT 0.525 419.920 546.000 423.960 ;
        RECT 4.400 418.520 546.000 419.920 ;
        RECT 0.525 414.480 546.000 418.520 ;
        RECT 4.400 413.080 546.000 414.480 ;
        RECT 0.525 409.040 546.000 413.080 ;
        RECT 4.400 407.640 546.000 409.040 ;
        RECT 0.525 403.600 546.000 407.640 ;
        RECT 4.400 402.200 546.000 403.600 ;
        RECT 0.525 398.160 546.000 402.200 ;
        RECT 4.400 396.760 546.000 398.160 ;
        RECT 0.525 392.720 546.000 396.760 ;
        RECT 4.400 391.320 546.000 392.720 ;
        RECT 0.525 387.280 546.000 391.320 ;
        RECT 4.400 385.880 546.000 387.280 ;
        RECT 0.525 385.240 546.000 385.880 ;
        RECT 0.525 383.840 545.600 385.240 ;
        RECT 0.525 381.840 546.000 383.840 ;
        RECT 4.400 380.440 546.000 381.840 ;
        RECT 0.525 376.400 546.000 380.440 ;
        RECT 4.400 375.000 546.000 376.400 ;
        RECT 0.525 370.960 546.000 375.000 ;
        RECT 4.400 369.560 546.000 370.960 ;
        RECT 0.525 365.520 546.000 369.560 ;
        RECT 4.400 364.120 546.000 365.520 ;
        RECT 0.525 360.080 546.000 364.120 ;
        RECT 4.400 358.680 546.000 360.080 ;
        RECT 0.525 354.640 546.000 358.680 ;
        RECT 4.400 353.240 546.000 354.640 ;
        RECT 0.525 349.200 546.000 353.240 ;
        RECT 4.400 347.800 546.000 349.200 ;
        RECT 0.525 343.760 546.000 347.800 ;
        RECT 4.400 342.360 546.000 343.760 ;
        RECT 0.525 338.320 546.000 342.360 ;
        RECT 4.400 336.920 546.000 338.320 ;
        RECT 0.525 332.880 546.000 336.920 ;
        RECT 4.400 331.480 546.000 332.880 ;
        RECT 0.525 327.440 546.000 331.480 ;
        RECT 4.400 326.040 546.000 327.440 ;
        RECT 0.525 322.000 546.000 326.040 ;
        RECT 4.400 320.600 546.000 322.000 ;
        RECT 0.525 316.560 546.000 320.600 ;
        RECT 4.400 315.160 546.000 316.560 ;
        RECT 0.525 311.120 546.000 315.160 ;
        RECT 4.400 309.720 546.000 311.120 ;
        RECT 0.525 305.680 546.000 309.720 ;
        RECT 4.400 304.280 546.000 305.680 ;
        RECT 0.525 300.240 546.000 304.280 ;
        RECT 4.400 298.840 546.000 300.240 ;
        RECT 0.525 294.800 546.000 298.840 ;
        RECT 4.400 293.400 546.000 294.800 ;
        RECT 0.525 289.360 546.000 293.400 ;
        RECT 4.400 287.960 546.000 289.360 ;
        RECT 0.525 283.920 546.000 287.960 ;
        RECT 4.400 282.520 546.000 283.920 ;
        RECT 0.525 278.480 546.000 282.520 ;
        RECT 4.400 277.080 546.000 278.480 ;
        RECT 0.525 275.760 546.000 277.080 ;
        RECT 0.525 274.360 545.600 275.760 ;
        RECT 0.525 273.040 546.000 274.360 ;
        RECT 4.400 271.640 546.000 273.040 ;
        RECT 0.525 267.600 546.000 271.640 ;
        RECT 4.400 266.200 546.000 267.600 ;
        RECT 0.525 262.160 546.000 266.200 ;
        RECT 4.400 260.760 546.000 262.160 ;
        RECT 0.525 256.720 546.000 260.760 ;
        RECT 4.400 255.320 546.000 256.720 ;
        RECT 0.525 251.280 546.000 255.320 ;
        RECT 4.400 249.880 546.000 251.280 ;
        RECT 0.525 245.840 546.000 249.880 ;
        RECT 4.400 244.440 546.000 245.840 ;
        RECT 0.525 240.400 546.000 244.440 ;
        RECT 4.400 239.000 546.000 240.400 ;
        RECT 0.525 234.960 546.000 239.000 ;
        RECT 4.400 233.560 546.000 234.960 ;
        RECT 0.525 229.520 546.000 233.560 ;
        RECT 4.400 228.120 546.000 229.520 ;
        RECT 0.525 224.080 546.000 228.120 ;
        RECT 4.400 222.680 546.000 224.080 ;
        RECT 0.525 218.640 546.000 222.680 ;
        RECT 4.400 217.240 546.000 218.640 ;
        RECT 0.525 213.200 546.000 217.240 ;
        RECT 4.400 211.800 546.000 213.200 ;
        RECT 0.525 207.760 546.000 211.800 ;
        RECT 4.400 206.360 546.000 207.760 ;
        RECT 0.525 202.320 546.000 206.360 ;
        RECT 4.400 200.920 546.000 202.320 ;
        RECT 0.525 196.880 546.000 200.920 ;
        RECT 4.400 195.480 546.000 196.880 ;
        RECT 0.525 191.440 546.000 195.480 ;
        RECT 4.400 190.040 546.000 191.440 ;
        RECT 0.525 186.000 546.000 190.040 ;
        RECT 4.400 184.600 546.000 186.000 ;
        RECT 0.525 180.560 546.000 184.600 ;
        RECT 4.400 179.160 546.000 180.560 ;
        RECT 0.525 175.120 546.000 179.160 ;
        RECT 4.400 173.720 546.000 175.120 ;
        RECT 0.525 169.680 546.000 173.720 ;
        RECT 4.400 168.280 546.000 169.680 ;
        RECT 0.525 166.280 546.000 168.280 ;
        RECT 0.525 164.880 545.600 166.280 ;
        RECT 0.525 164.240 546.000 164.880 ;
        RECT 4.400 162.840 546.000 164.240 ;
        RECT 0.525 158.800 546.000 162.840 ;
        RECT 4.400 157.400 546.000 158.800 ;
        RECT 0.525 153.360 546.000 157.400 ;
        RECT 4.400 151.960 546.000 153.360 ;
        RECT 0.525 147.920 546.000 151.960 ;
        RECT 4.400 146.520 546.000 147.920 ;
        RECT 0.525 142.480 546.000 146.520 ;
        RECT 4.400 141.080 546.000 142.480 ;
        RECT 0.525 137.040 546.000 141.080 ;
        RECT 4.400 135.640 546.000 137.040 ;
        RECT 0.525 131.600 546.000 135.640 ;
        RECT 4.400 130.200 546.000 131.600 ;
        RECT 0.525 126.160 546.000 130.200 ;
        RECT 4.400 124.760 546.000 126.160 ;
        RECT 0.525 120.720 546.000 124.760 ;
        RECT 4.400 119.320 546.000 120.720 ;
        RECT 0.525 115.280 546.000 119.320 ;
        RECT 4.400 113.880 546.000 115.280 ;
        RECT 0.525 109.840 546.000 113.880 ;
        RECT 4.400 108.440 546.000 109.840 ;
        RECT 0.525 104.400 546.000 108.440 ;
        RECT 4.400 103.000 546.000 104.400 ;
        RECT 0.525 98.960 546.000 103.000 ;
        RECT 4.400 97.560 546.000 98.960 ;
        RECT 0.525 93.520 546.000 97.560 ;
        RECT 4.400 92.120 546.000 93.520 ;
        RECT 0.525 88.080 546.000 92.120 ;
        RECT 4.400 86.680 546.000 88.080 ;
        RECT 0.525 82.640 546.000 86.680 ;
        RECT 4.400 81.240 546.000 82.640 ;
        RECT 0.525 77.200 546.000 81.240 ;
        RECT 4.400 75.800 546.000 77.200 ;
        RECT 0.525 71.760 546.000 75.800 ;
        RECT 4.400 70.360 546.000 71.760 ;
        RECT 0.525 66.320 546.000 70.360 ;
        RECT 4.400 64.920 546.000 66.320 ;
        RECT 0.525 60.880 546.000 64.920 ;
        RECT 4.400 59.480 546.000 60.880 ;
        RECT 0.525 56.800 546.000 59.480 ;
        RECT 0.525 55.440 545.600 56.800 ;
        RECT 4.400 55.400 545.600 55.440 ;
        RECT 4.400 54.040 546.000 55.400 ;
        RECT 0.525 50.000 546.000 54.040 ;
        RECT 4.400 48.600 546.000 50.000 ;
        RECT 0.525 44.560 546.000 48.600 ;
        RECT 4.400 43.160 546.000 44.560 ;
        RECT 0.525 39.120 546.000 43.160 ;
        RECT 4.400 37.720 546.000 39.120 ;
        RECT 0.525 33.680 546.000 37.720 ;
        RECT 4.400 32.280 546.000 33.680 ;
        RECT 0.525 28.240 546.000 32.280 ;
        RECT 4.400 26.840 546.000 28.240 ;
        RECT 0.525 22.800 546.000 26.840 ;
        RECT 4.400 21.400 546.000 22.800 ;
        RECT 0.525 17.360 546.000 21.400 ;
        RECT 4.400 15.960 546.000 17.360 ;
        RECT 0.525 10.715 546.000 15.960 ;
      LAYER met4 ;
        RECT 8.575 19.895 20.640 531.585 ;
        RECT 23.040 19.895 97.440 531.585 ;
        RECT 99.840 19.895 174.240 531.585 ;
        RECT 176.640 19.895 251.040 531.585 ;
        RECT 253.440 19.895 327.840 531.585 ;
        RECT 330.240 19.895 404.640 531.585 ;
        RECT 407.040 19.895 481.440 531.585 ;
        RECT 483.840 19.895 486.385 531.585 ;
  END
END wb_buttons_leds
END LIBRARY

