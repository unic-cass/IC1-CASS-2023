magic
tech sky130B
magscale 1 2
timestamp 1676037725
<< metal2 >>
rect -4079 12127 -689 12502
rect -4079 11871 -3966 12127
rect -3710 11871 -3442 12127
rect -3186 11871 -2888 12127
rect -2632 11871 -2334 12127
rect -2078 11871 -1810 12127
rect -1554 11871 -689 12127
rect -4079 11633 -689 11871
rect -4079 11377 -3966 11633
rect -3710 11377 -3442 11633
rect -3186 11377 -2888 11633
rect -2632 11377 -2334 11633
rect -2078 11377 -1810 11633
rect -1554 11377 -689 11633
rect -4079 11002 -689 11377
tri -689 11002 811 12502 sw
tri -1311 9000 691 11002 ne
rect 691 10500 811 11002
tri 811 10500 1313 11002 sw
rect 691 10124 4024 10500
rect 691 9868 1511 10124
rect 1767 9868 2035 10124
rect 2291 9868 2589 10124
rect 2845 9868 3143 10124
rect 3399 9868 3667 10124
rect 3923 9868 4024 10124
rect 691 9630 4024 9868
rect 691 9374 1511 9630
rect 1767 9374 2035 9630
rect 2291 9374 2589 9630
rect 2845 9374 3143 9630
rect 3399 9374 3667 9630
rect 3923 9374 4024 9630
rect 691 9000 4024 9374
rect 6408 375 15500 750
rect 6408 119 6552 375
rect 6808 119 7076 375
rect 7332 119 7630 375
rect 7886 119 15500 375
rect 6408 -119 15500 119
rect 6408 -375 6552 -119
rect 6808 -375 7076 -119
rect 7332 -375 7630 -119
rect 7886 -375 15500 -119
rect 6408 -750 15500 -375
tri -1311 -13004 691 -11002 se
rect 691 -11377 3925 -11002
rect 691 -11633 1410 -11377
rect 1666 -11633 1934 -11377
rect 2190 -11633 2488 -11377
rect 2744 -11633 3042 -11377
rect 3298 -11633 3566 -11377
rect 3822 -11633 3925 -11377
rect 691 -11871 3925 -11633
rect 691 -12127 1410 -11871
rect 1666 -12127 1934 -11871
rect 2190 -12127 2488 -11871
rect 2744 -12127 3042 -11871
rect 3298 -12127 3566 -11871
rect 3822 -12127 3925 -11871
rect 691 -12502 3925 -12127
rect 691 -13004 811 -12502
tri 811 -13004 1313 -12502 nw
rect -4123 -13377 -689 -13004
rect -4123 -13633 -4024 -13377
rect -3768 -13633 -3500 -13377
rect -3244 -13633 -2946 -13377
rect -2690 -13633 -2392 -13377
rect -2136 -13633 -1868 -13377
rect -1612 -13633 -689 -13377
rect -4123 -13871 -689 -13633
rect -4123 -14127 -4024 -13871
rect -3768 -14127 -3500 -13871
rect -3244 -14127 -2946 -13871
rect -2690 -14127 -2392 -13871
rect -2136 -14127 -1868 -13871
rect -1612 -14127 -689 -13871
rect -4123 -14504 -689 -14127
tri -689 -14504 811 -13004 nw
<< via2 >>
rect -3966 11871 -3710 12127
rect -3442 11871 -3186 12127
rect -2888 11871 -2632 12127
rect -2334 11871 -2078 12127
rect -1810 11871 -1554 12127
rect -3966 11377 -3710 11633
rect -3442 11377 -3186 11633
rect -2888 11377 -2632 11633
rect -2334 11377 -2078 11633
rect -1810 11377 -1554 11633
rect 1511 9868 1767 10124
rect 2035 9868 2291 10124
rect 2589 9868 2845 10124
rect 3143 9868 3399 10124
rect 3667 9868 3923 10124
rect 1511 9374 1767 9630
rect 2035 9374 2291 9630
rect 2589 9374 2845 9630
rect 3143 9374 3399 9630
rect 3667 9374 3923 9630
rect 6552 119 6808 375
rect 7076 119 7332 375
rect 7630 119 7886 375
rect 6552 -375 6808 -119
rect 7076 -375 7332 -119
rect 7630 -375 7886 -119
rect 1410 -11633 1666 -11377
rect 1934 -11633 2190 -11377
rect 2488 -11633 2744 -11377
rect 3042 -11633 3298 -11377
rect 3566 -11633 3822 -11377
rect 1410 -12127 1666 -11871
rect 1934 -12127 2190 -11871
rect 2488 -12127 2744 -11871
rect 3042 -12127 3298 -11871
rect 3566 -12127 3822 -11871
rect -4024 -13633 -3768 -13377
rect -3500 -13633 -3244 -13377
rect -2946 -13633 -2690 -13377
rect -2392 -13633 -2136 -13377
rect -1868 -13633 -1612 -13377
rect -4024 -14127 -3768 -13871
rect -3500 -14127 -3244 -13871
rect -2946 -14127 -2690 -13871
rect -2392 -14127 -2136 -13871
rect -1868 -14127 -1612 -13871
<< metal3 >>
tri -8131 12382 -6009 14504 se
rect -6009 14497 6009 14504
tri 6009 14497 6016 14504 sw
rect -6009 13004 6016 14497
tri -6009 12382 -5387 13004 nw
tri -5300 12382 -5180 12502 se
rect -5180 12382 -1739 12502
tri -10253 10260 -8131 12382 se
rect -8131 11673 -6718 12382
tri -6718 11673 -6009 12382 nw
tri -6009 11673 -5300 12382 se
rect -5300 12228 -1739 12382
tri -1739 12228 -1465 12502 sw
rect -5300 12127 -1453 12228
rect -5300 11871 -3966 12127
rect -3710 11871 -3442 12127
rect -3186 11871 -2888 12127
rect -2632 11871 -2334 12127
rect -2078 11871 -1810 12127
rect -1554 11871 -1453 12127
rect -5300 11673 -1453 11871
rect -8131 11089 -7302 11673
tri -7302 11089 -6718 11673 nw
tri -6593 11089 -6009 11673 se
rect -6009 11633 -1453 11673
rect -6009 11377 -3966 11633
rect -3710 11377 -3442 11633
rect -3186 11377 -2888 11633
rect -2632 11377 -2334 11633
rect -2078 11377 -1810 11633
rect -1554 11377 -1453 11633
rect -6009 11276 -1453 11377
rect -6009 11089 -1739 11276
rect -8131 10380 -8011 11089
tri -8011 10380 -7302 11089 nw
tri -7302 10380 -6593 11089 se
rect -6593 11002 -1739 11089
tri -1739 11002 -1465 11276 nw
rect -6593 10380 -5180 11002
tri -5180 10380 -4558 11002 nw
tri -1313 10500 689 12502 se
rect 689 12375 5180 12502
tri 5180 12375 5307 12502 sw
tri 5387 12375 6016 13004 ne
tri 6016 12375 8138 14497 sw
rect 689 11666 5307 12375
tri 5307 11666 6016 12375 sw
tri 6016 11666 6725 12375 ne
rect 6725 11666 8138 12375
rect 689 11002 6016 11666
rect 689 10500 809 11002
tri 809 10500 1311 11002 nw
tri 4558 10500 5060 11002 ne
rect 5060 10962 6016 11002
tri 6016 10962 6720 11666 sw
tri 6725 10962 7429 11666 ne
rect 7429 10962 8138 11666
rect 5060 10500 6720 10962
tri -4471 10380 -4351 10500 se
rect -4351 10380 -691 10500
tri -8131 10260 -8011 10380 nw
tri -7422 10260 -7302 10380 se
rect -7302 10260 -5889 10380
tri -12375 8138 -10253 10260 se
rect -10253 9551 -8840 10260
tri -8840 9551 -8131 10260 nw
tri -8131 9551 -7422 10260 se
rect -7422 9671 -5889 10260
tri -5889 9671 -5180 10380 nw
tri -5180 9671 -4471 10380 se
rect -4471 9671 -691 10380
rect -7422 9551 -6473 9671
rect -10253 8967 -9424 9551
tri -9424 8967 -8840 9551 nw
tri -8715 8967 -8131 9551 se
rect -8131 9087 -6473 9551
tri -6473 9087 -5889 9671 nw
tri -5764 9087 -5180 9671 se
rect -5180 9087 -691 9671
rect -8131 8967 -7182 9087
rect -10253 8258 -10133 8967
tri -10133 8258 -9424 8967 nw
tri -9424 8258 -8715 8967 se
rect -8715 8378 -7182 8967
tri -7182 8378 -6473 9087 nw
tri -6473 8378 -5764 9087 se
rect -5764 9000 -691 9087
tri -691 9000 809 10500 nw
tri 1410 10226 1684 10500 se
rect 1684 10226 4351 10500
rect 1410 10133 4351 10226
tri 4351 10133 4718 10500 sw
tri 5060 10133 5427 10500 ne
rect 5427 10253 6720 10500
tri 6720 10253 7429 10962 sw
tri 7429 10253 8138 10962 ne
tri 8138 10253 10260 12375 sw
rect 5427 10133 7429 10253
rect 1410 10124 4718 10133
rect 1410 9868 1511 10124
rect 1767 9868 2035 10124
rect 2291 9868 2589 10124
rect 2845 9868 3143 10124
rect 3399 9868 3667 10124
rect 3923 9868 4718 10124
rect 1410 9630 4718 9868
rect 1410 9374 1511 9630
rect 1767 9374 2035 9630
rect 2291 9374 2589 9630
rect 2845 9374 3143 9630
rect 3399 9374 3667 9630
rect 3923 9424 4718 9630
tri 4718 9424 5427 10133 sw
tri 5427 9424 6136 10133 ne
rect 6136 9544 7429 10133
tri 7429 9544 8138 10253 sw
tri 8138 9544 8847 10253 ne
rect 8847 9544 10260 10253
rect 6136 9424 8138 9544
rect 3923 9374 5427 9424
rect 1410 9274 5427 9374
tri 1410 9000 1684 9274 ne
rect 1684 9000 5427 9274
rect -5764 8378 -4471 9000
rect -8715 8258 -7302 8378
tri -7302 8258 -7182 8378 nw
tri -6593 8258 -6473 8378 se
rect -6473 8258 -4471 8378
tri -4471 8258 -3729 9000 nw
tri 3729 8378 4351 9000 ne
rect 4351 8715 5427 9000
tri 5427 8715 6136 9424 sw
tri 6136 8715 6845 9424 ne
rect 6845 8840 8138 9424
tri 8138 8840 8842 9544 sw
tri 8847 8840 9551 9544 ne
rect 9551 8840 10260 9544
rect 6845 8715 8842 8840
rect 4351 8378 6136 8715
tri -10253 8138 -10133 8258 nw
tri -9544 8138 -9424 8258 se
rect -9424 8138 -8011 8258
tri -14497 6016 -12375 8138 se
rect -12375 7429 -10962 8138
tri -10962 7429 -10253 8138 nw
tri -10253 7429 -9544 8138 se
rect -9544 7549 -8011 8138
tri -8011 7549 -7302 8258 nw
tri -7302 7549 -6593 8258 se
rect -6593 7549 -6473 8258
rect -9544 7429 -8595 7549
rect -12375 6845 -11546 7429
tri -11546 6845 -10962 7429 nw
tri -10837 6845 -10253 7429 se
rect -10253 6965 -8595 7429
tri -8595 6965 -8011 7549 nw
tri -7886 6965 -7302 7549 se
rect -7302 6965 -6473 7549
rect -10253 6845 -9304 6965
rect -12375 6136 -12255 6845
tri -12255 6136 -11546 6845 nw
tri -11546 6136 -10837 6845 se
rect -10837 6256 -9304 6845
tri -9304 6256 -8595 6965 nw
tri -8595 6256 -7886 6965 se
rect -7886 6256 -6473 6965
tri -6473 6256 -4471 8258 nw
tri 4351 7302 5427 8378 ne
rect 5427 8011 6136 8378
tri 6136 8011 6840 8715 sw
tri 6845 8011 7549 8715 ne
rect 7549 8131 8842 8715
tri 8842 8131 9551 8840 sw
tri 9551 8131 10260 8840 ne
tri 10260 8131 12382 10253 sw
rect 7549 8011 9551 8131
rect 5427 7302 6840 8011
tri 6840 7302 7549 8011 sw
tri 7549 7302 8258 8011 ne
rect 8258 7422 9551 8011
tri 9551 7422 10260 8131 sw
tri 10260 7422 10969 8131 ne
rect 10969 7422 12382 8131
rect 8258 7302 10260 7422
tri 5427 6473 6256 7302 ne
rect 6256 6593 7549 7302
tri 7549 6593 8258 7302 sw
tri 8258 6593 8967 7302 ne
rect 8967 6718 10260 7302
tri 10260 6718 10964 7422 sw
tri 10969 6718 11673 7422 ne
rect 11673 6718 12382 7422
rect 8967 6593 10964 6718
rect 6256 6473 8258 6593
rect -10837 6136 -9424 6256
tri -9424 6136 -9304 6256 nw
tri -8715 6136 -8595 6256 se
rect -8595 6136 -6593 6256
tri -6593 6136 -6473 6256 nw
tri -12375 6016 -12255 6136 nw
tri -11666 6016 -11546 6136 se
rect -11546 6016 -10133 6136
tri -14504 6009 -14497 6016 se
rect -14497 6009 -12382 6016
tri -12382 6009 -12375 6016 nw
tri -11673 6009 -11666 6016 se
rect -11666 6009 -10133 6016
rect -14504 -6009 -13004 6009
tri -13004 5387 -12382 6009 nw
tri -12382 5300 -11673 6009 se
rect -11673 5427 -10133 6009
tri -10133 5427 -9424 6136 nw
tri -9424 5427 -8715 6136 se
rect -8715 5427 -8378 6136
rect -11673 5300 -10380 5427
tri -12502 5180 -12382 5300 se
rect -12382 5180 -10380 5300
tri -10380 5180 -10133 5427 nw
tri -9671 5180 -9424 5427 se
rect -9424 5180 -8378 5427
rect -12502 -5180 -11002 5180
tri -11002 4558 -10380 5180 nw
tri -10380 4471 -9671 5180 se
rect -9671 4471 -8378 5180
tri -10500 4351 -10380 4471 se
rect -10380 4351 -8378 4471
tri -8378 4351 -6593 6136 nw
tri 6256 5180 7549 6473 ne
rect 7549 5889 8258 6473
tri 8258 5889 8962 6593 sw
tri 8967 5889 9671 6593 ne
rect 9671 6009 10964 6593
tri 10964 6009 11673 6718 sw
tri 11673 6009 12382 6718 ne
tri 12382 6009 14504 8131 sw
rect 9671 5889 11673 6009
rect 7549 5180 8962 5889
tri 8962 5180 9671 5889 sw
tri 9671 5180 10380 5889 ne
rect 10380 5300 11673 5889
tri 11673 5300 12382 6009 sw
tri 12382 5387 13004 6009 ne
rect 10380 5180 12382 5300
tri 12382 5180 12502 5300 sw
rect -10500 750 -9000 4351
tri -9000 3729 -8378 4351 nw
tri 7549 3729 9000 5180 ne
rect 9000 4471 9671 5180
tri 9671 4471 10380 5180 sw
tri 10380 4558 11002 5180 ne
rect 9000 4351 10380 4471
tri 10380 4351 10500 4471 sw
rect -10500 375 8000 750
rect -10500 119 6552 375
rect 6808 119 7076 375
rect 7332 119 7630 375
rect 7886 119 8000 375
rect -10500 -119 8000 119
rect -10500 -375 6552 -119
rect 6808 -375 7076 -119
rect 7332 -375 7630 -119
rect 7886 -375 8000 -119
rect -10500 -750 8000 -375
rect -10500 -4351 -9000 -750
tri -9000 -4351 -8378 -3729 sw
tri 8378 -4351 9000 -3729 se
rect 9000 -4351 10500 4351
tri -10500 -4471 -10380 -4351 ne
rect -10380 -4471 -8378 -4351
tri -11002 -5180 -10380 -4558 sw
tri -10380 -5180 -9671 -4471 ne
rect -9671 -5180 -8378 -4471
tri -12502 -5300 -12382 -5180 ne
rect -12382 -5300 -10380 -5180
tri -13004 -6009 -12382 -5387 sw
tri -12382 -6009 -11673 -5300 ne
rect -11673 -5889 -10380 -5300
tri -10380 -5889 -9671 -5180 sw
tri -9671 -5889 -8962 -5180 ne
rect -8962 -5889 -8378 -5180
rect -11673 -6009 -9671 -5889
tri -14504 -8131 -12382 -6009 ne
tri -12382 -6718 -11673 -6009 sw
tri -11673 -6718 -10964 -6009 ne
rect -10964 -6473 -9671 -6009
tri -9671 -6473 -9087 -5889 sw
tri -8962 -6473 -8378 -5889 ne
tri -8378 -6473 -6256 -4351 sw
tri 6473 -6256 8378 -4351 se
rect 8378 -4471 10380 -4351
tri 10380 -4471 10500 -4351 nw
rect 8378 -5180 9671 -4471
tri 9671 -5180 10380 -4471 nw
tri 10380 -5180 11002 -4558 se
rect 11002 -5180 12502 5180
rect 13004 3250 14504 6009
rect 13004 1750 15500 3250
rect 8378 -5427 9424 -5180
tri 9424 -5427 9671 -5180 nw
tri 10133 -5427 10380 -5180 se
rect 10380 -5300 12382 -5180
tri 12382 -5300 12502 -5180 nw
rect 13004 -3250 15500 -1750
rect 10380 -5427 11673 -5300
rect 8378 -6136 8715 -5427
tri 8715 -6136 9424 -5427 nw
tri 9424 -6136 10133 -5427 se
rect 10133 -6009 11673 -5427
tri 11673 -6009 12382 -5300 nw
tri 12382 -6009 13004 -5387 se
rect 13004 -6009 14504 -3250
rect 10133 -6136 11546 -6009
tri 11546 -6136 11673 -6009 nw
tri 12375 -6016 12382 -6009 se
rect 12382 -6016 14497 -6009
tri 14497 -6016 14504 -6009 nw
tri 12255 -6136 12375 -6016 se
rect 8378 -6256 8595 -6136
tri 8595 -6256 8715 -6136 nw
tri 9304 -6256 9424 -6136 se
rect 9424 -6256 10837 -6136
rect -10964 -6593 -9087 -6473
tri -9087 -6593 -8967 -6473 sw
tri -8378 -6593 -8258 -6473 ne
rect -8258 -6593 -6256 -6473
rect -10964 -6718 -8967 -6593
rect -12382 -7422 -11673 -6718
tri -11673 -7422 -10969 -6718 sw
tri -10964 -7422 -10260 -6718 ne
rect -10260 -7302 -8967 -6718
tri -8967 -7302 -8258 -6593 sw
tri -8258 -7302 -7549 -6593 ne
rect -7549 -7302 -6256 -6593
rect -10260 -7422 -8258 -7302
rect -12382 -8131 -10969 -7422
tri -10969 -8131 -10260 -7422 sw
tri -10260 -8131 -9551 -7422 ne
rect -9551 -8011 -8258 -7422
tri -8258 -8011 -7549 -7302 sw
tri -7549 -8011 -6840 -7302 ne
rect -6840 -8011 -6256 -7302
rect -9551 -8131 -7549 -8011
tri -12382 -10253 -10260 -8131 ne
tri -10260 -8840 -9551 -8131 sw
tri -9551 -8840 -8842 -8131 ne
rect -8842 -8595 -7549 -8131
tri -7549 -8595 -6965 -8011 sw
tri -6840 -8595 -6256 -8011 ne
tri -6256 -8595 -4134 -6473 sw
tri 4351 -8378 6473 -6256 se
rect 6473 -6965 7886 -6256
tri 7886 -6965 8595 -6256 nw
tri 8595 -6965 9304 -6256 se
rect 9304 -6845 10837 -6256
tri 10837 -6845 11546 -6136 nw
tri 11546 -6845 12255 -6136 se
rect 12255 -6845 12375 -6136
rect 9304 -6965 10253 -6845
rect 6473 -7549 7302 -6965
tri 7302 -7549 7886 -6965 nw
tri 8011 -7549 8595 -6965 se
rect 8595 -7429 10253 -6965
tri 10253 -7429 10837 -6845 nw
tri 10962 -7429 11546 -6845 se
rect 11546 -7429 12375 -6845
rect 8595 -7549 9544 -7429
rect 6473 -8258 6593 -7549
tri 6593 -8258 7302 -7549 nw
tri 7302 -8258 8011 -7549 se
rect 8011 -8138 9544 -7549
tri 9544 -8138 10253 -7429 nw
tri 10253 -8138 10962 -7429 se
rect 10962 -8138 12375 -7429
tri 12375 -8138 14497 -6016 nw
rect 8011 -8258 9424 -8138
tri 9424 -8258 9544 -8138 nw
tri 10133 -8258 10253 -8138 se
tri 6473 -8378 6593 -8258 nw
tri 7182 -8378 7302 -8258 se
rect 7302 -8378 8715 -8258
rect -8842 -8715 -6965 -8595
tri -6965 -8715 -6845 -8595 sw
tri -6256 -8715 -6136 -8595 ne
rect -6136 -8715 -4134 -8595
rect -8842 -8840 -6845 -8715
rect -10260 -9544 -9551 -8840
tri -9551 -9544 -8847 -8840 sw
tri -8842 -9544 -8138 -8840 ne
rect -8138 -9424 -6845 -8840
tri -6845 -9424 -6136 -8715 sw
tri -6136 -9424 -5427 -8715 ne
rect -5427 -9000 -4134 -8715
tri -4134 -9000 -3729 -8595 sw
tri 3729 -9000 4351 -8378 se
rect 4351 -9000 5764 -8378
rect -5427 -9087 5764 -9000
tri 5764 -9087 6473 -8378 nw
tri 6473 -9087 7182 -8378 se
rect 7182 -8967 8715 -8378
tri 8715 -8967 9424 -8258 nw
tri 9424 -8967 10133 -8258 se
rect 10133 -8967 10253 -8258
rect 7182 -9087 8131 -8967
rect -5427 -9424 5180 -9087
rect -8138 -9544 -6136 -9424
rect -10260 -10253 -8847 -9544
tri -8847 -10253 -8138 -9544 sw
tri -8138 -10253 -7429 -9544 ne
rect -7429 -10133 -6136 -9544
tri -6136 -10133 -5427 -9424 sw
tri -5427 -10133 -4718 -9424 ne
rect -4718 -9671 5180 -9424
tri 5180 -9671 5764 -9087 nw
tri 5889 -9671 6473 -9087 se
rect 6473 -9551 8131 -9087
tri 8131 -9551 8715 -8967 nw
tri 8840 -9551 9424 -8967 se
rect 9424 -9551 10253 -8967
rect 6473 -9671 7422 -9551
rect -4718 -10133 4471 -9671
rect -7429 -10253 -5427 -10133
tri -10260 -12375 -8138 -10253 ne
tri -8138 -10962 -7429 -10253 sw
tri -7429 -10962 -6720 -10253 ne
rect -6720 -10500 -5427 -10253
tri -5427 -10500 -5060 -10133 sw
tri -4718 -10500 -4351 -10133 ne
rect -4351 -10380 4471 -10133
tri 4471 -10380 5180 -9671 nw
tri 5180 -10380 5889 -9671 se
rect 5889 -10260 7422 -9671
tri 7422 -10260 8131 -9551 nw
tri 8131 -10260 8840 -9551 se
rect 8840 -10260 10253 -9551
tri 10253 -10260 12375 -8138 nw
rect 5889 -10380 7302 -10260
tri 7302 -10380 7422 -10260 nw
tri 8011 -10380 8131 -10260 se
rect -4351 -10500 4351 -10380
tri 4351 -10500 4471 -10380 nw
rect -6720 -10962 -5060 -10500
rect -8138 -11666 -7429 -10962
tri -7429 -11666 -6725 -10962 sw
tri -6720 -11666 -6016 -10962 ne
rect -6016 -11004 -5060 -10962
tri -5060 -11004 -4556 -10500 sw
tri 4558 -11002 5180 -10380 se
rect 5180 -11002 6593 -10380
rect -6016 -11666 -689 -11004
rect -8138 -12375 -6725 -11666
tri -6725 -12375 -6016 -11666 sw
tri -6016 -12375 -5307 -11666 ne
rect -5307 -12375 -689 -11666
tri -8138 -14497 -6016 -12375 ne
tri -6016 -12502 -5889 -12375 sw
tri -5307 -12502 -5180 -12375 ne
rect -5180 -12502 -689 -12375
tri -689 -12502 809 -11004 sw
tri 1311 -11276 1585 -11002 se
rect 1585 -11089 6593 -11002
tri 6593 -11089 7302 -10380 nw
tri 7302 -11089 8011 -10380 se
rect 8011 -11089 8131 -10380
rect 1585 -11276 6009 -11089
rect 1311 -11377 6009 -11276
rect 1311 -11633 1410 -11377
rect 1666 -11633 1934 -11377
rect 2190 -11633 2488 -11377
rect 2744 -11633 3042 -11377
rect 3298 -11633 3566 -11377
rect 3822 -11633 6009 -11377
rect 1311 -11673 6009 -11633
tri 6009 -11673 6593 -11089 nw
tri 6718 -11673 7302 -11089 se
rect 7302 -11673 8131 -11089
rect 1311 -11871 5300 -11673
rect 1311 -12127 1410 -11871
rect 1666 -12127 1934 -11871
rect 2190 -12127 2488 -11871
rect 2744 -12127 3042 -11871
rect 3298 -12127 3566 -11871
rect 3822 -12127 5300 -11871
rect 1311 -12228 5300 -12127
tri 1311 -12502 1585 -12228 ne
rect 1585 -12382 5300 -12228
tri 5300 -12382 6009 -11673 nw
tri 6009 -12382 6718 -11673 se
rect 6718 -12382 8131 -11673
tri 8131 -12382 10253 -10260 nw
rect 1585 -12502 5180 -12382
tri 5180 -12502 5300 -12382 nw
rect -6016 -13004 -5889 -12502
tri -5889 -13004 -5387 -12502 sw
rect -6016 -13278 -1783 -13004
tri -1783 -13278 -1509 -13004 sw
rect -6016 -13377 -1509 -13278
rect -6016 -13633 -4024 -13377
rect -3768 -13633 -3500 -13377
rect -3244 -13633 -2946 -13377
rect -2690 -13633 -2392 -13377
rect -2136 -13633 -1868 -13377
rect -1612 -13633 -1509 -13377
rect -6016 -13871 -1509 -13633
rect -6016 -14127 -4024 -13871
rect -3768 -14127 -3500 -13871
rect -3244 -14127 -2946 -13871
rect -2690 -14127 -2392 -13871
rect -2136 -14127 -1868 -13871
rect -1612 -14127 -1509 -13871
rect -6016 -14230 -1509 -14127
rect -6016 -14497 -1783 -14230
tri -6016 -14504 -6009 -14497 ne
rect -6009 -14504 -1783 -14497
tri -1783 -14504 -1509 -14230 nw
tri -1313 -14504 689 -12502 ne
rect 689 -13004 809 -12502
tri 809 -13004 1311 -12502 sw
tri 5387 -13004 6009 -12382 se
rect 689 -14504 6009 -13004
tri 6009 -14504 8131 -12382 nw
<< comment >>
tri -6009 6009 -2490 14504 ne
rect -2490 6009 2490 14504
tri 2490 6009 6009 14504 nw
tri -14504 1031 -2490 6009 sw
tri -2490 1031 -427 6009 ne
rect -427 1032 428 6009
tri 428 1032 2490 6009 nw
tri 2491 1032 14504 6009 se
rect -427 1031 73 1032
rect -14504 176 -2489 1031
tri -2489 176 -427 1031 sw
tri -427 176 -73 1031 ne
rect -73 177 73 1031
tri 73 177 428 1032 nw
tri 428 177 2490 1032 se
rect 2490 177 14504 1032
rect -73 176 12 177
rect -14504 30 -425 176
tri -425 30 -73 176 sw
tri -73 30 -12 176 ne
rect -12 30 12 176
tri 12 30 73 177 nw
tri 73 30 427 177 se
rect 427 30 14504 177
rect -14504 4 -73 30
tri -73 4 -12 30 sw
tri -12 4 -2 30 ne
rect -2 5 2 30
tri 2 5 12 30 nw
tri 12 5 72 30 se
rect 72 5 14504 30
rect -2 4 0 5
rect -14504 0 -10 4
tri -10 0 -2 4 sw
tri -2 0 0 4 ne
tri 0 1 2 5 nw
tri 2 1 12 5 se
rect 12 1 14504 5
tri 0 0 2 1 se
rect 2 0 14504 1
rect -14504 -1 -2 0
tri -2 -1 0 0 nw
tri 0 -1 1 0 ne
rect 1 -1 14504 0
rect -14504 -5 -12 -1
tri -12 -5 -2 -1 nw
tri -2 -5 0 -1 se
tri 0 -2 1 -1 sw
tri 1 -2 3 -1 ne
rect 3 -2 14504 -1
rect 0 -5 1 -2
rect -14504 -30 -72 -5
tri -72 -30 -12 -5 nw
tri -12 -30 -2 -5 se
rect -2 -6 1 -5
tri 1 -6 3 -2 sw
tri 4 -6 13 -2 ne
rect 13 -6 14504 -2
rect -2 -30 3 -6
rect -14504 -177 -427 -30
tri -427 -177 -73 -30 nw
tri -73 -177 -12 -30 se
rect -12 -31 3 -30
tri 3 -31 13 -6 sw
tri 14 -31 74 -6 ne
rect 74 -31 14504 -6
rect -12 -177 13 -31
rect -14504 -1032 -2490 -177
tri -2490 -1032 -428 -177 nw
tri -428 -1032 -73 -177 se
rect -73 -178 13 -177
tri 13 -178 74 -31 sw
tri 74 -178 428 -31 ne
rect 428 -178 14504 -31
rect -73 -1032 74 -178
tri 74 -1032 428 -178 sw
tri 429 -1032 2490 -178 ne
rect 2490 -1032 14504 -178
tri -14504 -6009 -2491 -1032 nw
tri -2490 -6009 -428 -1032 se
rect -428 -6009 428 -1032
tri 428 -6009 2490 -1032 sw
tri 2490 -6009 14504 -1032 ne
tri -6009 -14504 -2490 -6009 se
rect -2490 -14504 2490 -6009
tri 2490 -14504 6009 -6009 sw
<< properties >>
string GDS_END 10392512
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 10385804
string gencell sky130_fd_pr__rf_test_coil1
string library sky130
string parameter m=1
string path 343.850 -150.225 343.850 -43.750 
<< end >>
