magic
tech sky130B
timestamp 1676037725
<< properties >>
string GDS_END 29563964
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 29563256
<< end >>
