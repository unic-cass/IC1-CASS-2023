magic
tech sky130A
magscale 1 2
timestamp 1698611444
<< obsli1 >>
rect 1104 2159 85652 86513
<< obsm1 >>
rect 474 1572 85712 86760
<< metal2 >>
rect 2410 88182 2466 88982
rect 4894 88182 4950 88982
rect 7378 88182 7434 88982
rect 9862 88182 9918 88982
rect 12346 88182 12402 88982
rect 14830 88182 14886 88982
rect 17314 88182 17370 88982
rect 19798 88182 19854 88982
rect 22282 88182 22338 88982
rect 24766 88182 24822 88982
rect 27250 88182 27306 88982
rect 29734 88182 29790 88982
rect 32218 88182 32274 88982
rect 34702 88182 34758 88982
rect 37186 88182 37242 88982
rect 39670 88182 39726 88982
rect 42154 88182 42210 88982
rect 44638 88182 44694 88982
rect 47122 88182 47178 88982
rect 49606 88182 49662 88982
rect 52090 88182 52146 88982
rect 54574 88182 54630 88982
rect 57058 88182 57114 88982
rect 59542 88182 59598 88982
rect 62026 88182 62082 88982
rect 64510 88182 64566 88982
rect 66994 88182 67050 88982
rect 69478 88182 69534 88982
rect 71962 88182 72018 88982
rect 74446 88182 74502 88982
rect 76930 88182 76986 88982
rect 79414 88182 79470 88982
rect 81898 88182 81954 88982
rect 84382 88182 84438 88982
rect 8758 0 8814 800
rect 26054 0 26110 800
rect 43350 0 43406 800
rect 60646 0 60702 800
rect 77942 0 77998 800
<< obsm2 >>
rect 480 88126 2354 88210
rect 2522 88126 4838 88210
rect 5006 88126 7322 88210
rect 7490 88126 9806 88210
rect 9974 88126 12290 88210
rect 12458 88126 14774 88210
rect 14942 88126 17258 88210
rect 17426 88126 19742 88210
rect 19910 88126 22226 88210
rect 22394 88126 24710 88210
rect 24878 88126 27194 88210
rect 27362 88126 29678 88210
rect 29846 88126 32162 88210
rect 32330 88126 34646 88210
rect 34814 88126 37130 88210
rect 37298 88126 39614 88210
rect 39782 88126 42098 88210
rect 42266 88126 44582 88210
rect 44750 88126 47066 88210
rect 47234 88126 49550 88210
rect 49718 88126 52034 88210
rect 52202 88126 54518 88210
rect 54686 88126 57002 88210
rect 57170 88126 59486 88210
rect 59654 88126 61970 88210
rect 62138 88126 64454 88210
rect 64622 88126 66938 88210
rect 67106 88126 69422 88210
rect 69590 88126 71906 88210
rect 72074 88126 74390 88210
rect 74558 88126 76874 88210
rect 77042 88126 79358 88210
rect 79526 88126 81842 88210
rect 82010 88126 84326 88210
rect 84494 88126 85542 88210
rect 480 856 85542 88126
rect 480 734 8702 856
rect 8870 734 25998 856
rect 26166 734 43294 856
rect 43462 734 60590 856
rect 60758 734 77886 856
rect 78054 734 85542 856
<< metal3 >>
rect 0 87048 800 87168
rect 86038 86776 86838 86896
rect 0 85688 800 85808
rect 0 84328 800 84448
rect 86038 83240 86838 83360
rect 0 82968 800 83088
rect 0 81608 800 81728
rect 0 80248 800 80368
rect 86038 79704 86838 79824
rect 0 78888 800 79008
rect 0 77528 800 77648
rect 0 76168 800 76288
rect 86038 76168 86838 76288
rect 0 74808 800 74928
rect 0 73448 800 73568
rect 86038 72632 86838 72752
rect 0 72088 800 72208
rect 0 70728 800 70848
rect 0 69368 800 69488
rect 86038 69096 86838 69216
rect 0 68008 800 68128
rect 0 66648 800 66768
rect 86038 65560 86838 65680
rect 0 65288 800 65408
rect 0 63928 800 64048
rect 0 62568 800 62688
rect 86038 62024 86838 62144
rect 0 61208 800 61328
rect 0 59848 800 59968
rect 0 58488 800 58608
rect 86038 58488 86838 58608
rect 0 57128 800 57248
rect 0 55768 800 55888
rect 86038 54952 86838 55072
rect 0 54408 800 54528
rect 0 53048 800 53168
rect 0 51688 800 51808
rect 86038 51416 86838 51536
rect 0 50328 800 50448
rect 0 48968 800 49088
rect 86038 47880 86838 48000
rect 0 47608 800 47728
rect 0 46248 800 46368
rect 0 44888 800 45008
rect 86038 44344 86838 44464
rect 0 43528 800 43648
rect 0 42168 800 42288
rect 0 40808 800 40928
rect 86038 40808 86838 40928
rect 0 39448 800 39568
rect 0 38088 800 38208
rect 86038 37272 86838 37392
rect 0 36728 800 36848
rect 0 35368 800 35488
rect 0 34008 800 34128
rect 86038 33736 86838 33856
rect 0 32648 800 32768
rect 0 31288 800 31408
rect 86038 30200 86838 30320
rect 0 29928 800 30048
rect 0 28568 800 28688
rect 0 27208 800 27328
rect 86038 26664 86838 26784
rect 0 25848 800 25968
rect 0 24488 800 24608
rect 0 23128 800 23248
rect 86038 23128 86838 23248
rect 0 21768 800 21888
rect 0 20408 800 20528
rect 86038 19592 86838 19712
rect 0 19048 800 19168
rect 0 17688 800 17808
rect 0 16328 800 16448
rect 86038 16056 86838 16176
rect 0 14968 800 15088
rect 0 13608 800 13728
rect 86038 12520 86838 12640
rect 0 12248 800 12368
rect 0 10888 800 11008
rect 0 9528 800 9648
rect 86038 8984 86838 9104
rect 0 8168 800 8288
rect 0 6808 800 6928
rect 0 5448 800 5568
rect 86038 5448 86838 5568
rect 0 4088 800 4208
rect 0 2728 800 2848
rect 86038 1912 86838 2032
rect 0 1368 800 1488
<< obsm3 >>
rect 880 86976 86038 87138
rect 880 86968 85958 86976
rect 606 86696 85958 86968
rect 606 85888 86038 86696
rect 880 85608 86038 85888
rect 606 84528 86038 85608
rect 880 84248 86038 84528
rect 606 83440 86038 84248
rect 606 83168 85958 83440
rect 880 83160 85958 83168
rect 880 82888 86038 83160
rect 606 81808 86038 82888
rect 880 81528 86038 81808
rect 606 80448 86038 81528
rect 880 80168 86038 80448
rect 606 79904 86038 80168
rect 606 79624 85958 79904
rect 606 79088 86038 79624
rect 880 78808 86038 79088
rect 606 77728 86038 78808
rect 880 77448 86038 77728
rect 606 76368 86038 77448
rect 880 76088 85958 76368
rect 606 75008 86038 76088
rect 880 74728 86038 75008
rect 606 73648 86038 74728
rect 880 73368 86038 73648
rect 606 72832 86038 73368
rect 606 72552 85958 72832
rect 606 72288 86038 72552
rect 880 72008 86038 72288
rect 606 70928 86038 72008
rect 880 70648 86038 70928
rect 606 69568 86038 70648
rect 880 69296 86038 69568
rect 880 69288 85958 69296
rect 606 69016 85958 69288
rect 606 68208 86038 69016
rect 880 67928 86038 68208
rect 606 66848 86038 67928
rect 880 66568 86038 66848
rect 606 65760 86038 66568
rect 606 65488 85958 65760
rect 880 65480 85958 65488
rect 880 65208 86038 65480
rect 606 64128 86038 65208
rect 880 63848 86038 64128
rect 606 62768 86038 63848
rect 880 62488 86038 62768
rect 606 62224 86038 62488
rect 606 61944 85958 62224
rect 606 61408 86038 61944
rect 880 61128 86038 61408
rect 606 60048 86038 61128
rect 880 59768 86038 60048
rect 606 58688 86038 59768
rect 880 58408 85958 58688
rect 606 57328 86038 58408
rect 880 57048 86038 57328
rect 606 55968 86038 57048
rect 880 55688 86038 55968
rect 606 55152 86038 55688
rect 606 54872 85958 55152
rect 606 54608 86038 54872
rect 880 54328 86038 54608
rect 606 53248 86038 54328
rect 880 52968 86038 53248
rect 606 51888 86038 52968
rect 880 51616 86038 51888
rect 880 51608 85958 51616
rect 606 51336 85958 51608
rect 606 50528 86038 51336
rect 880 50248 86038 50528
rect 606 49168 86038 50248
rect 880 48888 86038 49168
rect 606 48080 86038 48888
rect 606 47808 85958 48080
rect 880 47800 85958 47808
rect 880 47528 86038 47800
rect 606 46448 86038 47528
rect 880 46168 86038 46448
rect 606 45088 86038 46168
rect 880 44808 86038 45088
rect 606 44544 86038 44808
rect 606 44264 85958 44544
rect 606 43728 86038 44264
rect 880 43448 86038 43728
rect 606 42368 86038 43448
rect 880 42088 86038 42368
rect 606 41008 86038 42088
rect 880 40728 85958 41008
rect 606 39648 86038 40728
rect 880 39368 86038 39648
rect 606 38288 86038 39368
rect 880 38008 86038 38288
rect 606 37472 86038 38008
rect 606 37192 85958 37472
rect 606 36928 86038 37192
rect 880 36648 86038 36928
rect 606 35568 86038 36648
rect 880 35288 86038 35568
rect 606 34208 86038 35288
rect 880 33936 86038 34208
rect 880 33928 85958 33936
rect 606 33656 85958 33928
rect 606 32848 86038 33656
rect 880 32568 86038 32848
rect 606 31488 86038 32568
rect 880 31208 86038 31488
rect 606 30400 86038 31208
rect 606 30128 85958 30400
rect 880 30120 85958 30128
rect 880 29848 86038 30120
rect 606 28768 86038 29848
rect 880 28488 86038 28768
rect 606 27408 86038 28488
rect 880 27128 86038 27408
rect 606 26864 86038 27128
rect 606 26584 85958 26864
rect 606 26048 86038 26584
rect 880 25768 86038 26048
rect 606 24688 86038 25768
rect 880 24408 86038 24688
rect 606 23328 86038 24408
rect 880 23048 85958 23328
rect 606 21968 86038 23048
rect 880 21688 86038 21968
rect 606 20608 86038 21688
rect 880 20328 86038 20608
rect 606 19792 86038 20328
rect 606 19512 85958 19792
rect 606 19248 86038 19512
rect 880 18968 86038 19248
rect 606 17888 86038 18968
rect 880 17608 86038 17888
rect 606 16528 86038 17608
rect 880 16256 86038 16528
rect 880 16248 85958 16256
rect 606 15976 85958 16248
rect 606 15168 86038 15976
rect 880 14888 86038 15168
rect 606 13808 86038 14888
rect 880 13528 86038 13808
rect 606 12720 86038 13528
rect 606 12448 85958 12720
rect 880 12440 85958 12448
rect 880 12168 86038 12440
rect 606 11088 86038 12168
rect 880 10808 86038 11088
rect 606 9728 86038 10808
rect 880 9448 86038 9728
rect 606 9184 86038 9448
rect 606 8904 85958 9184
rect 606 8368 86038 8904
rect 880 8088 86038 8368
rect 606 7008 86038 8088
rect 880 6728 86038 7008
rect 606 5648 86038 6728
rect 880 5368 85958 5648
rect 606 4288 86038 5368
rect 880 4008 86038 4288
rect 606 2928 86038 4008
rect 880 2648 86038 2928
rect 606 2112 86038 2648
rect 606 1832 85958 2112
rect 606 1568 86038 1832
rect 880 1395 86038 1568
<< metal4 >>
rect 2344 2128 2664 86544
rect 17704 2128 18024 86544
rect 33064 2128 33384 86544
rect 48424 2128 48744 86544
rect 63784 2128 64104 86544
rect 79144 2128 79464 86544
<< obsm4 >>
rect 526 2048 2264 85781
rect 2744 2048 17624 85781
rect 18104 2048 32984 85781
rect 33464 2048 48344 85781
rect 48824 2048 63704 85781
rect 64184 2048 79064 85781
rect 79544 2048 83010 85781
rect 526 1939 83010 2048
<< obsm5 >>
rect 484 9020 83052 68500
<< labels >>
rlabel metal3 s 86038 1912 86838 2032 6 buttons
port 1 nsew signal input
rlabel metal2 s 2410 88182 2466 88982 6 clk
port 2 nsew signal input
rlabel metal2 s 7378 88182 7434 88982 6 i_wb_addr[0]
port 3 nsew signal input
rlabel metal2 s 32218 88182 32274 88982 6 i_wb_addr[10]
port 4 nsew signal input
rlabel metal2 s 34702 88182 34758 88982 6 i_wb_addr[11]
port 5 nsew signal input
rlabel metal2 s 37186 88182 37242 88982 6 i_wb_addr[12]
port 6 nsew signal input
rlabel metal2 s 39670 88182 39726 88982 6 i_wb_addr[13]
port 7 nsew signal input
rlabel metal2 s 42154 88182 42210 88982 6 i_wb_addr[14]
port 8 nsew signal input
rlabel metal2 s 44638 88182 44694 88982 6 i_wb_addr[15]
port 9 nsew signal input
rlabel metal2 s 47122 88182 47178 88982 6 i_wb_addr[16]
port 10 nsew signal input
rlabel metal2 s 49606 88182 49662 88982 6 i_wb_addr[17]
port 11 nsew signal input
rlabel metal2 s 52090 88182 52146 88982 6 i_wb_addr[18]
port 12 nsew signal input
rlabel metal2 s 54574 88182 54630 88982 6 i_wb_addr[19]
port 13 nsew signal input
rlabel metal2 s 9862 88182 9918 88982 6 i_wb_addr[1]
port 14 nsew signal input
rlabel metal2 s 57058 88182 57114 88982 6 i_wb_addr[20]
port 15 nsew signal input
rlabel metal2 s 59542 88182 59598 88982 6 i_wb_addr[21]
port 16 nsew signal input
rlabel metal2 s 62026 88182 62082 88982 6 i_wb_addr[22]
port 17 nsew signal input
rlabel metal2 s 64510 88182 64566 88982 6 i_wb_addr[23]
port 18 nsew signal input
rlabel metal2 s 66994 88182 67050 88982 6 i_wb_addr[24]
port 19 nsew signal input
rlabel metal2 s 69478 88182 69534 88982 6 i_wb_addr[25]
port 20 nsew signal input
rlabel metal2 s 71962 88182 72018 88982 6 i_wb_addr[26]
port 21 nsew signal input
rlabel metal2 s 74446 88182 74502 88982 6 i_wb_addr[27]
port 22 nsew signal input
rlabel metal2 s 76930 88182 76986 88982 6 i_wb_addr[28]
port 23 nsew signal input
rlabel metal2 s 79414 88182 79470 88982 6 i_wb_addr[29]
port 24 nsew signal input
rlabel metal2 s 12346 88182 12402 88982 6 i_wb_addr[2]
port 25 nsew signal input
rlabel metal2 s 81898 88182 81954 88982 6 i_wb_addr[30]
port 26 nsew signal input
rlabel metal2 s 84382 88182 84438 88982 6 i_wb_addr[31]
port 27 nsew signal input
rlabel metal2 s 14830 88182 14886 88982 6 i_wb_addr[3]
port 28 nsew signal input
rlabel metal2 s 17314 88182 17370 88982 6 i_wb_addr[4]
port 29 nsew signal input
rlabel metal2 s 19798 88182 19854 88982 6 i_wb_addr[5]
port 30 nsew signal input
rlabel metal2 s 22282 88182 22338 88982 6 i_wb_addr[6]
port 31 nsew signal input
rlabel metal2 s 24766 88182 24822 88982 6 i_wb_addr[7]
port 32 nsew signal input
rlabel metal2 s 27250 88182 27306 88982 6 i_wb_addr[8]
port 33 nsew signal input
rlabel metal2 s 29734 88182 29790 88982 6 i_wb_addr[9]
port 34 nsew signal input
rlabel metal2 s 8758 0 8814 800 6 i_wb_cyc
port 35 nsew signal input
rlabel metal3 s 0 1368 800 1488 6 i_wb_data[0]
port 36 nsew signal input
rlabel metal3 s 0 14968 800 15088 6 i_wb_data[10]
port 37 nsew signal input
rlabel metal3 s 0 16328 800 16448 6 i_wb_data[11]
port 38 nsew signal input
rlabel metal3 s 0 17688 800 17808 6 i_wb_data[12]
port 39 nsew signal input
rlabel metal3 s 0 19048 800 19168 6 i_wb_data[13]
port 40 nsew signal input
rlabel metal3 s 0 20408 800 20528 6 i_wb_data[14]
port 41 nsew signal input
rlabel metal3 s 0 21768 800 21888 6 i_wb_data[15]
port 42 nsew signal input
rlabel metal3 s 0 23128 800 23248 6 i_wb_data[16]
port 43 nsew signal input
rlabel metal3 s 0 24488 800 24608 6 i_wb_data[17]
port 44 nsew signal input
rlabel metal3 s 0 25848 800 25968 6 i_wb_data[18]
port 45 nsew signal input
rlabel metal3 s 0 27208 800 27328 6 i_wb_data[19]
port 46 nsew signal input
rlabel metal3 s 0 2728 800 2848 6 i_wb_data[1]
port 47 nsew signal input
rlabel metal3 s 0 28568 800 28688 6 i_wb_data[20]
port 48 nsew signal input
rlabel metal3 s 0 29928 800 30048 6 i_wb_data[21]
port 49 nsew signal input
rlabel metal3 s 0 31288 800 31408 6 i_wb_data[22]
port 50 nsew signal input
rlabel metal3 s 0 32648 800 32768 6 i_wb_data[23]
port 51 nsew signal input
rlabel metal3 s 0 34008 800 34128 6 i_wb_data[24]
port 52 nsew signal input
rlabel metal3 s 0 35368 800 35488 6 i_wb_data[25]
port 53 nsew signal input
rlabel metal3 s 0 36728 800 36848 6 i_wb_data[26]
port 54 nsew signal input
rlabel metal3 s 0 38088 800 38208 6 i_wb_data[27]
port 55 nsew signal input
rlabel metal3 s 0 39448 800 39568 6 i_wb_data[28]
port 56 nsew signal input
rlabel metal3 s 0 40808 800 40928 6 i_wb_data[29]
port 57 nsew signal input
rlabel metal3 s 0 4088 800 4208 6 i_wb_data[2]
port 58 nsew signal input
rlabel metal3 s 0 42168 800 42288 6 i_wb_data[30]
port 59 nsew signal input
rlabel metal3 s 0 43528 800 43648 6 i_wb_data[31]
port 60 nsew signal input
rlabel metal3 s 0 5448 800 5568 6 i_wb_data[3]
port 61 nsew signal input
rlabel metal3 s 0 6808 800 6928 6 i_wb_data[4]
port 62 nsew signal input
rlabel metal3 s 0 8168 800 8288 6 i_wb_data[5]
port 63 nsew signal input
rlabel metal3 s 0 9528 800 9648 6 i_wb_data[6]
port 64 nsew signal input
rlabel metal3 s 0 10888 800 11008 6 i_wb_data[7]
port 65 nsew signal input
rlabel metal3 s 0 12248 800 12368 6 i_wb_data[8]
port 66 nsew signal input
rlabel metal3 s 0 13608 800 13728 6 i_wb_data[9]
port 67 nsew signal input
rlabel metal2 s 26054 0 26110 800 6 i_wb_stb
port 68 nsew signal input
rlabel metal2 s 43350 0 43406 800 6 i_wb_we
port 69 nsew signal input
rlabel metal3 s 86038 5448 86838 5568 6 led_enb[0]
port 70 nsew signal output
rlabel metal3 s 86038 40808 86838 40928 6 led_enb[10]
port 71 nsew signal output
rlabel metal3 s 86038 44344 86838 44464 6 led_enb[11]
port 72 nsew signal output
rlabel metal3 s 86038 8984 86838 9104 6 led_enb[1]
port 73 nsew signal output
rlabel metal3 s 86038 12520 86838 12640 6 led_enb[2]
port 74 nsew signal output
rlabel metal3 s 86038 16056 86838 16176 6 led_enb[3]
port 75 nsew signal output
rlabel metal3 s 86038 19592 86838 19712 6 led_enb[4]
port 76 nsew signal output
rlabel metal3 s 86038 23128 86838 23248 6 led_enb[5]
port 77 nsew signal output
rlabel metal3 s 86038 26664 86838 26784 6 led_enb[6]
port 78 nsew signal output
rlabel metal3 s 86038 30200 86838 30320 6 led_enb[7]
port 79 nsew signal output
rlabel metal3 s 86038 33736 86838 33856 6 led_enb[8]
port 80 nsew signal output
rlabel metal3 s 86038 37272 86838 37392 6 led_enb[9]
port 81 nsew signal output
rlabel metal3 s 86038 47880 86838 48000 6 leds[0]
port 82 nsew signal output
rlabel metal3 s 86038 83240 86838 83360 6 leds[10]
port 83 nsew signal output
rlabel metal3 s 86038 86776 86838 86896 6 leds[11]
port 84 nsew signal output
rlabel metal3 s 86038 51416 86838 51536 6 leds[1]
port 85 nsew signal output
rlabel metal3 s 86038 54952 86838 55072 6 leds[2]
port 86 nsew signal output
rlabel metal3 s 86038 58488 86838 58608 6 leds[3]
port 87 nsew signal output
rlabel metal3 s 86038 62024 86838 62144 6 leds[4]
port 88 nsew signal output
rlabel metal3 s 86038 65560 86838 65680 6 leds[5]
port 89 nsew signal output
rlabel metal3 s 86038 69096 86838 69216 6 leds[6]
port 90 nsew signal output
rlabel metal3 s 86038 72632 86838 72752 6 leds[7]
port 91 nsew signal output
rlabel metal3 s 86038 76168 86838 76288 6 leds[8]
port 92 nsew signal output
rlabel metal3 s 86038 79704 86838 79824 6 leds[9]
port 93 nsew signal output
rlabel metal2 s 60646 0 60702 800 6 o_wb_ack
port 94 nsew signal output
rlabel metal3 s 0 44888 800 45008 6 o_wb_data[0]
port 95 nsew signal output
rlabel metal3 s 0 58488 800 58608 6 o_wb_data[10]
port 96 nsew signal output
rlabel metal3 s 0 59848 800 59968 6 o_wb_data[11]
port 97 nsew signal output
rlabel metal3 s 0 61208 800 61328 6 o_wb_data[12]
port 98 nsew signal output
rlabel metal3 s 0 62568 800 62688 6 o_wb_data[13]
port 99 nsew signal output
rlabel metal3 s 0 63928 800 64048 6 o_wb_data[14]
port 100 nsew signal output
rlabel metal3 s 0 65288 800 65408 6 o_wb_data[15]
port 101 nsew signal output
rlabel metal3 s 0 66648 800 66768 6 o_wb_data[16]
port 102 nsew signal output
rlabel metal3 s 0 68008 800 68128 6 o_wb_data[17]
port 103 nsew signal output
rlabel metal3 s 0 69368 800 69488 6 o_wb_data[18]
port 104 nsew signal output
rlabel metal3 s 0 70728 800 70848 6 o_wb_data[19]
port 105 nsew signal output
rlabel metal3 s 0 46248 800 46368 6 o_wb_data[1]
port 106 nsew signal output
rlabel metal3 s 0 72088 800 72208 6 o_wb_data[20]
port 107 nsew signal output
rlabel metal3 s 0 73448 800 73568 6 o_wb_data[21]
port 108 nsew signal output
rlabel metal3 s 0 74808 800 74928 6 o_wb_data[22]
port 109 nsew signal output
rlabel metal3 s 0 76168 800 76288 6 o_wb_data[23]
port 110 nsew signal output
rlabel metal3 s 0 77528 800 77648 6 o_wb_data[24]
port 111 nsew signal output
rlabel metal3 s 0 78888 800 79008 6 o_wb_data[25]
port 112 nsew signal output
rlabel metal3 s 0 80248 800 80368 6 o_wb_data[26]
port 113 nsew signal output
rlabel metal3 s 0 81608 800 81728 6 o_wb_data[27]
port 114 nsew signal output
rlabel metal3 s 0 82968 800 83088 6 o_wb_data[28]
port 115 nsew signal output
rlabel metal3 s 0 84328 800 84448 6 o_wb_data[29]
port 116 nsew signal output
rlabel metal3 s 0 47608 800 47728 6 o_wb_data[2]
port 117 nsew signal output
rlabel metal3 s 0 85688 800 85808 6 o_wb_data[30]
port 118 nsew signal output
rlabel metal3 s 0 87048 800 87168 6 o_wb_data[31]
port 119 nsew signal output
rlabel metal3 s 0 48968 800 49088 6 o_wb_data[3]
port 120 nsew signal output
rlabel metal3 s 0 50328 800 50448 6 o_wb_data[4]
port 121 nsew signal output
rlabel metal3 s 0 51688 800 51808 6 o_wb_data[5]
port 122 nsew signal output
rlabel metal3 s 0 53048 800 53168 6 o_wb_data[6]
port 123 nsew signal output
rlabel metal3 s 0 54408 800 54528 6 o_wb_data[7]
port 124 nsew signal output
rlabel metal3 s 0 55768 800 55888 6 o_wb_data[8]
port 125 nsew signal output
rlabel metal3 s 0 57128 800 57248 6 o_wb_data[9]
port 126 nsew signal output
rlabel metal2 s 77942 0 77998 800 6 o_wb_stall
port 127 nsew signal output
rlabel metal2 s 4894 88182 4950 88982 6 reset
port 128 nsew signal input
rlabel metal4 s 2344 2128 2664 86544 6 vccd1
port 129 nsew power bidirectional
rlabel metal4 s 33064 2128 33384 86544 6 vccd1
port 129 nsew power bidirectional
rlabel metal4 s 63784 2128 64104 86544 6 vccd1
port 129 nsew power bidirectional
rlabel metal4 s 17704 2128 18024 86544 6 vssd1
port 130 nsew ground bidirectional
rlabel metal4 s 48424 2128 48744 86544 6 vssd1
port 130 nsew ground bidirectional
rlabel metal4 s 79144 2128 79464 86544 6 vssd1
port 130 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 86838 88982
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 28991702
string GDS_FILE /wb_buttons_leds/openlane/wb_buttons_leds/runs/RUN_2023.10.29_19.42.28/results/signoff/wb_buttons_leds.magic.gds
string GDS_START 1413422
<< end >>

