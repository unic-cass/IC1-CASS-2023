magic
tech sky130A
timestamp 1676037725
<< properties >>
string GDS_END 3276418
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 3274878
<< end >>
