* NGSPICE file created from wb_buttons_leds.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_4 abstract view
.subckt sky130_fd_sc_hd__a21bo_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_2 abstract view
.subckt sky130_fd_sc_hd__a311oi_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_2 abstract view
.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_4 abstract view
.subckt sky130_fd_sc_hd__o32ai_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_2 abstract view
.subckt sky130_fd_sc_hd__a32oi_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_1 abstract view
.subckt sky130_fd_sc_hd__a32oi_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_2 abstract view
.subckt sky130_fd_sc_hd__o311ai_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_2 abstract view
.subckt sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

.subckt wb_buttons_leds buttons clk i_wb_addr[0] i_wb_addr[10] i_wb_addr[11] i_wb_addr[12]
+ i_wb_addr[13] i_wb_addr[14] i_wb_addr[15] i_wb_addr[16] i_wb_addr[17] i_wb_addr[18]
+ i_wb_addr[19] i_wb_addr[1] i_wb_addr[20] i_wb_addr[21] i_wb_addr[22] i_wb_addr[23]
+ i_wb_addr[24] i_wb_addr[25] i_wb_addr[26] i_wb_addr[27] i_wb_addr[28] i_wb_addr[29]
+ i_wb_addr[2] i_wb_addr[30] i_wb_addr[31] i_wb_addr[3] i_wb_addr[4] i_wb_addr[5]
+ i_wb_addr[6] i_wb_addr[7] i_wb_addr[8] i_wb_addr[9] i_wb_cyc i_wb_data[0] i_wb_data[10]
+ i_wb_data[11] i_wb_data[12] i_wb_data[13] i_wb_data[14] i_wb_data[15] i_wb_data[16]
+ i_wb_data[17] i_wb_data[18] i_wb_data[19] i_wb_data[1] i_wb_data[20] i_wb_data[21]
+ i_wb_data[22] i_wb_data[23] i_wb_data[24] i_wb_data[25] i_wb_data[26] i_wb_data[27]
+ i_wb_data[28] i_wb_data[29] i_wb_data[2] i_wb_data[30] i_wb_data[31] i_wb_data[3]
+ i_wb_data[4] i_wb_data[5] i_wb_data[6] i_wb_data[7] i_wb_data[8] i_wb_data[9] i_wb_stb
+ i_wb_we led_enb[0] led_enb[10] led_enb[11] led_enb[1] led_enb[2] led_enb[3] led_enb[4]
+ led_enb[5] led_enb[6] led_enb[7] led_enb[8] led_enb[9] leds[0] leds[10] leds[11]
+ leds[1] leds[2] leds[3] leds[4] leds[5] leds[6] leds[7] leds[8] leds[9] o_wb_ack
+ o_wb_data[0] o_wb_data[10] o_wb_data[11] o_wb_data[12] o_wb_data[13] o_wb_data[14]
+ o_wb_data[15] o_wb_data[16] o_wb_data[17] o_wb_data[18] o_wb_data[19] o_wb_data[1]
+ o_wb_data[20] o_wb_data[21] o_wb_data[22] o_wb_data[23] o_wb_data[24] o_wb_data[25]
+ o_wb_data[26] o_wb_data[27] o_wb_data[28] o_wb_data[29] o_wb_data[2] o_wb_data[30]
+ o_wb_data[31] o_wb_data[3] o_wb_data[4] o_wb_data[5] o_wb_data[6] o_wb_data[7] o_wb_data[8]
+ o_wb_data[9] o_wb_stall reset vccd1 vssd1
XFILLER_140_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09671_ _09631_/Y _09666_/B _09674_/B _09670_/X vssd1 vssd1 vccd1 vccd1 _09819_/A
+ sky130_fd_sc_hd__a211oi_2
XFILLER_95_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_556 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09105_ _17425_/A _17423_/A _09172_/B _09502_/B vssd1 vssd1 vccd1 vccd1 _09106_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_163_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09036_ _17081_/A _09031_/A _09031_/B vssd1 vssd1 vccd1 vccd1 _09039_/A sky130_fd_sc_hd__o21ba_1
XFILLER_164_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_355 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout820 _09265_/C vssd1 vssd1 vccd1 vccd1 _15208_/A sky130_fd_sc_hd__buf_2
XFILLER_131_252 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout831 _17486_/Q vssd1 vssd1 vccd1 vccd1 _14851_/A sky130_fd_sc_hd__buf_2
X_09938_ _10560_/A _10072_/B _09803_/C vssd1 vssd1 vccd1 vccd1 _09939_/B sky130_fd_sc_hd__a21oi_1
Xfanout842 _17485_/Q vssd1 vssd1 vccd1 vccd1 _11387_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_120_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout853 _09128_/B vssd1 vssd1 vccd1 vccd1 _12127_/C sky130_fd_sc_hd__clkbuf_4
Xfanout864 _17306_/A1 vssd1 vssd1 vccd1 vccd1 _12127_/D sky130_fd_sc_hd__clkbuf_4
Xfanout875 _09981_/D vssd1 vssd1 vccd1 vccd1 _10067_/B sky130_fd_sc_hd__buf_2
XFILLER_133_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout886 _11592_/B vssd1 vssd1 vccd1 vccd1 _15042_/B sky130_fd_sc_hd__buf_2
X_09869_ _09870_/A _09870_/B _09870_/C vssd1 vssd1 vccd1 vccd1 _09869_/X sky130_fd_sc_hd__a21o_1
XFILLER_92_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout897 _11468_/D vssd1 vssd1 vccd1 vccd1 _15008_/A sky130_fd_sc_hd__buf_2
XTAP_3202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11900_ _17385_/A _17383_/A _12258_/B _11900_/D vssd1 vssd1 vccd1 vccd1 _11901_/B
+ sky130_fd_sc_hd__and4_1
XTAP_3235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12880_ _12881_/A _12881_/B vssd1 vssd1 vccd1 vccd1 _13040_/B sky130_fd_sc_hd__nor2_1
XFILLER_45_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11831_ _11837_/A _11831_/B vssd1 vssd1 vccd1 vccd1 _11831_/Y sky130_fd_sc_hd__nand2_1
XFILLER_61_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14550_ _14599_/B _14708_/D vssd1 vssd1 vccd1 vccd1 _14679_/B sky130_fd_sc_hd__nand2_1
XTAP_2578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11762_ _11762_/A _11762_/B vssd1 vssd1 vccd1 vccd1 _11762_/X sky130_fd_sc_hd__and2_1
XTAP_2589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13501_ _13501_/A _13501_/B vssd1 vssd1 vccd1 vccd1 _13503_/A sky130_fd_sc_hd__nor2_1
XFILLER_158_105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10713_ _10713_/A _10713_/B vssd1 vssd1 vccd1 vccd1 _10715_/C sky130_fd_sc_hd__xnor2_1
XTAP_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14481_ _15457_/C _12864_/A _14733_/S vssd1 vssd1 vccd1 vccd1 _14481_/X sky130_fd_sc_hd__mux2_1
XTAP_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11693_ _11693_/A vssd1 vssd1 vccd1 vccd1 _11693_/Y sky130_fd_sc_hd__inv_2
XTAP_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16220_ _08776_/C _17075_/A2 _16218_/X _16219_/Y vssd1 vssd1 vccd1 vccd1 _16221_/A
+ sky130_fd_sc_hd__a211o_1
X_13432_ _13431_/A _13431_/B _13431_/C vssd1 vssd1 vccd1 vccd1 _13443_/B sky130_fd_sc_hd__o21ai_2
XFILLER_13_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10644_ _10644_/A _10649_/A _10644_/C vssd1 vssd1 vccd1 vccd1 _10653_/B sky130_fd_sc_hd__or3_1
XFILLER_13_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16151_ _16040_/B _16245_/A _16149_/X vssd1 vssd1 vccd1 vccd1 _16153_/A sky130_fd_sc_hd__a21oi_1
XFILLER_139_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13363_ _13363_/A _13363_/B vssd1 vssd1 vccd1 vccd1 _13364_/B sky130_fd_sc_hd__and2_1
X_10575_ _10567_/A _10572_/A _10573_/X _10574_/Y vssd1 vssd1 vccd1 vccd1 _10575_/Y
+ sky130_fd_sc_hd__o211ai_4
X_15102_ _15102_/A _15102_/B vssd1 vssd1 vccd1 vccd1 _15102_/Y sky130_fd_sc_hd__nand2_1
X_12314_ _12314_/A _12314_/B vssd1 vssd1 vccd1 vccd1 _12316_/C sky130_fd_sc_hd__nand2_1
XFILLER_155_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16082_ _15577_/Y _16361_/A _15954_/A vssd1 vssd1 vccd1 vccd1 _16082_/X sky130_fd_sc_hd__o21a_1
XFILLER_155_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13294_ _13295_/A _13295_/B _13295_/C vssd1 vssd1 vccd1 vccd1 _13308_/A sky130_fd_sc_hd__a21o_1
XFILLER_170_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15033_ _12025_/B _11813_/B _14765_/B _15033_/A3 _14942_/A _15095_/B vssd1 vssd1
+ vccd1 vccd1 _15034_/B sky130_fd_sc_hd__mux4_1
X_12245_ _13028_/A _12871_/B vssd1 vssd1 vccd1 vccd1 _12247_/B sky130_fd_sc_hd__nand2_1
XFILLER_5_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12176_ _17415_/A _12338_/C vssd1 vssd1 vccd1 vccd1 _12177_/B sky130_fd_sc_hd__nand2_1
XFILLER_68_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11127_ _11257_/A _11257_/B vssd1 vssd1 vccd1 vccd1 _11130_/C sky130_fd_sc_hd__nand2_1
X_16984_ _17083_/A _17040_/A _16984_/C vssd1 vssd1 vccd1 vccd1 _16986_/B sky130_fd_sc_hd__and3_1
XFILLER_122_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11058_ _11058_/A _11058_/B vssd1 vssd1 vccd1 vccd1 _11059_/C sky130_fd_sc_hd__xnor2_1
X_15935_ _15935_/A _15935_/B vssd1 vssd1 vccd1 vccd1 _15937_/B sky130_fd_sc_hd__xnor2_1
XFILLER_95_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10009_ _10009_/A _10009_/B _10009_/C vssd1 vssd1 vccd1 vccd1 _10010_/B sky130_fd_sc_hd__nand3_1
X_15866_ _15866_/A _15866_/B _15866_/C vssd1 vssd1 vccd1 vccd1 _15867_/B sky130_fd_sc_hd__or3_1
XFILLER_97_1036 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17605_ fanout934/X _17605_/D vssd1 vssd1 vccd1 vccd1 _17605_/Q sky130_fd_sc_hd__dfxtp_1
X_14817_ _14775_/X _14816_/X _12560_/A vssd1 vssd1 vccd1 vccd1 _16577_/A sky130_fd_sc_hd__a21bo_1
XFILLER_92_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15797_ _15797_/A _15797_/B vssd1 vssd1 vccd1 vccd1 _15797_/Y sky130_fd_sc_hd__nand2_1
X_17536_ fanout947/X _17536_/D vssd1 vssd1 vccd1 vccd1 _17536_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_91_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14748_ _14748_/A _14748_/B vssd1 vssd1 vccd1 vccd1 _14750_/B sky130_fd_sc_hd__or2_1
XFILLER_17_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17467_ fanout955/X _17467_/D vssd1 vssd1 vccd1 vccd1 _17467_/Q sky130_fd_sc_hd__dfxtp_1
X_14679_ _14649_/A _14679_/B vssd1 vssd1 vccd1 vccd1 _14680_/C sky130_fd_sc_hd__nand2b_1
XFILLER_20_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16418_ _16419_/A _16419_/B vssd1 vssd1 vccd1 vccd1 _16519_/B sky130_fd_sc_hd__or2_1
X_17398_ input44/X _17422_/A2 _17397_/X _17422_/C1 vssd1 vssd1 vccd1 vccd1 _17527_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_164_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16349_ _16266_/A _16266_/B _16267_/Y vssd1 vssd1 vccd1 vccd1 _16363_/B sky130_fd_sc_hd__a21bo_1
XFILLER_172_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout127 _17273_/A2 vssd1 vssd1 vccd1 vccd1 _17291_/A2 sky130_fd_sc_hd__buf_2
XFILLER_102_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout138 _15734_/B vssd1 vssd1 vccd1 vccd1 _16315_/C sky130_fd_sc_hd__clkbuf_4
Xfanout149 _14912_/Y vssd1 vssd1 vccd1 vccd1 _15097_/A sky130_fd_sc_hd__buf_2
X_09723_ _09723_/A _09723_/B vssd1 vssd1 vccd1 vccd1 _09725_/C sky130_fd_sc_hd__or2_1
XFILLER_74_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09654_ _09655_/A _09653_/Y _09654_/C _11808_/B vssd1 vssd1 vccd1 vccd1 _09784_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_103_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_24 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_876 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09585_ _09728_/B _12500_/B _11861_/B _09873_/A vssd1 vssd1 vccd1 vccd1 _09585_/Y
+ sky130_fd_sc_hd__a22oi_1
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_171 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_54 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10360_ _10591_/A _11027_/A _10479_/B _10594_/B vssd1 vssd1 vccd1 vccd1 _10374_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_164_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09019_ _08905_/A _08905_/C _08905_/B vssd1 vssd1 vccd1 vccd1 _09051_/B sky130_fd_sc_hd__a21o_1
XFILLER_136_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10291_ _14787_/A _10745_/D _10786_/B _14786_/A vssd1 vssd1 vccd1 vccd1 _10291_/Y
+ sky130_fd_sc_hd__a22oi_1
X_12030_ _12025_/A _09350_/B _14948_/B vssd1 vssd1 vccd1 vccd1 _12031_/B sky130_fd_sc_hd__a21o_1
XFILLER_105_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout650 _13908_/B vssd1 vssd1 vccd1 vccd1 _13735_/D sky130_fd_sc_hd__buf_2
Xfanout661 _16974_/A vssd1 vssd1 vccd1 vccd1 _14545_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_93_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout672 _11808_/B vssd1 vssd1 vccd1 vccd1 _12275_/D sky130_fd_sc_hd__clkbuf_4
Xfanout683 fanout690/X vssd1 vssd1 vccd1 vccd1 _13464_/B sky130_fd_sc_hd__buf_2
X_13981_ _13982_/A _13982_/B vssd1 vssd1 vccd1 vccd1 _14072_/A sky130_fd_sc_hd__and2b_1
XFILLER_77_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout694 fanout699/X vssd1 vssd1 vccd1 vccd1 _13691_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_59_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15720_ _11700_/Y _16106_/A _15701_/X _15719_/X vssd1 vssd1 vccd1 vccd1 _15720_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_101_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12932_ _13117_/B _12932_/B vssd1 vssd1 vccd1 vccd1 _12933_/C sky130_fd_sc_hd__nand2_1
XTAP_3021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15651_ _15651_/A _15651_/B vssd1 vssd1 vccd1 vccd1 _15742_/B sky130_fd_sc_hd__xnor2_1
XTAP_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12863_ _12861_/X _12862_/X _13840_/S vssd1 vssd1 vccd1 vccd1 _12864_/A sky130_fd_sc_hd__mux2_1
XTAP_3076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14602_ _14601_/A _14601_/B _14601_/C vssd1 vssd1 vccd1 vccd1 _14646_/A sky130_fd_sc_hd__o21ai_1
XTAP_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11814_ _14982_/B _14981_/B _11837_/A vssd1 vssd1 vccd1 vccd1 _11814_/Y sky130_fd_sc_hd__o21ai_1
XTAP_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15582_ _15582_/A _15582_/B vssd1 vssd1 vccd1 vccd1 _15584_/B sky130_fd_sc_hd__xnor2_1
X_12794_ _12794_/A _12794_/B vssd1 vssd1 vccd1 vccd1 _12796_/A sky130_fd_sc_hd__nor2_1
XTAP_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17321_ input39/X _17321_/B _17321_/C vssd1 vssd1 vccd1 vccd1 _17321_/X sky130_fd_sc_hd__or3_1
XTAP_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14533_ _14533_/A _14533_/B _14533_/C vssd1 vssd1 vccd1 vccd1 _14534_/B sky130_fd_sc_hd__and3_1
XTAP_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11745_ _11745_/A _11745_/B vssd1 vssd1 vccd1 vccd1 _11747_/B sky130_fd_sc_hd__xnor2_1
XFILLER_42_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17252_ _17593_/Q _17291_/A2 _17291_/B1 vssd1 vssd1 vccd1 vccd1 _17252_/X sky130_fd_sc_hd__a21o_1
X_14464_ _14463_/B _14463_/C _14463_/A vssd1 vssd1 vccd1 vccd1 _14465_/B sky130_fd_sc_hd__a21o_1
XFILLER_174_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11676_ _11676_/A _15011_/A vssd1 vssd1 vccd1 vccd1 _11679_/A sky130_fd_sc_hd__nor2_1
XFILLER_30_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16203_ _16203_/A _16203_/B _16099_/X vssd1 vssd1 vccd1 vccd1 _16203_/X sky130_fd_sc_hd__or3b_1
X_13415_ _13415_/A _13415_/B vssd1 vssd1 vccd1 vccd1 _13417_/C sky130_fd_sc_hd__nor2_1
X_10627_ _10713_/A _10713_/B vssd1 vssd1 vccd1 vccd1 _10627_/X sky130_fd_sc_hd__and2_1
X_17183_ input14/X input3/X vssd1 vssd1 vccd1 vccd1 _17428_/C sky130_fd_sc_hd__nor2_1
XFILLER_127_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14395_ _14396_/A _14396_/B vssd1 vssd1 vccd1 vccd1 _14395_/Y sky130_fd_sc_hd__nor2_1
XFILLER_10_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16134_ _16136_/A _16136_/B vssd1 vssd1 vccd1 vccd1 _16234_/C sky130_fd_sc_hd__nand2_1
XFILLER_127_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13346_ _13346_/A _13346_/B _13346_/C vssd1 vssd1 vccd1 vccd1 _13347_/B sky130_fd_sc_hd__and3_1
XFILLER_154_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10558_ _10560_/B _11027_/C _11027_/D _10560_/A vssd1 vssd1 vccd1 vccd1 _10561_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_170_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16065_ _16355_/A _16065_/B vssd1 vssd1 vccd1 vccd1 _16066_/B sky130_fd_sc_hd__nand2_1
X_13277_ _14757_/S _14735_/A1 _12218_/A _13276_/Y _14636_/A vssd1 vssd1 vccd1 vccd1
+ _13277_/X sky130_fd_sc_hd__a311o_1
XFILLER_170_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10489_ _10489_/A _10489_/B vssd1 vssd1 vccd1 vccd1 _10496_/A sky130_fd_sc_hd__xnor2_1
X_15016_ _16582_/A _15001_/X _15015_/X vssd1 vssd1 vccd1 vccd1 _15016_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_170_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12228_ _11824_/Y _11852_/B _12700_/B vssd1 vssd1 vccd1 vccd1 _12229_/C sky130_fd_sc_hd__mux2_1
XFILLER_123_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12159_ _17409_/A _12487_/D vssd1 vssd1 vccd1 vccd1 _12161_/C sky130_fd_sc_hd__nand2_1
XFILLER_1_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16967_ _16858_/Y _16914_/A _16914_/B vssd1 vssd1 vccd1 vccd1 _16967_/X sky130_fd_sc_hd__o21ba_1
XFILLER_37_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15918_ _15918_/A _16129_/A _16743_/C _17043_/B vssd1 vssd1 vccd1 vccd1 _15918_/X
+ sky130_fd_sc_hd__and4_1
X_16898_ _16897_/A _16897_/B _16897_/C vssd1 vssd1 vccd1 vccd1 _16900_/B sky130_fd_sc_hd__o21ai_1
XFILLER_65_854 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15849_ _16165_/A _16165_/B vssd1 vssd1 vccd1 vccd1 _15850_/B sky130_fd_sc_hd__nand2_1
XFILLER_80_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09370_ _09370_/A _09370_/B _09370_/C vssd1 vssd1 vccd1 vccd1 _09387_/B sky130_fd_sc_hd__nand3_1
XFILLER_80_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17519_ fanout942/X _17519_/D vssd1 vssd1 vccd1 vccd1 _17519_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_71_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_34 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09706_ _09706_/A _09706_/B vssd1 vssd1 vccd1 vccd1 _09709_/A sky130_fd_sc_hd__nor2_1
XFILLER_55_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwb_buttons_leds_968 vssd1 vssd1 vccd1 vccd1 wb_buttons_leds_968/HI led_enb[10] sky130_fd_sc_hd__conb_1
XFILLER_55_353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09637_ _09797_/A _14770_/A _10067_/B _10446_/B vssd1 vssd1 vccd1 vccd1 _09640_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_83_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09568_ _10255_/A _10897_/B vssd1 vssd1 vccd1 vccd1 _16989_/A sky130_fd_sc_hd__nand2_4
XFILLER_43_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09499_ _09620_/A _09500_/B vssd1 vssd1 vccd1 vccd1 _09499_/Y sky130_fd_sc_hd__nand2_1
XFILLER_24_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11530_ _11534_/B _11530_/B _11530_/C vssd1 vssd1 vccd1 vccd1 _11574_/A sky130_fd_sc_hd__and3_1
XFILLER_135_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11461_ _11460_/B _11461_/B vssd1 vssd1 vccd1 vccd1 _11703_/B sky130_fd_sc_hd__and2b_1
XFILLER_139_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13200_ _13369_/A _13200_/B vssd1 vssd1 vccd1 vccd1 _13202_/C sky130_fd_sc_hd__nor2_1
XFILLER_20_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10412_ _14786_/A _14787_/A _10786_/B _10743_/D vssd1 vssd1 vccd1 vccd1 _10415_/A
+ sky130_fd_sc_hd__and4_1
X_11392_ _11393_/B _11393_/C _11393_/A vssd1 vssd1 vccd1 vccd1 _11453_/A sky130_fd_sc_hd__o21ai_1
XFILLER_136_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14180_ _14180_/A _14180_/B vssd1 vssd1 vccd1 vccd1 _14181_/C sky130_fd_sc_hd__xnor2_1
XFILLER_87_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13131_ _12956_/A _12960_/A _13264_/A _13130_/Y vssd1 vssd1 vccd1 vccd1 _13264_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_109_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10343_ _10342_/A _10342_/B _10342_/C vssd1 vssd1 vccd1 vccd1 _10343_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_152_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13062_ _13061_/A _13061_/B _13061_/C vssd1 vssd1 vccd1 vccd1 _13063_/B sky130_fd_sc_hd__a21o_1
X_10274_ _10271_/A _10014_/D _10272_/X _10269_/X _10145_/B vssd1 vssd1 vccd1 vccd1
+ _10276_/B sky130_fd_sc_hd__a32o_1
XFILLER_105_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12013_ _12013_/A _12013_/B vssd1 vssd1 vccd1 vccd1 _12014_/B sky130_fd_sc_hd__and2_1
XFILLER_105_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16821_ _16822_/A _16822_/B vssd1 vssd1 vccd1 vccd1 _16897_/A sky130_fd_sc_hd__nor2_1
XFILLER_38_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout480 _17521_/Q vssd1 vssd1 vccd1 vccd1 _13182_/A sky130_fd_sc_hd__buf_2
XFILLER_94_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout491 _09728_/B vssd1 vssd1 vccd1 vccd1 _17383_/A sky130_fd_sc_hd__clkbuf_4
X_16752_ _16751_/A _16751_/B _16751_/C vssd1 vssd1 vccd1 vccd1 _16835_/A sky130_fd_sc_hd__a21oi_1
XFILLER_59_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13964_ _13964_/A _13964_/B vssd1 vssd1 vccd1 vccd1 _13971_/A sky130_fd_sc_hd__xnor2_1
XFILLER_93_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15703_ _15709_/A _16571_/B _15262_/A vssd1 vssd1 vccd1 vccd1 _15705_/B sky130_fd_sc_hd__or3b_1
X_12915_ _12915_/A _12915_/B _12915_/C vssd1 vssd1 vccd1 vccd1 _12916_/B sky130_fd_sc_hd__and3_1
XFILLER_46_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16683_ _16880_/A _16760_/B vssd1 vssd1 vccd1 vccd1 _16684_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13895_ _14318_/A _14318_/B _14426_/D _14360_/D vssd1 vssd1 vccd1 vccd1 _13896_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_94_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15634_ _16917_/A _15621_/Y _15633_/Y _15613_/Y vssd1 vssd1 vccd1 vccd1 _15634_/Y
+ sky130_fd_sc_hd__a211oi_1
XFILLER_64_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12846_ _12844_/X _12845_/X _13833_/S vssd1 vssd1 vccd1 vccd1 _12847_/B sky130_fd_sc_hd__mux2_1
XTAP_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15565_ _16317_/B _16533_/A _16695_/A _15647_/A vssd1 vssd1 vccd1 vccd1 _15568_/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12777_ _12778_/A _12778_/B _12778_/C vssd1 vssd1 vccd1 vccd1 _12779_/A sky130_fd_sc_hd__a21oi_1
XTAP_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17304_ _17304_/A1 _17322_/A2 _17303_/X _17358_/C1 vssd1 vssd1 vccd1 vccd1 _17481_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14516_ _14518_/A _14518_/B _14518_/C vssd1 vssd1 vccd1 vccd1 _14519_/B sky130_fd_sc_hd__a21o_1
X_11728_ _11725_/A _11725_/B _11725_/C vssd1 vssd1 vccd1 vccd1 _11729_/C sky130_fd_sc_hd__a21oi_1
XFILLER_30_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15496_ _15496_/A _15496_/B vssd1 vssd1 vccd1 vccd1 _15498_/A sky130_fd_sc_hd__nor2_1
XFILLER_147_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17235_ _17555_/Q _17274_/B vssd1 vssd1 vccd1 vccd1 _17235_/X sky130_fd_sc_hd__and2_1
XFILLER_174_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14447_ _14508_/A _14446_/C _14446_/A vssd1 vssd1 vccd1 vccd1 _14459_/B sky130_fd_sc_hd__a21o_1
XFILLER_80_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11659_ _11659_/A _11659_/B vssd1 vssd1 vccd1 vccd1 _11681_/B sky130_fd_sc_hd__xnor2_1
XFILLER_30_798 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17166_ _17166_/A _17166_/B _17166_/C vssd1 vssd1 vccd1 vccd1 _17166_/X sky130_fd_sc_hd__and3_1
XFILLER_7_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14378_ _14378_/A _14378_/B _14378_/C vssd1 vssd1 vccd1 vccd1 _14379_/B sky130_fd_sc_hd__and3_1
XFILLER_171_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16117_ _15715_/A _17164_/B _17164_/D _15628_/A vssd1 vssd1 vccd1 vccd1 _16117_/X
+ sky130_fd_sc_hd__o31a_1
X_13329_ _13329_/A _13329_/B _13329_/C vssd1 vssd1 vccd1 vccd1 _13330_/B sky130_fd_sc_hd__nand3_1
XFILLER_6_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17097_ _17096_/A _17096_/B _17096_/C vssd1 vssd1 vccd1 vccd1 _17097_/X sky130_fd_sc_hd__o21a_1
XFILLER_50_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16048_ _16048_/A _16048_/B vssd1 vssd1 vccd1 vccd1 _16051_/A sky130_fd_sc_hd__xnor2_1
XFILLER_143_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08870_ _08844_/X _08908_/A _08868_/X _08869_/Y vssd1 vssd1 vccd1 vccd1 _08873_/C
+ sky130_fd_sc_hd__o211ai_4
XFILLER_9_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09422_ _09423_/A _09423_/B vssd1 vssd1 vccd1 vccd1 _09441_/A sky130_fd_sc_hd__nand2b_1
XFILLER_53_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_665 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09353_ _09353_/A _09491_/A vssd1 vssd1 vccd1 vccd1 _09355_/B sky130_fd_sc_hd__nor2_1
XFILLER_40_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_570 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09284_ _13302_/A _12500_/B vssd1 vssd1 vccd1 vccd1 _09421_/A sky130_fd_sc_hd__and2_1
XFILLER_166_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08999_ _08999_/A _08999_/B vssd1 vssd1 vccd1 vccd1 _09001_/A sky130_fd_sc_hd__nor2_1
XFILLER_90_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_662 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10961_ _11010_/B _10961_/B _11043_/B vssd1 vssd1 vccd1 vccd1 _10978_/A sky130_fd_sc_hd__or3_1
XFILLER_44_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12700_ _12845_/S _12700_/B _12700_/C _14912_/B vssd1 vssd1 vccd1 vccd1 _13628_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_44_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13680_ _13680_/A _13680_/B _13680_/C vssd1 vssd1 vccd1 vccd1 _13681_/B sky130_fd_sc_hd__nor3_1
XFILLER_70_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10892_ _11148_/A _10892_/B vssd1 vssd1 vccd1 vccd1 _10893_/C sky130_fd_sc_hd__and2_1
X_12631_ _12631_/A _12631_/B _12631_/C vssd1 vssd1 vccd1 vccd1 _12631_/Y sky130_fd_sc_hd__nor3_2
XFILLER_169_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15350_ _15350_/A _15350_/B vssd1 vssd1 vccd1 vccd1 _15352_/B sky130_fd_sc_hd__xnor2_1
X_12562_ _12561_/A _12561_/B _12561_/C vssd1 vssd1 vccd1 vccd1 _12730_/A sky130_fd_sc_hd__o21ai_1
XFILLER_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14301_ _14680_/A _14599_/B _14301_/C _14485_/D vssd1 vssd1 vccd1 vccd1 _14302_/B
+ sky130_fd_sc_hd__and4_1
X_11513_ _11475_/A _11475_/C _11475_/B vssd1 vssd1 vccd1 vccd1 _11514_/C sky130_fd_sc_hd__a21oi_1
XFILLER_8_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15281_ _15281_/A _15281_/B vssd1 vssd1 vccd1 vccd1 _15283_/B sky130_fd_sc_hd__xnor2_1
XFILLER_11_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12493_ _12492_/A _12492_/B _12492_/C vssd1 vssd1 vccd1 vccd1 _12494_/B sky130_fd_sc_hd__o21a_1
X_17020_ _16966_/B _16969_/B _16966_/A vssd1 vssd1 vccd1 vccd1 _17066_/B sky130_fd_sc_hd__o21bai_1
XFILLER_7_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14232_ _14232_/A _14232_/B vssd1 vssd1 vccd1 vccd1 _14235_/A sky130_fd_sc_hd__xor2_1
X_11444_ _11444_/A _11444_/B _11444_/C vssd1 vssd1 vccd1 vccd1 _11444_/Y sky130_fd_sc_hd__nand3_2
XFILLER_7_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14163_ _14237_/A _14237_/B vssd1 vssd1 vccd1 vccd1 _14165_/B sky130_fd_sc_hd__xor2_1
X_11375_ _11553_/B _11518_/C _11325_/A _11324_/D vssd1 vssd1 vccd1 vccd1 _11376_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_164_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13114_ _13114_/A _13114_/B vssd1 vssd1 vccd1 vccd1 _13115_/B sky130_fd_sc_hd__nor2_1
XFILLER_152_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10326_ _10559_/A _10594_/B _10326_/C vssd1 vssd1 vccd1 vccd1 _10329_/B sky130_fd_sc_hd__nand3_1
XFILLER_113_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14094_ _14254_/A _14094_/B _14094_/C vssd1 vssd1 vccd1 vccd1 _14200_/B sky130_fd_sc_hd__and3_1
XFILLER_112_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13045_ _13046_/A _13046_/B _13046_/C vssd1 vssd1 vccd1 vccd1 _13047_/A sky130_fd_sc_hd__a21o_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10257_ _10257_/A _10257_/B vssd1 vssd1 vccd1 vccd1 _10372_/B sky130_fd_sc_hd__nor2_1
XFILLER_105_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10188_ _10188_/A _10188_/B _10188_/C vssd1 vssd1 vccd1 vccd1 _10188_/Y sky130_fd_sc_hd__nand3_1
XFILLER_67_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16804_ _17070_/B _16795_/Y _16797_/X _16007_/A _16803_/X vssd1 vssd1 vccd1 vccd1
+ _16804_/X sky130_fd_sc_hd__o221a_1
XFILLER_93_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14996_ _10255_/B _10270_/B _10142_/B _10014_/D _09925_/A _10182_/C vssd1 vssd1 vccd1
+ vccd1 _14998_/B sky130_fd_sc_hd__mux4_1
XFILLER_47_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13947_ _13948_/A _13948_/C vssd1 vssd1 vccd1 vccd1 _13947_/Y sky130_fd_sc_hd__nand2_1
XFILLER_46_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16735_ _16735_/A _16735_/B vssd1 vssd1 vccd1 vccd1 _16735_/Y sky130_fd_sc_hd__nor2_1
XFILLER_93_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16666_ _16667_/A _16938_/D vssd1 vssd1 vccd1 vccd1 _16670_/B sky130_fd_sc_hd__nor2_1
XFILLER_46_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13878_ _13878_/A _13878_/B vssd1 vssd1 vccd1 vccd1 _13880_/A sky130_fd_sc_hd__nor2_1
XFILLER_50_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15617_ _15617_/A _16571_/B _15262_/B vssd1 vssd1 vccd1 vccd1 _15618_/B sky130_fd_sc_hd__or3b_1
X_12829_ _12826_/A _12827_/Y _12676_/A _12677_/Y vssd1 vssd1 vccd1 vccd1 _12829_/Y
+ sky130_fd_sc_hd__a211oi_1
X_16597_ _16597_/A _16597_/B vssd1 vssd1 vccd1 vccd1 _16600_/A sky130_fd_sc_hd__xnor2_1
XFILLER_62_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15548_ _15548_/A vssd1 vssd1 vccd1 vccd1 _17552_/D sky130_fd_sc_hd__clkinv_2
XFILLER_148_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15479_ _15564_/A _15479_/B vssd1 vssd1 vccd1 vccd1 _15481_/B sky130_fd_sc_hd__nand2_1
X_17218_ _17440_/Q _17275_/A2 _17216_/X _17217_/X _17364_/C1 vssd1 vssd1 vccd1 vccd1
+ _17440_/D sky130_fd_sc_hd__o221a_1
XFILLER_163_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17149_ _17119_/B _17086_/A _17038_/C _16315_/A vssd1 vssd1 vccd1 vccd1 _17149_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_116_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09971_ _09964_/A _09962_/X _09923_/A _09957_/A vssd1 vssd1 vccd1 vccd1 _10091_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_115_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08922_ _08922_/A _08922_/B vssd1 vssd1 vccd1 vccd1 _08923_/B sky130_fd_sc_hd__nor2_1
XFILLER_130_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_851 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08853_ _17379_/A _11895_/B _11895_/D _11902_/B vssd1 vssd1 vccd1 vccd1 _08854_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_97_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08784_ _08791_/A _08791_/B _09058_/C _09446_/D vssd1 vssd1 vccd1 vccd1 _08798_/A
+ sky130_fd_sc_hd__and4_1
XTAP_2908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_963 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09405_ _17401_/A _09267_/D _09268_/A _09266_/Y vssd1 vssd1 vccd1 vccd1 _09411_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_164_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09336_ _09344_/A _09316_/X _09334_/A _09335_/Y vssd1 vssd1 vccd1 vccd1 _09339_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_139_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09267_ _09268_/A _09266_/Y _12070_/A _09267_/D vssd1 vssd1 vccd1 vccd1 _09411_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_138_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09198_ _12795_/A _09555_/C _09198_/C vssd1 vssd1 vccd1 vccd1 _09227_/B sky130_fd_sc_hd__nand3_1
XFILLER_101_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11160_ _11160_/A _11160_/B vssd1 vssd1 vccd1 vccd1 _11162_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10111_ _10112_/A _10110_/Y _10111_/C _10111_/D vssd1 vssd1 vccd1 vccd1 _10234_/A
+ sky130_fd_sc_hd__and4bb_1
X_11091_ _11080_/A _11080_/C _11080_/D _11080_/B vssd1 vssd1 vccd1 vccd1 _11145_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_121_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_916 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10042_ _10042_/A _10046_/A _10042_/C vssd1 vssd1 vccd1 vccd1 _10050_/B sky130_fd_sc_hd__or3_1
XFILLER_121_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_724 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14850_ _14850_/A _15314_/A _15314_/B vssd1 vssd1 vccd1 vccd1 _15463_/B sky130_fd_sc_hd__and3_1
XFILLER_152_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13801_ _13801_/A _13801_/B vssd1 vssd1 vccd1 vccd1 _13803_/A sky130_fd_sc_hd__nor2_1
XFILLER_35_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14781_ _16809_/A _15898_/A vssd1 vssd1 vccd1 vccd1 _15895_/B sky130_fd_sc_hd__or2_1
X_11993_ _11993_/A _12155_/B _11993_/C vssd1 vssd1 vccd1 vccd1 _12197_/A sky130_fd_sc_hd__nor3_1
XFILLER_29_695 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16520_ _16625_/A _16520_/B vssd1 vssd1 vccd1 vccd1 _16522_/B sky130_fd_sc_hd__nor2_1
XFILLER_17_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13732_ _13936_/A _13732_/B vssd1 vssd1 vccd1 vccd1 _13828_/B sky130_fd_sc_hd__or2_1
X_10944_ _10995_/B _10902_/B _10902_/C vssd1 vssd1 vccd1 vccd1 _10945_/B sky130_fd_sc_hd__o21ai_1
XFILLER_43_131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_676 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16451_ _16354_/B _16356_/B _16354_/A vssd1 vssd1 vccd1 vccd1 _16453_/B sky130_fd_sc_hd__o21ba_1
X_13663_ _14213_/B _13764_/D _13664_/D _13966_/A vssd1 vssd1 vccd1 vccd1 _13665_/A
+ sky130_fd_sc_hd__a22oi_1
X_10875_ _10933_/A _11122_/B _10875_/C _10962_/B vssd1 vssd1 vccd1 vccd1 _10878_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_71_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15402_ _15402_/A _15402_/B _16695_/A vssd1 vssd1 vccd1 vccd1 _15484_/A sky130_fd_sc_hd__and3_1
XFILLER_31_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12614_ _12611_/X _12612_/Y _12458_/A _12458_/Y vssd1 vssd1 vccd1 vccd1 _12631_/B
+ sky130_fd_sc_hd__o211a_1
X_16382_ _16382_/A _16382_/B vssd1 vssd1 vccd1 vccd1 _16562_/B sky130_fd_sc_hd__or2_1
X_13594_ _13595_/A _13595_/B vssd1 vssd1 vccd1 vccd1 _13594_/X sky130_fd_sc_hd__and2b_1
XFILLER_157_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_523 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15333_ _16226_/B _16536_/A _15334_/A vssd1 vssd1 vccd1 vccd1 _15408_/B sky130_fd_sc_hd__and3_1
XFILLER_129_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12545_ _12543_/X _12544_/X _13833_/S vssd1 vssd1 vccd1 vccd1 _12545_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15264_ _15143_/X _15262_/X _15305_/C vssd1 vssd1 vccd1 vccd1 _16446_/A sky130_fd_sc_hd__a21bo_4
XFILLER_172_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12476_ _12476_/A _12476_/B _12476_/C vssd1 vssd1 vccd1 vccd1 _12477_/B sky130_fd_sc_hd__and3_1
X_17003_ _17003_/A _17003_/B _17003_/C vssd1 vssd1 vccd1 vccd1 _17004_/B sky130_fd_sc_hd__nand3_1
X_14215_ _14215_/A _14360_/D vssd1 vssd1 vccd1 vccd1 _14216_/B sky130_fd_sc_hd__nand2_1
X_11427_ _11427_/A _11506_/B _11427_/C _15402_/A vssd1 vssd1 vccd1 vccd1 _11430_/A
+ sky130_fd_sc_hd__and4_1
XANTENNA_5 _17523_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15195_ _08743_/A _15171_/Y _15173_/Y _15194_/X vssd1 vssd1 vccd1 vccd1 _15195_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_153_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14146_ _14229_/B _14146_/B vssd1 vssd1 vccd1 vccd1 _14148_/B sky130_fd_sc_hd__nor2_1
X_11358_ _11359_/A _11359_/B vssd1 vssd1 vccd1 vccd1 _11416_/B sky130_fd_sc_hd__nor2_1
XFILLER_99_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10309_ _10753_/A _10309_/B _10309_/C vssd1 vssd1 vccd1 vccd1 _10312_/A sky130_fd_sc_hd__and3_1
X_14077_ _14077_/A _14077_/B vssd1 vssd1 vccd1 vccd1 _14078_/B sky130_fd_sc_hd__or2_1
X_11289_ _11348_/A _11253_/B _11351_/A vssd1 vssd1 vccd1 vccd1 _11295_/B sky130_fd_sc_hd__o21ai_1
X_13028_ _13028_/A _13632_/D vssd1 vssd1 vccd1 vccd1 _13029_/B sky130_fd_sc_hd__nand2_1
XFILLER_6_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_919 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14979_ _15096_/S _14979_/B vssd1 vssd1 vccd1 vccd1 _14979_/Y sky130_fd_sc_hd__nor2_1
XFILLER_63_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16718_ _16715_/Y _16717_/Y _16911_/A vssd1 vssd1 vccd1 vccd1 _16718_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_19_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_643 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_440 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16649_ _16649_/A _16649_/B _16649_/C vssd1 vssd1 vccd1 vccd1 _16649_/X sky130_fd_sc_hd__and3_1
XFILLER_34_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09121_ _09015_/X _09017_/Y _09119_/A _09119_/Y vssd1 vssd1 vccd1 vccd1 _09122_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_148_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09052_ _09052_/A _09052_/B vssd1 vssd1 vccd1 vccd1 _09053_/B sky130_fd_sc_hd__nor2_1
XFILLER_148_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_792 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09954_ _10078_/A _10078_/B _09936_/A vssd1 vssd1 vccd1 vccd1 _09956_/B sky130_fd_sc_hd__a21o_1
XFILLER_131_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08905_ _08905_/A _08905_/B _08905_/C vssd1 vssd1 vccd1 vccd1 _09051_/A sky130_fd_sc_hd__nand3_2
XFILLER_103_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_724 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09885_ _09885_/A _09885_/B _09885_/C vssd1 vssd1 vccd1 vccd1 _10029_/A sky130_fd_sc_hd__and3_1
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08836_ _08913_/A _09728_/B _09321_/D _09319_/C vssd1 vssd1 vccd1 vccd1 _08862_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_58_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08767_ _17401_/A _09030_/C _08754_/C _08754_/D vssd1 vssd1 vccd1 vccd1 _08768_/B
+ sky130_fd_sc_hd__a22oi_1
XFILLER_57_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_621 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_635 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10660_ _10660_/A _10757_/A vssd1 vssd1 vccd1 vccd1 _10669_/B sky130_fd_sc_hd__nor2_1
XFILLER_167_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09319_ _17379_/A _11895_/B _09319_/C _09319_/D vssd1 vssd1 vccd1 vccd1 _09328_/A
+ sky130_fd_sc_hd__and4_1
X_10591_ _10591_/A _11027_/A _11006_/C _11027_/C vssd1 vssd1 vccd1 vccd1 _10592_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_167_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12330_ _12498_/B _12330_/B vssd1 vssd1 vccd1 vccd1 _12333_/A sky130_fd_sc_hd__nand2_1
XFILLER_127_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12261_ _12261_/A _12261_/B vssd1 vssd1 vccd1 vccd1 _12263_/B sky130_fd_sc_hd__xnor2_1
XFILLER_147_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14000_ _14001_/A _14001_/B vssd1 vssd1 vccd1 vccd1 _14092_/A sky130_fd_sc_hd__nand2_1
XFILLER_141_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11212_ _11212_/A _11212_/B vssd1 vssd1 vccd1 vccd1 _11216_/A sky130_fd_sc_hd__xnor2_2
XFILLER_134_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_924 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12192_ _12192_/A _12192_/B vssd1 vssd1 vccd1 vccd1 _12193_/C sky130_fd_sc_hd__xnor2_1
X_11143_ _11144_/A _11146_/B _11143_/C _11143_/D vssd1 vssd1 vccd1 vccd1 _11237_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_150_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput75 _17468_/Q vssd1 vssd1 vccd1 vccd1 leds[2] sky130_fd_sc_hd__clkbuf_1
XFILLER_122_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput86 _17445_/Q vssd1 vssd1 vccd1 vccd1 o_wb_data[11] sky130_fd_sc_hd__clkbuf_1
Xoutput97 _17455_/Q vssd1 vssd1 vccd1 vccd1 o_wb_data[21] sky130_fd_sc_hd__clkbuf_1
X_11074_ _11074_/A _11074_/B vssd1 vssd1 vccd1 vccd1 _11075_/C sky130_fd_sc_hd__nand2_1
X_15951_ _16165_/A _16355_/B vssd1 vssd1 vccd1 vccd1 _15953_/B sky130_fd_sc_hd__nand2_1
XFILLER_89_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14902_ _17119_/A _16880_/A _16758_/A _15147_/A vssd1 vssd1 vccd1 vccd1 _14967_/D
+ sky130_fd_sc_hd__or4b_1
XFILLER_49_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10025_ _09865_/B _09975_/X _09991_/Y _10005_/X vssd1 vssd1 vccd1 vccd1 _10025_/Y
+ sky130_fd_sc_hd__a211oi_1
XFILLER_76_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15882_ _15883_/A _15883_/B _15881_/Y vssd1 vssd1 vccd1 vccd1 _15884_/A sky130_fd_sc_hd__o21bai_1
XFILLER_48_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14833_ _17476_/D _17477_/D vssd1 vssd1 vccd1 vccd1 _14933_/B sky130_fd_sc_hd__or2_2
XFILLER_64_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17552_ fanout937/X _17552_/D vssd1 vssd1 vccd1 vccd1 _17552_/Q sky130_fd_sc_hd__dfxtp_1
X_14764_ _14765_/A _14765_/B vssd1 vssd1 vccd1 vccd1 _14764_/Y sky130_fd_sc_hd__nor2_1
XFILLER_17_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11976_ _12804_/B _12174_/D _12129_/B _17419_/A vssd1 vssd1 vccd1 vccd1 _11978_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_147_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16503_ _16503_/A _16670_/A vssd1 vssd1 vccd1 vccd1 _16503_/Y sky130_fd_sc_hd__nand2_1
X_13715_ _13601_/A _13604_/A _13818_/A _13714_/Y vssd1 vssd1 vccd1 vccd1 _13818_/B
+ sky130_fd_sc_hd__o211ai_1
X_10927_ _11074_/A _10928_/B vssd1 vssd1 vccd1 vccd1 _10927_/X sky130_fd_sc_hd__or2_1
X_17483_ fanout948/X _17483_/D vssd1 vssd1 vccd1 vccd1 _17483_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14695_ _14723_/B _14695_/B vssd1 vssd1 vccd1 vccd1 _14699_/A sky130_fd_sc_hd__or2_1
XFILLER_71_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16434_ _16511_/B _16434_/B vssd1 vssd1 vccd1 vccd1 _16436_/B sky130_fd_sc_hd__or2_1
X_13646_ _13749_/A _13645_/B _13645_/C vssd1 vssd1 vccd1 vccd1 _13648_/B sky130_fd_sc_hd__a21o_1
XFILLER_72_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10858_ _10859_/B _10859_/C _10859_/A vssd1 vssd1 vccd1 vccd1 _10861_/A sky130_fd_sc_hd__a21o_1
XFILLER_72_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16365_ _16365_/A _16365_/B vssd1 vssd1 vccd1 vccd1 _16367_/B sky130_fd_sc_hd__or2_1
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13577_ _13577_/A _13577_/B vssd1 vssd1 vccd1 vccd1 _13579_/A sky130_fd_sc_hd__nor2_1
X_10789_ _10792_/A _10897_/B _10901_/A _10787_/Y vssd1 vssd1 vccd1 vccd1 _10796_/B
+ sky130_fd_sc_hd__o2bb2a_1
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15316_ _15314_/A _15713_/B1 _14929_/X _14801_/B vssd1 vssd1 vccd1 vccd1 _15316_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_118_718 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_364 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12528_ _12528_/A _12528_/B _12528_/C vssd1 vssd1 vccd1 vccd1 _12530_/A sky130_fd_sc_hd__nor3_1
X_16296_ _16389_/A _16296_/B vssd1 vssd1 vccd1 vccd1 _16296_/Y sky130_fd_sc_hd__nand2_1
XFILLER_9_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15247_ _15175_/B _15116_/B _15110_/B _14906_/B vssd1 vssd1 vccd1 vccd1 _15248_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_145_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12459_ _12267_/Y _12290_/X _12457_/X _12458_/Y vssd1 vssd1 vccd1 vccd1 _12481_/A
+ sky130_fd_sc_hd__o211ai_4
X_15178_ _15174_/Y _15175_/X _15176_/Y _15177_/Y _16111_/A vssd1 vssd1 vccd1 vccd1
+ _15178_/X sky130_fd_sc_hd__a311o_1
XFILLER_67_1044 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14129_ _15457_/A _14127_/X _14128_/X vssd1 vssd1 vccd1 vccd1 _14129_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_113_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout309 _14962_/A vssd1 vssd1 vccd1 vccd1 _15175_/A sky130_fd_sc_hd__buf_4
XFILLER_99_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09670_ _09530_/X _09541_/X _09668_/A _09668_/Y vssd1 vssd1 vccd1 vccd1 _09670_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_94_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_749 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09104_ _17423_/A _09172_/B _09502_/B _17425_/A vssd1 vssd1 vccd1 vccd1 _09106_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_164_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09035_ _09048_/B _09048_/C _09048_/A vssd1 vssd1 vccd1 vccd1 _09050_/A sky130_fd_sc_hd__a21o_1
XFILLER_163_367 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout810 _15624_/A vssd1 vssd1 vccd1 vccd1 _15617_/A sky130_fd_sc_hd__clkbuf_4
Xfanout821 _09265_/C vssd1 vssd1 vccd1 vccd1 _10971_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_131_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09937_ _10560_/B _09937_/B vssd1 vssd1 vccd1 vccd1 _09953_/A sky130_fd_sc_hd__nand2_1
Xfanout832 _17486_/Q vssd1 vssd1 vccd1 vccd1 _10920_/B sky130_fd_sc_hd__buf_4
Xfanout843 _12463_/D vssd1 vssd1 vccd1 vccd1 _09937_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_120_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout854 _09128_/B vssd1 vssd1 vccd1 vccd1 _10072_/B sky130_fd_sc_hd__clkbuf_4
Xfanout865 _09979_/C vssd1 vssd1 vccd1 vccd1 _10203_/B sky130_fd_sc_hd__buf_2
XFILLER_58_543 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout876 _17304_/A1 vssd1 vssd1 vccd1 vccd1 _09981_/D sky130_fd_sc_hd__buf_2
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09868_ _09868_/A _09868_/B vssd1 vssd1 vccd1 vccd1 _09870_/C sky130_fd_sc_hd__or2_1
Xfanout887 _15402_/A vssd1 vssd1 vccd1 vccd1 _11592_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_133_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout898 _11468_/D vssd1 vssd1 vccd1 vccd1 _11629_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08819_ _17387_/A _09319_/D _08798_/A _08786_/Y vssd1 vssd1 vccd1 vccd1 _08821_/C
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_58_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09799_ _09801_/B _09798_/Y _10321_/A _10067_/B vssd1 vssd1 vccd1 vccd1 _09941_/A
+ sky130_fd_sc_hd__and4bb_1
XTAP_3247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11830_ _12923_/D _12770_/D _12050_/S vssd1 vssd1 vccd1 vccd1 _11831_/B sky130_fd_sc_hd__mux2_1
XTAP_2524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11761_ _11756_/A _11755_/B _11759_/A vssd1 vssd1 vccd1 vccd1 _11762_/B sky130_fd_sc_hd__a21o_1
XFILLER_60_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13500_ _13500_/A _13500_/B _13500_/C vssd1 vssd1 vccd1 vccd1 _13501_/B sky130_fd_sc_hd__nor3_1
XTAP_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10712_ _10729_/A _10729_/B vssd1 vssd1 vccd1 vccd1 _10712_/X sky130_fd_sc_hd__or2_1
XFILLER_14_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_668 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14480_ _14763_/S _14478_/X _14479_/Y _14423_/Y vssd1 vssd1 vccd1 vccd1 _17598_/D
+ sky130_fd_sc_hd__a31o_1
XTAP_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11692_ _15524_/C _11692_/B _11670_/C vssd1 vssd1 vccd1 vccd1 _11693_/A sky130_fd_sc_hd__or3b_1
XTAP_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13431_ _13431_/A _13431_/B _13431_/C vssd1 vssd1 vccd1 vccd1 _13443_/A sky130_fd_sc_hd__or3_1
X_10643_ _10644_/A _10644_/C vssd1 vssd1 vccd1 vccd1 _10649_/B sky130_fd_sc_hd__nor2_1
XFILLER_42_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16150_ _16667_/A _16827_/B vssd1 vssd1 vccd1 vccd1 _16245_/A sky130_fd_sc_hd__nor2_1
XFILLER_167_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13362_ _13363_/A _13363_/B vssd1 vssd1 vccd1 vccd1 _13482_/A sky130_fd_sc_hd__nor2_1
XFILLER_42_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10574_ _10458_/X _10472_/Y _10557_/X _10572_/X vssd1 vssd1 vccd1 vccd1 _10574_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_158_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15101_ _10657_/B _10308_/B _10431_/B _14863_/B _14914_/S _14958_/A vssd1 vssd1 vccd1
+ vccd1 _15102_/B sky130_fd_sc_hd__mux4_1
XFILLER_158_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12313_ _12312_/A _12312_/B _12312_/C vssd1 vssd1 vccd1 vccd1 _12314_/B sky130_fd_sc_hd__a21o_1
XFILLER_158_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16081_ _16081_/A _16081_/B vssd1 vssd1 vccd1 vccd1 _16089_/A sky130_fd_sc_hd__nand2_1
X_13293_ _13411_/B _13293_/B vssd1 vssd1 vccd1 vccd1 _13295_/C sky130_fd_sc_hd__nand2_1
XFILLER_170_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15032_ _12700_/C _12032_/Y _15100_/A _14948_/A vssd1 vssd1 vccd1 vccd1 _16011_/C
+ sky130_fd_sc_hd__o211ai_4
X_12244_ _12244_/A _12429_/A vssd1 vssd1 vccd1 vccd1 _12247_/A sky130_fd_sc_hd__or2_1
XFILLER_142_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_62 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12175_ _12175_/A _12175_/B vssd1 vssd1 vccd1 vccd1 _12177_/A sky130_fd_sc_hd__nor2_1
XFILLER_122_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11126_ _11126_/A _11126_/B vssd1 vssd1 vccd1 vccd1 _11257_/B sky130_fd_sc_hd__xnor2_1
XFILLER_1_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16983_ _16983_/A _17038_/B vssd1 vssd1 vccd1 vccd1 _16984_/C sky130_fd_sc_hd__nand2_1
XFILLER_3_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11057_ _11057_/A _11057_/B _11057_/C vssd1 vssd1 vccd1 vccd1 _11059_/B sky130_fd_sc_hd__nand3_1
X_15934_ _16416_/A _16041_/B vssd1 vssd1 vccd1 vccd1 _15935_/B sky130_fd_sc_hd__nor2_1
XFILLER_110_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_82 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10008_ _10009_/A _10009_/B _10009_/C vssd1 vssd1 vccd1 vccd1 _10010_/A sky130_fd_sc_hd__a21o_1
X_15865_ _15866_/A _15866_/B _15866_/C vssd1 vssd1 vccd1 vccd1 _15867_/A sky130_fd_sc_hd__o21ai_1
XFILLER_36_226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17604_ fanout936/X _17604_/D vssd1 vssd1 vccd1 vccd1 _17604_/Q sky130_fd_sc_hd__dfxtp_1
X_14816_ _16397_/B _16398_/A _12235_/C vssd1 vssd1 vccd1 vccd1 _14816_/X sky130_fd_sc_hd__a21o_1
X_15796_ _15811_/A _16571_/B _16136_/A vssd1 vssd1 vccd1 vccd1 _15797_/B sky130_fd_sc_hd__or3b_1
X_17535_ fanout944/X _17535_/D vssd1 vssd1 vccd1 vccd1 _17535_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_44_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11959_ _11958_/A _11958_/B _11958_/C vssd1 vssd1 vccd1 vccd1 _12169_/A sky130_fd_sc_hd__o21ai_1
X_14747_ _14747_/A _14747_/B _14747_/C vssd1 vssd1 vccd1 vccd1 _14748_/B sky130_fd_sc_hd__and3_1
XFILLER_32_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17466_ fanout955/X _17466_/D vssd1 vssd1 vccd1 vccd1 _17466_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14678_ _14678_/A _14678_/B vssd1 vssd1 vccd1 vccd1 _14682_/A sky130_fd_sc_hd__nor2_1
X_16417_ _16417_/A _16519_/A vssd1 vssd1 vccd1 vccd1 _16419_/B sky130_fd_sc_hd__nand2_1
X_13629_ _14210_/B _13627_/X _13628_/Y _15457_/B _14482_/B1 vssd1 vssd1 vccd1 vccd1
+ _13629_/X sky130_fd_sc_hd__o221a_1
XFILLER_34_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17397_ _17397_/A _17421_/B vssd1 vssd1 vccd1 vccd1 _17397_/X sky130_fd_sc_hd__or2_1
XFILLER_146_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16348_ _16462_/A _16348_/B vssd1 vssd1 vccd1 vccd1 _16367_/A sky130_fd_sc_hd__nand2b_1
XFILLER_118_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16279_ _16279_/A _16279_/B _16279_/C vssd1 vssd1 vccd1 vccd1 _16280_/B sky130_fd_sc_hd__nor3_1
XFILLER_145_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout128 _17273_/A2 vssd1 vssd1 vccd1 vccd1 _17282_/A2 sky130_fd_sc_hd__clkbuf_2
Xfanout139 _15074_/B vssd1 vssd1 vccd1 vccd1 _16226_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_86_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09722_ _09722_/A _09722_/B vssd1 vssd1 vccd1 vccd1 _09723_/B sky130_fd_sc_hd__nor2_1
XFILLER_55_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09653_ _15254_/S _09926_/B _14982_/B vssd1 vssd1 vccd1 vccd1 _09653_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_27_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09584_ _09873_/A _09728_/B _12500_/B _11861_/B vssd1 vssd1 vccd1 vccd1 _09587_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_55_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09018_ _08930_/A _08930_/C _08930_/B vssd1 vssd1 vccd1 vccd1 _09018_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_88_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10290_ _14786_/A _14787_/A _10745_/D _10743_/C vssd1 vssd1 vccd1 vccd1 _10293_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_145_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout640 _17507_/Q vssd1 vssd1 vccd1 vccd1 _15033_/A3 sky130_fd_sc_hd__buf_4
XFILLER_120_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout651 _17505_/Q vssd1 vssd1 vccd1 vccd1 _13908_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_59_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout662 _17504_/Q vssd1 vssd1 vccd1 vccd1 _16974_/A sky130_fd_sc_hd__clkbuf_4
X_13980_ _13980_/A _13980_/B vssd1 vssd1 vccd1 vccd1 _13982_/B sky130_fd_sc_hd__xnor2_1
XFILLER_19_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout673 _17503_/Q vssd1 vssd1 vccd1 vccd1 _11808_/B sky130_fd_sc_hd__buf_4
XFILLER_58_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout684 _16789_/A vssd1 vssd1 vccd1 vccd1 _14360_/D sky130_fd_sc_hd__clkbuf_4
Xfanout695 _12256_/D vssd1 vssd1 vccd1 vccd1 _09321_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_58_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12931_ _12931_/A _12931_/B vssd1 vssd1 vccd1 vccd1 _12932_/B sky130_fd_sc_hd__or2_1
XFILLER_46_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15650_ _15651_/A _15651_/B vssd1 vssd1 vccd1 vccd1 _15762_/A sky130_fd_sc_hd__and2_1
XFILLER_18_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12862_ _12386_/X _12389_/X _12865_/S vssd1 vssd1 vccd1 vccd1 _12862_/X sky130_fd_sc_hd__mux2_1
XTAP_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11813_ _12025_/A _11813_/B vssd1 vssd1 vccd1 vccd1 _14981_/B sky130_fd_sc_hd__and2_1
X_14601_ _14601_/A _14601_/B _14601_/C vssd1 vssd1 vccd1 vccd1 _14603_/A sky130_fd_sc_hd__or3_1
XTAP_3099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15581_ _15750_/A _16589_/B vssd1 vssd1 vccd1 vccd1 _15582_/B sky130_fd_sc_hd__nand2_1
X_12793_ _12792_/A _12792_/B _12792_/C vssd1 vssd1 vccd1 vccd1 _12794_/B sky130_fd_sc_hd__o21a_1
XTAP_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17320_ _09272_/D _17322_/A2 _17319_/X _17426_/C1 vssd1 vssd1 vccd1 vccd1 _17489_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14532_ _14585_/A _14532_/B vssd1 vssd1 vccd1 vccd1 _14629_/A sky130_fd_sc_hd__and2_1
XTAP_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11744_ _11745_/A _11745_/B vssd1 vssd1 vccd1 vccd1 _11750_/A sky130_fd_sc_hd__nand2b_1
XFILLER_15_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_947 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14463_ _14463_/A _14463_/B _14463_/C vssd1 vssd1 vccd1 vccd1 _14465_/A sky130_fd_sc_hd__nand3_1
X_17251_ _17451_/Q _17290_/A2 _17249_/X _17250_/X _17284_/C1 vssd1 vssd1 vccd1 vccd1
+ _17451_/D sky130_fd_sc_hd__o221a_1
X_11675_ _15056_/A _11675_/B _11675_/C vssd1 vssd1 vccd1 vccd1 _15011_/A sky130_fd_sc_hd__or3_1
XFILLER_174_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13414_ _13658_/A _13414_/B _13852_/B _13844_/C vssd1 vssd1 vccd1 vccd1 _13415_/B
+ sky130_fd_sc_hd__and4_1
X_16202_ _16098_/A _16101_/Y _16203_/B vssd1 vssd1 vccd1 vccd1 _16292_/B sky130_fd_sc_hd__a21oi_2
X_10626_ _10626_/A _10626_/B vssd1 vssd1 vccd1 vccd1 _10713_/B sky130_fd_sc_hd__nor2_1
X_17182_ input29/X wire215/X vssd1 vssd1 vccd1 vccd1 _17198_/C sky130_fd_sc_hd__and2b_1
XFILLER_168_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14394_ _14394_/A _14394_/B vssd1 vssd1 vccd1 vccd1 _14396_/B sky130_fd_sc_hd__or2_1
X_16133_ _16133_/A _16133_/B vssd1 vssd1 vccd1 vccd1 _16142_/A sky130_fd_sc_hd__xnor2_1
XFILLER_128_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13345_ _13346_/A _13346_/B _13346_/C vssd1 vssd1 vccd1 vccd1 _13347_/A sky130_fd_sc_hd__a21oi_1
XFILLER_154_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10557_ _10571_/A _10571_/B vssd1 vssd1 vccd1 vccd1 _10557_/X sky130_fd_sc_hd__or2_1
XFILLER_128_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16064_ _16064_/A _16064_/B vssd1 vssd1 vccd1 vccd1 _16066_/A sky130_fd_sc_hd__nor2_1
XFILLER_6_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13276_ _14757_/S _13276_/B vssd1 vssd1 vccd1 vccd1 _13276_/Y sky130_fd_sc_hd__nor2_1
XFILLER_154_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10488_ _10489_/A _10489_/B vssd1 vssd1 vccd1 vccd1 _10503_/A sky130_fd_sc_hd__nand2b_1
XFILLER_154_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15015_ _15628_/A _17143_/A1 _11854_/X _15013_/Y vssd1 vssd1 vccd1 vccd1 _15015_/X
+ sky130_fd_sc_hd__o31a_1
X_12227_ _12219_/X _12226_/X _14356_/S vssd1 vssd1 vccd1 vccd1 _12227_/X sky130_fd_sc_hd__mux2_1
XFILLER_97_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_104 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12158_ _17413_/A _12787_/B _12320_/D _12158_/D vssd1 vssd1 vccd1 vccd1 _12325_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_2_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11109_ _11075_/A _11075_/B _11075_/C vssd1 vssd1 vccd1 vccd1 _11110_/C sky130_fd_sc_hd__o21ai_1
XFILLER_68_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12089_ _12089_/A _12089_/B vssd1 vssd1 vccd1 vccd1 _12091_/A sky130_fd_sc_hd__nor2_1
X_16966_ _16966_/A _16966_/B vssd1 vssd1 vccd1 vccd1 _16969_/A sky130_fd_sc_hd__or2_1
XFILLER_77_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15917_ _16129_/A _17043_/B vssd1 vssd1 vccd1 vccd1 _15917_/Y sky130_fd_sc_hd__nand2_1
X_16897_ _16897_/A _16897_/B _16897_/C vssd1 vssd1 vccd1 vccd1 _16900_/A sky130_fd_sc_hd__or3_1
XFILLER_37_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15848_ _15848_/A _15848_/B vssd1 vssd1 vccd1 vccd1 _15850_/A sky130_fd_sc_hd__nor2_1
XFILLER_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15779_ _15690_/A _15779_/B vssd1 vssd1 vccd1 vccd1 _15781_/B sky130_fd_sc_hd__nand2b_1
XFILLER_17_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17518_ fanout942/X _17518_/D vssd1 vssd1 vccd1 vccd1 _17518_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_33_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17449_ fanout954/X _17449_/D vssd1 vssd1 vccd1 vccd1 _17449_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09705_ _09718_/B _09718_/C _09718_/A vssd1 vssd1 vccd1 vccd1 _09720_/A sky130_fd_sc_hd__a21o_1
XFILLER_114_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwb_buttons_leds_958 vssd1 vssd1 vccd1 vccd1 wb_buttons_leds_958/HI led_enb[0] sky130_fd_sc_hd__conb_1
X_09636_ _09636_/A _09636_/B vssd1 vssd1 vccd1 vccd1 _09642_/A sky130_fd_sc_hd__nor2_1
Xwb_buttons_leds_969 vssd1 vssd1 vccd1 vccd1 wb_buttons_leds_969/HI led_enb[11] sky130_fd_sc_hd__conb_1
XFILLER_43_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_398 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09567_ _16933_/A _16982_/B vssd1 vssd1 vccd1 vccd1 _09567_/Y sky130_fd_sc_hd__nor2_1
XFILLER_130_67 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09498_ _09498_/A _09498_/B vssd1 vssd1 vccd1 vccd1 _09500_/B sky130_fd_sc_hd__or2_1
XFILLER_90_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11460_ _11460_/A _11460_/B _11460_/C vssd1 vssd1 vccd1 vccd1 _11461_/B sky130_fd_sc_hd__or3_2
XFILLER_128_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10411_ _10411_/A _10411_/B vssd1 vssd1 vccd1 vccd1 _10427_/A sky130_fd_sc_hd__xnor2_1
XFILLER_139_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11391_ _11520_/C _14895_/B _11436_/B vssd1 vssd1 vccd1 vccd1 _11393_/C sky130_fd_sc_hd__and3_1
XFILLER_87_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_827 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13130_ _13127_/X _13128_/Y _12987_/X _12993_/A vssd1 vssd1 vccd1 vccd1 _13130_/Y
+ sky130_fd_sc_hd__a211oi_1
X_10342_ _10342_/A _10342_/B _10342_/C vssd1 vssd1 vccd1 vccd1 _10345_/A sky130_fd_sc_hd__and3_1
XFILLER_136_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13061_ _13061_/A _13061_/B _13061_/C vssd1 vssd1 vccd1 vccd1 _13063_/A sky130_fd_sc_hd__nand3_1
XFILLER_3_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10273_ _15707_/A _15622_/A _10272_/X vssd1 vssd1 vccd1 vccd1 _10391_/B sky130_fd_sc_hd__o21a_1
X_12012_ _12013_/A _12013_/B vssd1 vssd1 vccd1 vccd1 _12375_/A sky130_fd_sc_hd__nor2_1
XFILLER_78_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16820_ _16750_/A _16750_/B _16883_/C _16670_/C vssd1 vssd1 vccd1 vccd1 _16822_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_93_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout470 _11790_/A vssd1 vssd1 vccd1 vccd1 _10126_/B sky130_fd_sc_hd__buf_4
XFILLER_19_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout481 _17521_/Q vssd1 vssd1 vccd1 vccd1 _12275_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_59_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16751_ _16751_/A _16751_/B _16751_/C vssd1 vssd1 vccd1 vccd1 _16753_/A sky130_fd_sc_hd__and3_1
XFILLER_19_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout492 _09299_/B vssd1 vssd1 vccd1 vccd1 _09728_/B sky130_fd_sc_hd__buf_4
XFILLER_93_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13963_ _13964_/A _13964_/B vssd1 vssd1 vccd1 vccd1 _14058_/A sky130_fd_sc_hd__nand2b_1
XFILLER_93_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_332 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15702_ _15262_/A _16644_/B _15206_/A vssd1 vssd1 vccd1 vccd1 _15705_/A sky130_fd_sc_hd__a21o_1
X_12914_ _12915_/A _12915_/B _12915_/C vssd1 vssd1 vccd1 vccd1 _13072_/B sky130_fd_sc_hd__a21oi_1
X_16682_ _16680_/X _16682_/B vssd1 vssd1 vccd1 vccd1 _16684_/A sky130_fd_sc_hd__nand2b_1
X_13894_ _14318_/A _14360_/D _16864_/A vssd1 vssd1 vccd1 vccd1 _13896_/A sky130_fd_sc_hd__a21boi_1
XFILLER_46_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12845_ _12211_/X _12224_/X _12845_/S vssd1 vssd1 vccd1 vccd1 _12845_/X sky130_fd_sc_hd__mux2_1
XTAP_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15633_ _15456_/B _15623_/X _15632_/X vssd1 vssd1 vccd1 vccd1 _15633_/Y sky130_fd_sc_hd__o21ai_1
XTAP_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12776_ _12931_/A _12776_/B vssd1 vssd1 vccd1 vccd1 _12778_/C sky130_fd_sc_hd__or2_1
XFILLER_15_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15564_ _15564_/A _15564_/B vssd1 vssd1 vccd1 vccd1 _15588_/A sky130_fd_sc_hd__xor2_1
XTAP_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17303_ input61/X _17321_/B _17321_/C vssd1 vssd1 vccd1 vccd1 _17303_/X sky130_fd_sc_hd__or3_1
XTAP_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11727_ _11732_/A _11727_/B vssd1 vssd1 vccd1 vccd1 _11729_/B sky130_fd_sc_hd__nand2_1
X_14515_ _14569_/B _14515_/B vssd1 vssd1 vccd1 vccd1 _14518_/C sky130_fd_sc_hd__nand2_1
XFILLER_148_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15495_ _16056_/A _16589_/B _15213_/C vssd1 vssd1 vccd1 vccd1 _15496_/B sky130_fd_sc_hd__a21oi_1
XFILLER_30_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17234_ _17587_/Q _17273_/A2 _17273_/B1 vssd1 vssd1 vccd1 vccd1 _17234_/X sky130_fd_sc_hd__a21o_1
X_11658_ _15715_/A _15008_/B _11681_/A _11658_/D vssd1 vssd1 vccd1 vccd1 _11678_/A
+ sky130_fd_sc_hd__nand4_1
X_14446_ _14446_/A _14508_/A _14446_/C vssd1 vssd1 vccd1 vccd1 _14518_/A sky130_fd_sc_hd__nand3_1
X_10609_ _10610_/B _10610_/A vssd1 vssd1 vccd1 vccd1 _10615_/B sky130_fd_sc_hd__nand2b_1
XFILLER_128_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14377_ _14378_/A _14378_/B _14378_/C vssd1 vssd1 vccd1 vccd1 _14446_/A sky130_fd_sc_hd__a21oi_1
X_17165_ _16735_/A _14758_/B _17163_/X _17164_/X vssd1 vssd1 vccd1 vccd1 _17166_/C
+ sky130_fd_sc_hd__o211a_1
X_11589_ _11630_/A _11563_/D _11564_/A _11562_/Y vssd1 vssd1 vccd1 vccd1 _11590_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_116_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_602 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13328_ _13329_/A _13329_/B _13329_/C vssd1 vssd1 vccd1 vccd1 _13330_/A sky130_fd_sc_hd__a21o_1
X_16116_ _15097_/X _15100_/Y _15102_/Y _15123_/Y _15312_/S _15116_/A vssd1 vssd1 vccd1
+ vccd1 _16116_/X sky130_fd_sc_hd__mux4_1
XFILLER_115_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17096_ _17096_/A _17096_/B _17096_/C vssd1 vssd1 vccd1 vccd1 _17096_/Y sky130_fd_sc_hd__nor3_1
XFILLER_115_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16047_ _16048_/A _16048_/B vssd1 vssd1 vccd1 vccd1 _16047_/X sky130_fd_sc_hd__and2b_1
X_13259_ _13093_/B _13095_/B _13093_/A vssd1 vssd1 vccd1 vccd1 _13260_/A sky130_fd_sc_hd__o21ba_1
XFILLER_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16949_ _16950_/B _16950_/A vssd1 vssd1 vccd1 vccd1 _17003_/B sky130_fd_sc_hd__nand2b_1
XFILLER_65_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_983 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09421_ _09421_/A _09421_/B vssd1 vssd1 vccd1 vccd1 _09423_/B sky130_fd_sc_hd__xnor2_1
XFILLER_80_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09352_ _09353_/A _09351_/Y _14982_/A _11813_/B vssd1 vssd1 vccd1 vccd1 _09491_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_80_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09283_ _11006_/A _10897_/B vssd1 vssd1 vccd1 vccd1 _17119_/B sky130_fd_sc_hd__nand2_4
XFILLER_60_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_871 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08998_ _17373_/A _11930_/B _12439_/D _12447_/B vssd1 vssd1 vccd1 vccd1 _08999_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_75_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_950 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10960_ _10907_/B _10909_/B _10907_/A vssd1 vssd1 vccd1 vccd1 _11043_/B sky130_fd_sc_hd__o21ba_1
XFILLER_44_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09619_ _09619_/A _09619_/B _09656_/A vssd1 vssd1 vccd1 vccd1 _09620_/B sky130_fd_sc_hd__or3_1
X_10891_ _10891_/A _10891_/B _10891_/C vssd1 vssd1 vccd1 vccd1 _10892_/B sky130_fd_sc_hd__or3_1
XFILLER_16_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12630_ _12631_/A _12631_/B _12631_/C vssd1 vssd1 vccd1 vccd1 _12630_/X sky130_fd_sc_hd__o21a_1
XFILLER_43_357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_891 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12561_ _12561_/A _12561_/B _12561_/C vssd1 vssd1 vccd1 vccd1 _12563_/A sky130_fd_sc_hd__or3_1
XFILLER_54_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_587 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11512_ _11512_/A _11512_/B _11512_/C vssd1 vssd1 vccd1 vccd1 _11558_/A sky130_fd_sc_hd__nand3_2
XFILLER_129_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14300_ _14680_/A _14545_/D vssd1 vssd1 vccd1 vccd1 _14367_/A sky130_fd_sc_hd__nand2_1
XFILLER_156_215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15280_ _15281_/A _15281_/B vssd1 vssd1 vccd1 vccd1 _15428_/A sky130_fd_sc_hd__nor2_1
X_12492_ _12492_/A _12492_/B _12492_/C vssd1 vssd1 vccd1 vccd1 _12494_/A sky130_fd_sc_hd__nor3_1
XFILLER_8_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14231_ _14154_/A _14156_/B _14154_/B vssd1 vssd1 vccd1 vccd1 _14232_/B sky130_fd_sc_hd__o21ba_1
X_11443_ _11435_/A _11435_/B _11435_/C vssd1 vssd1 vccd1 vccd1 _11444_/C sky130_fd_sc_hd__a21o_1
XFILLER_171_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14162_ _14162_/A _14162_/B vssd1 vssd1 vccd1 vccd1 _14237_/B sky130_fd_sc_hd__nor2_1
XFILLER_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11374_ _11423_/B _11592_/B _11373_/B _11370_/X vssd1 vssd1 vccd1 vccd1 _11376_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_152_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13113_ _13114_/A _13114_/B vssd1 vssd1 vccd1 vccd1 _13248_/B sky130_fd_sc_hd__and2_1
XFILLER_153_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10325_ _10325_/A _10325_/B vssd1 vssd1 vccd1 vccd1 _10326_/C sky130_fd_sc_hd__and2_1
X_14093_ _14200_/A _14093_/B vssd1 vssd1 vccd1 vccd1 _14094_/C sky130_fd_sc_hd__nor2_1
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13044_ _13181_/B _13044_/B vssd1 vssd1 vccd1 vccd1 _13046_/C sky130_fd_sc_hd__and2_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10256_ _10126_/B _10920_/B _10799_/B _10254_/A vssd1 vssd1 vccd1 vccd1 _10257_/B
+ sky130_fd_sc_hd__a22oi_1
XFILLER_121_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_8 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10187_ _10188_/A _10188_/B _10188_/C vssd1 vssd1 vccd1 vccd1 _10187_/X sky130_fd_sc_hd__and3_1
XFILLER_67_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16803_ _17140_/A _14864_/B _16798_/Y _16802_/X vssd1 vssd1 vccd1 vccd1 _16803_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_94_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14995_ _14992_/Y _14994_/Y _15103_/S vssd1 vssd1 vccd1 vccd1 _14995_/X sky130_fd_sc_hd__mux2_1
XFILLER_19_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16734_ _13459_/A _17075_/A2 _16733_/X vssd1 vssd1 vccd1 vccd1 _16734_/X sky130_fd_sc_hd__a21o_1
X_13946_ _13948_/B _13948_/C _14094_/B _13948_/A vssd1 vssd1 vccd1 vccd1 _13949_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_62_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16665_ _16665_/A _16665_/B vssd1 vssd1 vccd1 vccd1 _16673_/A sky130_fd_sc_hd__xor2_1
XFILLER_61_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13877_ _13977_/A _13977_/B _14213_/D _14141_/D vssd1 vssd1 vccd1 vccd1 _13878_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_61_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15616_ _15262_/B _16209_/B _15617_/A vssd1 vssd1 vccd1 vccd1 _15616_/Y sky130_fd_sc_hd__a21boi_1
X_12828_ _12676_/A _12677_/Y _12826_/A _12827_/Y vssd1 vssd1 vccd1 vccd1 _12991_/A
+ sky130_fd_sc_hd__o211a_1
X_16596_ _16748_/C _16596_/B vssd1 vssd1 vccd1 vccd1 _16597_/B sky130_fd_sc_hd__xnor2_1
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15547_ _15541_/A _16806_/A2 _15523_/X _15546_/X vssd1 vssd1 vccd1 vccd1 _15548_/A
+ sky130_fd_sc_hd__a22o_1
X_12759_ _12759_/A _12759_/B vssd1 vssd1 vccd1 vccd1 _12761_/C sky130_fd_sc_hd__xnor2_1
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_930 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15478_ _16226_/C _16505_/A _15473_/X _15476_/Y vssd1 vssd1 vccd1 vccd1 _15479_/B
+ sky130_fd_sc_hd__a22o_1
X_17217_ _17549_/Q _17274_/B vssd1 vssd1 vccd1 vccd1 _17217_/X sky130_fd_sc_hd__and2_1
XFILLER_163_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14429_ _14430_/A _14430_/B vssd1 vssd1 vccd1 vccd1 _14497_/B sky130_fd_sc_hd__nor2_1
XFILLER_144_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17148_ _17134_/B _16977_/A _17131_/X _17147_/X vssd1 vssd1 vccd1 vccd1 _17573_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_115_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_495 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09970_ _09970_/A _09970_/B vssd1 vssd1 vccd1 vccd1 _10097_/A sky130_fd_sc_hd__or2_1
X_17079_ _16917_/A _17067_/Y _17068_/X _17078_/X vssd1 vssd1 vccd1 vccd1 _17079_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_171_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08921_ _09078_/A _08947_/B _12258_/B _12256_/C vssd1 vssd1 vccd1 vccd1 _08922_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_118_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08852_ _11895_/B _11895_/D _11902_/B _17379_/A vssd1 vssd1 vccd1 vccd1 _08854_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_112_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_747 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08783_ _08783_/A _08783_/B _08783_/C vssd1 vssd1 vccd1 vccd1 _08801_/B sky130_fd_sc_hd__or3_1
XFILLER_57_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_791 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09404_ _09404_/A _09404_/B vssd1 vssd1 vccd1 vccd1 _09434_/A sky130_fd_sc_hd__xnor2_1
XFILLER_80_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09335_ _09335_/A vssd1 vssd1 vccd1 vccd1 _09335_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09266_ _17399_/A _09555_/D _12174_/D _17403_/A vssd1 vssd1 vccd1 vccd1 _09266_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_139_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09197_ _09227_/A _09197_/B vssd1 vssd1 vccd1 vccd1 _09198_/C sky130_fd_sc_hd__and2_1
XFILLER_5_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10110_ _10109_/B _10594_/B _17479_/Q _10236_/A vssd1 vssd1 vccd1 vccd1 _10110_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_171_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11090_ _11090_/A _11090_/B vssd1 vssd1 vccd1 vccd1 _11153_/A sky130_fd_sc_hd__nor2_1
XFILLER_136_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10041_ _10042_/A _10042_/C vssd1 vssd1 vccd1 vccd1 _10046_/B sky130_fd_sc_hd__nor2_1
XFILLER_88_563 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_31 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13800_ _13800_/A _13800_/B _13800_/C vssd1 vssd1 vccd1 vccd1 _13801_/B sky130_fd_sc_hd__and3_1
XFILLER_29_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11992_ _12155_/A _11991_/B _11971_/X vssd1 vssd1 vccd1 vccd1 _11993_/C sky130_fd_sc_hd__o21ba_1
XFILLER_63_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14780_ _16317_/A _16014_/A vssd1 vssd1 vccd1 vccd1 _16005_/B sky130_fd_sc_hd__or2_1
XFILLER_56_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10943_ _10943_/A _10943_/B _10943_/C vssd1 vssd1 vccd1 vccd1 _10946_/B sky130_fd_sc_hd__nand3_1
X_13731_ _13936_/A _13732_/B vssd1 vssd1 vccd1 vccd1 _13731_/Y sky130_fd_sc_hd__nand2_1
XFILLER_17_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_143 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16450_ _16450_/A _16450_/B vssd1 vssd1 vccd1 vccd1 _16453_/A sky130_fd_sc_hd__xor2_1
X_10874_ _10874_/A _10879_/A _10874_/C vssd1 vssd1 vccd1 vccd1 _10883_/B sky130_fd_sc_hd__or3_1
X_13662_ _13662_/A _13662_/B _13662_/C vssd1 vssd1 vccd1 vccd1 _13671_/B sky130_fd_sc_hd__or3_1
XFILLER_31_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15401_ _15402_/A _15402_/B _16533_/A vssd1 vssd1 vccd1 vccd1 _15404_/B sky130_fd_sc_hd__and3_1
XFILLER_43_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12613_ _12458_/A _12458_/Y _12611_/X _12612_/Y vssd1 vssd1 vccd1 vccd1 _12631_/A
+ sky130_fd_sc_hd__a211oi_4
XFILLER_43_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16381_ _16381_/A _16381_/B vssd1 vssd1 vccd1 vccd1 _16385_/A sky130_fd_sc_hd__xor2_2
XFILLER_31_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13593_ _13688_/A _13593_/B vssd1 vssd1 vccd1 vccd1 _13595_/B sky130_fd_sc_hd__nor2_1
XFILLER_129_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12544_ _11805_/X _11843_/X _12845_/S vssd1 vssd1 vccd1 vccd1 _12544_/X sky130_fd_sc_hd__mux2_1
X_15332_ _16226_/B _16536_/A vssd1 vssd1 vccd1 vccd1 _15334_/B sky130_fd_sc_hd__nand2_1
XFILLER_157_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15263_ _15143_/X _15262_/X _15305_/C vssd1 vssd1 vccd1 vccd1 _15263_/Y sky130_fd_sc_hd__a21boi_2
X_12475_ _12476_/A _12476_/B _12476_/C vssd1 vssd1 vccd1 vccd1 _12477_/A sky130_fd_sc_hd__a21oi_1
XFILLER_8_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17002_ _17003_/A _17003_/B _17003_/C vssd1 vssd1 vccd1 vccd1 _17090_/A sky130_fd_sc_hd__a21o_1
XFILLER_8_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11426_ _11426_/A _11426_/B _11426_/C vssd1 vssd1 vccd1 vccd1 _11433_/A sky130_fd_sc_hd__nand3_1
X_14214_ _14214_/A _14214_/B vssd1 vssd1 vccd1 vccd1 _14216_/A sky130_fd_sc_hd__nor2_1
XANTENNA_6 _17523_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15194_ _15237_/A1 _11853_/Y _12401_/B _15178_/X _15193_/X vssd1 vssd1 vccd1 vccd1
+ _15194_/X sky130_fd_sc_hd__o311a_1
XFILLER_137_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_944 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14145_ _14145_/A _14145_/B vssd1 vssd1 vccd1 vccd1 _14146_/B sky130_fd_sc_hd__and2_1
X_11357_ _11357_/A _11357_/B vssd1 vssd1 vccd1 vccd1 _11359_/B sky130_fd_sc_hd__xor2_1
XFILLER_152_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10308_ _10430_/A _10308_/B vssd1 vssd1 vccd1 vccd1 _10309_/C sky130_fd_sc_hd__and2_1
X_14076_ _14077_/A _14077_/B vssd1 vssd1 vccd1 vccd1 _14188_/A sky130_fd_sc_hd__nand2_1
X_11288_ _11288_/A _11291_/B _11288_/C vssd1 vssd1 vccd1 vccd1 _11351_/A sky130_fd_sc_hd__nand3_1
XFILLER_98_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13027_ _13027_/A _13027_/B vssd1 vssd1 vccd1 vccd1 _13029_/A sky130_fd_sc_hd__nor2_1
X_10239_ _10366_/A _11027_/C _10365_/B _10236_/X vssd1 vssd1 vccd1 vccd1 _10246_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_6_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14978_ _14978_/A _14978_/B vssd1 vssd1 vccd1 vccd1 _14978_/Y sky130_fd_sc_hd__nor2_1
XFILLER_63_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16717_ _16566_/Y _16854_/C _16716_/Y vssd1 vssd1 vccd1 vccd1 _16717_/Y sky130_fd_sc_hd__a21oi_1
X_13929_ _13929_/A _13929_/B vssd1 vssd1 vccd1 vccd1 _13932_/A sky130_fd_sc_hd__xor2_1
XFILLER_63_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16648_ _17156_/B _16648_/B _16648_/C vssd1 vssd1 vccd1 vccd1 _16648_/X sky130_fd_sc_hd__or3_1
XFILLER_22_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_1030 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16579_ _16579_/A _16651_/B _16579_/C vssd1 vssd1 vccd1 vccd1 _16579_/X sky130_fd_sc_hd__or3_1
XFILLER_148_502 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09120_ _09119_/A _09119_/Y _09015_/X _09017_/Y vssd1 vssd1 vccd1 vccd1 _09122_/A
+ sky130_fd_sc_hd__a211oi_2
X_09051_ _09051_/A _09051_/B _09051_/C vssd1 vssd1 vccd1 vccd1 _09071_/A sky130_fd_sc_hd__and3_1
XFILLER_163_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_571 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09953_ _09953_/A _09953_/B vssd1 vssd1 vccd1 vccd1 _10078_/B sky130_fd_sc_hd__xnor2_1
XFILLER_44_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08904_ _08904_/A _08904_/B _08904_/C vssd1 vssd1 vccd1 vccd1 _08905_/C sky130_fd_sc_hd__nand3_1
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09884_ _09884_/A _09884_/B vssd1 vssd1 vccd1 vccd1 _09885_/C sky130_fd_sc_hd__xnor2_1
XFILLER_97_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08835_ _09728_/B _09321_/D _09319_/C _08913_/A vssd1 vssd1 vccd1 vccd1 _08835_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_97_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_844 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08766_ _08766_/A _08766_/B vssd1 vssd1 vccd1 vccd1 _08783_/A sky130_fd_sc_hd__xnor2_4
XFILLER_39_983 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_474 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_88 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09318_ _09318_/A _09318_/B vssd1 vssd1 vccd1 vccd1 _09332_/A sky130_fd_sc_hd__nand2_1
XFILLER_167_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10590_ _11027_/A _11006_/C _11027_/C _10591_/A vssd1 vssd1 vccd1 vccd1 _10593_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_167_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09249_ _09248_/B _09248_/C _09248_/A vssd1 vssd1 vccd1 vccd1 _09249_/X sky130_fd_sc_hd__a21o_1
XFILLER_166_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12260_ _12261_/A _12261_/B vssd1 vssd1 vccd1 vccd1 _12454_/A sky130_fd_sc_hd__nand2b_1
XFILLER_108_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11211_ _11719_/B _11211_/B vssd1 vssd1 vccd1 vccd1 _11217_/A sky130_fd_sc_hd__nand2_1
XFILLER_108_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12191_ _12192_/A _12192_/B vssd1 vssd1 vccd1 vccd1 _12191_/X sky130_fd_sc_hd__and2b_1
XFILLER_162_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_722 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11142_ _11110_/A _11110_/C _11110_/B vssd1 vssd1 vccd1 vccd1 _11143_/D sky130_fd_sc_hd__a21o_1
XFILLER_134_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput76 _17469_/Q vssd1 vssd1 vccd1 vccd1 leds[3] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput87 _17446_/Q vssd1 vssd1 vccd1 vccd1 o_wb_data[12] sky130_fd_sc_hd__clkbuf_1
XFILLER_110_608 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11073_ _11107_/A _11073_/B vssd1 vssd1 vccd1 vccd1 _11074_/B sky130_fd_sc_hd__or2_1
X_15950_ _15577_/Y _16361_/A _15949_/X vssd1 vssd1 vccd1 vccd1 _15953_/A sky130_fd_sc_hd__o21ai_1
Xoutput98 _17456_/Q vssd1 vssd1 vccd1 vccd1 o_wb_data[22] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14901_ _16758_/A _16938_/A vssd1 vssd1 vccd1 vccd1 _15205_/A sky130_fd_sc_hd__or2_1
XFILLER_0_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10024_ _10023_/B _10023_/C _10023_/A vssd1 vssd1 vccd1 vccd1 _10027_/C sky130_fd_sc_hd__a21o_1
XFILLER_163_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15881_ _15881_/A _15881_/B vssd1 vssd1 vccd1 vccd1 _15881_/Y sky130_fd_sc_hd__xnor2_1
X_14832_ _14832_/A _17153_/A vssd1 vssd1 vccd1 vccd1 _17151_/B sky130_fd_sc_hd__or2_1
XFILLER_91_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_279 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17551_ fanout938/X _17551_/D vssd1 vssd1 vccd1 vccd1 _17551_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14763_ _14758_/Y _14762_/Y _14763_/S vssd1 vssd1 vccd1 vccd1 _17606_/D sky130_fd_sc_hd__mux2_1
XFILLER_91_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11975_ _08989_/A _08991_/B _08989_/B vssd1 vssd1 vccd1 vccd1 _11982_/A sky130_fd_sc_hd__o21ba_1
XFILLER_72_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16502_ _16595_/A _16813_/B vssd1 vssd1 vccd1 vccd1 _16670_/A sky130_fd_sc_hd__nor2_2
XFILLER_60_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13714_ _13713_/A _13713_/B _13713_/C vssd1 vssd1 vccd1 vccd1 _13714_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_72_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10926_ _10926_/A _10926_/B vssd1 vssd1 vccd1 vccd1 _10928_/B sky130_fd_sc_hd__xnor2_1
XFILLER_147_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17482_ fanout949/X _17482_/D vssd1 vssd1 vccd1 vccd1 _17482_/Q sky130_fd_sc_hd__dfxtp_1
X_14694_ _14693_/A _14693_/B _14693_/C vssd1 vssd1 vccd1 vccd1 _14695_/B sky130_fd_sc_hd__a21oi_1
XFILLER_16_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16433_ _16152_/A _16809_/C _16432_/C vssd1 vssd1 vccd1 vccd1 _16434_/B sky130_fd_sc_hd__a21oi_1
X_10857_ _10859_/B _10859_/C _10859_/A vssd1 vssd1 vccd1 vccd1 _10857_/Y sky130_fd_sc_hd__a21oi_1
X_13645_ _13749_/A _13645_/B _13645_/C vssd1 vssd1 vccd1 vccd1 _13749_/B sky130_fd_sc_hd__nand3_1
XFILLER_71_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16364_ _16363_/B _16364_/B vssd1 vssd1 vccd1 vccd1 _16365_/B sky130_fd_sc_hd__and2b_1
XFILLER_82_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10788_ _10901_/A _10787_/Y _10792_/A _10897_/B vssd1 vssd1 vccd1 vccd1 _10901_/B
+ sky130_fd_sc_hd__and4bb_1
XFILLER_9_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13576_ _13576_/A _13576_/B _13576_/C vssd1 vssd1 vccd1 vccd1 _13577_/B sky130_fd_sc_hd__and3_1
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15315_ _16015_/A _15381_/B _15315_/C vssd1 vssd1 vccd1 vccd1 _15315_/X sky130_fd_sc_hd__or3_1
XFILLER_145_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12527_ _12355_/A _12355_/B _12356_/X vssd1 vssd1 vccd1 vccd1 _12528_/C sky130_fd_sc_hd__o21ba_1
X_16295_ _16295_/A _16295_/B vssd1 vssd1 vccd1 vccd1 _16296_/B sky130_fd_sc_hd__xnor2_1
XFILLER_172_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15246_ _12858_/Y _15252_/B _15245_/X _16011_/A vssd1 vssd1 vccd1 vccd1 _15246_/X
+ sky130_fd_sc_hd__o22a_1
X_12458_ _12458_/A _12458_/B _12626_/B _12458_/D vssd1 vssd1 vccd1 vccd1 _12458_/Y
+ sky130_fd_sc_hd__nand4_4
X_11409_ _11408_/A _11458_/A vssd1 vssd1 vccd1 vccd1 _11411_/B sky130_fd_sc_hd__and2b_1
X_12389_ _12022_/Y _12024_/Y _14948_/A vssd1 vssd1 vccd1 vccd1 _12389_/X sky130_fd_sc_hd__mux2_1
X_15177_ _15174_/Y _15175_/X _15176_/Y vssd1 vssd1 vccd1 vccd1 _15177_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_113_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14128_ _12219_/X _14210_/B _14482_/B1 vssd1 vssd1 vccd1 vccd1 _14128_/X sky130_fd_sc_hd__o21a_1
XFILLER_114_958 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14059_ _14058_/A _14058_/B _14060_/A vssd1 vssd1 vccd1 vccd1 _14192_/A sky130_fd_sc_hd__a21o_1
XFILLER_79_360 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_875 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09103_ _09103_/A _09103_/B vssd1 vssd1 vccd1 vccd1 _09110_/A sky130_fd_sc_hd__xnor2_1
XFILLER_149_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09034_ _09262_/A _09262_/B vssd1 vssd1 vccd1 vccd1 _09048_/C sky130_fd_sc_hd__nand2_1
XFILLER_163_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout800 _10525_/D vssd1 vssd1 vccd1 vccd1 _15709_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_132_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout811 _11281_/B vssd1 vssd1 vccd1 vccd1 _15624_/A sky130_fd_sc_hd__buf_4
XFILLER_132_777 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout822 _10255_/B vssd1 vssd1 vccd1 vccd1 _10736_/D sky130_fd_sc_hd__clkbuf_2
X_09936_ _09936_/A _09936_/B vssd1 vssd1 vccd1 vccd1 _10078_/A sky130_fd_sc_hd__nor2_1
Xfanout833 _17486_/Q vssd1 vssd1 vccd1 vccd1 _10875_/C sky130_fd_sc_hd__buf_2
Xfanout844 _12463_/D vssd1 vssd1 vccd1 vccd1 _09985_/D sky130_fd_sc_hd__clkbuf_2
Xfanout855 _09128_/B vssd1 vssd1 vccd1 vccd1 _09838_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_86_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout866 _17306_/A1 vssd1 vssd1 vccd1 vccd1 _09979_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_98_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout877 _17304_/A1 vssd1 vssd1 vccd1 vccd1 _11920_/D sky130_fd_sc_hd__buf_2
X_09867_ _09867_/A _09867_/B vssd1 vssd1 vccd1 vccd1 _09868_/B sky130_fd_sc_hd__nor2_1
XFILLER_97_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_555 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout888 _17302_/A1 vssd1 vssd1 vccd1 vccd1 _15402_/A sky130_fd_sc_hd__clkbuf_4
Xfanout899 fanout904/X vssd1 vssd1 vccd1 vccd1 _11468_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08818_ _08812_/A _08814_/B _08812_/B vssd1 vssd1 vccd1 vccd1 _08822_/A sky130_fd_sc_hd__o21ba_1
XTAP_3226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09798_ _09514_/B _10446_/B _15003_/B _09942_/A vssd1 vssd1 vccd1 vccd1 _09798_/Y
+ sky130_fd_sc_hd__a22oi_1
XTAP_3237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08749_ _12070_/A _11859_/D vssd1 vssd1 vccd1 vccd1 _08750_/B sky130_fd_sc_hd__nand2_1
XTAP_2525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11760_ _16727_/B _16795_/A _16568_/B _16641_/A vssd1 vssd1 vccd1 vccd1 _11760_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_27_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10711_ _10711_/A _10711_/B vssd1 vssd1 vccd1 vccd1 _10729_/B sky130_fd_sc_hd__xnor2_2
XFILLER_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11691_ _15303_/A _11691_/B vssd1 vssd1 vccd1 vccd1 _11691_/Y sky130_fd_sc_hd__nor2_1
XTAP_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10642_ _10745_/C _10534_/D _10535_/A _10533_/Y vssd1 vssd1 vccd1 vccd1 _10644_/C
+ sky130_fd_sc_hd__o2bb2a_1
X_13430_ _13430_/A _13430_/B vssd1 vssd1 vccd1 vccd1 _13431_/C sky130_fd_sc_hd__and2_1
XFILLER_13_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13361_ _13361_/A _13361_/B vssd1 vssd1 vccd1 vccd1 _13363_/B sky130_fd_sc_hd__nor2_1
XFILLER_127_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10573_ _10557_/X _10572_/X _10458_/X _10472_/Y vssd1 vssd1 vccd1 vccd1 _10573_/X
+ sky130_fd_sc_hd__a211o_2
XFILLER_167_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15100_ _15100_/A _15100_/B vssd1 vssd1 vccd1 vccd1 _15100_/Y sky130_fd_sc_hd__nand2_1
X_12312_ _12312_/A _12312_/B _12312_/C vssd1 vssd1 vccd1 vccd1 _12314_/A sky130_fd_sc_hd__nand3_1
X_16080_ _16080_/A _16080_/B _16080_/C vssd1 vssd1 vccd1 vccd1 _16081_/B sky130_fd_sc_hd__or3_1
X_13292_ _13292_/A _13292_/B vssd1 vssd1 vccd1 vccd1 _13293_/B sky130_fd_sc_hd__or2_1
XFILLER_166_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12243_ _12722_/A _12722_/B _13450_/C _13334_/C vssd1 vssd1 vccd1 vccd1 _12429_/A
+ sky130_fd_sc_hd__and4_1
X_15031_ _15030_/A _15089_/S _15093_/A _15030_/D vssd1 vssd1 vccd1 vccd1 _15031_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_154_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12174_ _17419_/A _17417_/A _12338_/D _12174_/D vssd1 vssd1 vccd1 vccd1 _12175_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_174_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11125_ _11125_/A _11264_/A vssd1 vssd1 vccd1 vccd1 _11257_/A sky130_fd_sc_hd__or2_1
XFILLER_111_917 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16982_ _16982_/A _16982_/B _17038_/C vssd1 vssd1 vccd1 vccd1 _17040_/A sky130_fd_sc_hd__or3_1
XFILLER_95_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11056_ _11157_/B _11055_/B _11055_/C _11055_/D vssd1 vssd1 vccd1 vccd1 _11056_/Y
+ sky130_fd_sc_hd__a22oi_2
X_15933_ _15933_/A _15933_/B vssd1 vssd1 vccd1 vccd1 _15935_/A sky130_fd_sc_hd__nand2_1
XFILLER_95_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10007_ _10007_/A _10007_/B vssd1 vssd1 vccd1 vccd1 _10009_/C sky130_fd_sc_hd__xnor2_1
XFILLER_92_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15864_ _15864_/A _15864_/B vssd1 vssd1 vccd1 vccd1 _15866_/C sky130_fd_sc_hd__xnor2_1
XFILLER_77_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17603_ fanout934/X _17603_/D vssd1 vssd1 vccd1 vccd1 _17603_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14815_ _16302_/B _16302_/C _16302_/A vssd1 vssd1 vccd1 vccd1 _16398_/A sky130_fd_sc_hd__a21bo_1
XFILLER_92_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15795_ _16136_/A _16209_/B _15811_/A vssd1 vssd1 vccd1 vccd1 _15797_/A sky130_fd_sc_hd__a21bo_1
X_17534_ fanout943/X _17534_/D vssd1 vssd1 vccd1 vccd1 _17534_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_923 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14746_ _14747_/A _14747_/B _14747_/C vssd1 vssd1 vccd1 vccd1 _14748_/A sky130_fd_sc_hd__a21oi_1
X_11958_ _11958_/A _11958_/B _11958_/C vssd1 vssd1 vccd1 vccd1 _11960_/A sky130_fd_sc_hd__or3_1
XFILLER_32_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10909_ _10909_/A _10909_/B vssd1 vssd1 vccd1 vccd1 _11073_/B sky130_fd_sc_hd__xnor2_1
X_17465_ fanout936/X _17465_/D vssd1 vssd1 vccd1 vccd1 _17465_/Q sky130_fd_sc_hd__dfxtp_2
X_14677_ _14677_/A _14677_/B vssd1 vssd1 vccd1 vccd1 _14688_/A sky130_fd_sc_hd__xnor2_1
X_11889_ _12118_/B _11889_/B vssd1 vssd1 vccd1 vccd1 _11891_/C sky130_fd_sc_hd__nand2_1
X_16416_ _16416_/A _16497_/A _16662_/C _16662_/D vssd1 vssd1 vccd1 vccd1 _16519_/A
+ sky130_fd_sc_hd__or4_1
XFILLER_149_129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13628_ _13831_/S _13628_/B vssd1 vssd1 vccd1 vccd1 _13628_/Y sky130_fd_sc_hd__nand2_1
XFILLER_158_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17396_ input43/X _17422_/A2 _17395_/X _17408_/C1 vssd1 vssd1 vccd1 vccd1 _17526_/D
+ sky130_fd_sc_hd__o211a_1
X_16347_ _16347_/A _16347_/B _16345_/X vssd1 vssd1 vccd1 vccd1 _16348_/B sky130_fd_sc_hd__or3b_1
XFILLER_118_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13559_ _13559_/A vssd1 vssd1 vccd1 vccd1 _13559_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16278_ _16279_/B _16279_/C _16279_/A vssd1 vssd1 vccd1 vccd1 _16280_/A sky130_fd_sc_hd__o21a_1
XFILLER_146_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15229_ _15230_/A _15230_/B vssd1 vssd1 vccd1 vccd1 _15231_/A sky130_fd_sc_hd__or2_1
XFILLER_172_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_327 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout129 _17225_/A2 vssd1 vssd1 vccd1 vccd1 _17273_/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_68_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09721_ _09721_/A _09721_/B _09739_/B vssd1 vssd1 vccd1 vccd1 _09768_/B sky130_fd_sc_hd__and3_1
XFILLER_80_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09652_ _15254_/S _12025_/B _09652_/C vssd1 vssd1 vccd1 vccd1 _09655_/A sky130_fd_sc_hd__and3_1
XFILLER_95_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_994 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09583_ _09583_/A _09583_/B vssd1 vssd1 vccd1 vccd1 _09589_/A sky130_fd_sc_hd__nor2_1
XFILLER_83_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09017_ _09016_/A _09016_/B _09016_/C vssd1 vssd1 vccd1 vccd1 _09017_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_163_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout630 _17139_/A vssd1 vssd1 vccd1 vccd1 _12592_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_144_55 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout641 _14008_/B vssd1 vssd1 vccd1 vccd1 _13738_/B sky130_fd_sc_hd__buf_2
Xfanout652 _17028_/A vssd1 vssd1 vccd1 vccd1 _14366_/B sky130_fd_sc_hd__clkbuf_4
X_09919_ _09919_/A _09919_/B vssd1 vssd1 vccd1 vccd1 _09920_/B sky130_fd_sc_hd__or2_1
XFILLER_120_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout663 _12445_/D vssd1 vssd1 vccd1 vccd1 _11895_/D sky130_fd_sc_hd__clkbuf_4
Xfanout674 _17502_/Q vssd1 vssd1 vccd1 vccd1 _14065_/B sky130_fd_sc_hd__buf_4
XFILLER_59_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout685 fanout690/X vssd1 vssd1 vccd1 vccd1 _16789_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_101_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12930_ _12931_/A _12931_/B vssd1 vssd1 vccd1 vccd1 _13117_/B sky130_fd_sc_hd__nand2_1
Xfanout696 fanout699/X vssd1 vssd1 vccd1 vccd1 _12256_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_59_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12861_ _12383_/X _12385_/X _12865_/S vssd1 vssd1 vccd1 vccd1 _12861_/X sky130_fd_sc_hd__mux2_1
XTAP_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_355 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14600_ _14600_/A _14600_/B vssd1 vssd1 vccd1 vccd1 _14601_/C sky130_fd_sc_hd__nor2_1
XTAP_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11812_ _14978_/A _14979_/B _12046_/A vssd1 vssd1 vccd1 vccd1 _12546_/C sky130_fd_sc_hd__o21a_1
XTAP_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15580_ _15580_/A _15580_/B vssd1 vssd1 vccd1 vccd1 _15582_/A sky130_fd_sc_hd__nor2_1
XFILLER_27_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12792_ _12792_/A _12792_/B _12792_/C vssd1 vssd1 vccd1 vccd1 _12794_/A sky130_fd_sc_hd__nor3_1
XTAP_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14531_ _14531_/A _14531_/B _14531_/C vssd1 vssd1 vccd1 vccd1 _14532_/B sky130_fd_sc_hd__or3_1
XTAP_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11743_ _11732_/A _11732_/C _11732_/B vssd1 vssd1 vccd1 vccd1 _11745_/B sky130_fd_sc_hd__o21bai_1
XTAP_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17250_ _17560_/Q _17289_/B vssd1 vssd1 vccd1 vccd1 _17250_/X sky130_fd_sc_hd__and2_1
XFILLER_159_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14462_ _14518_/B _14460_/X _14382_/A _14395_/Y vssd1 vssd1 vccd1 vccd1 _14463_/C
+ sky130_fd_sc_hd__a211o_1
XTAP_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11674_ _11674_/A _11674_/B vssd1 vssd1 vccd1 vccd1 _15235_/A sky130_fd_sc_hd__or2_1
XFILLER_30_959 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16201_ _16382_/A _16201_/B vssd1 vssd1 vccd1 vccd1 _16203_/B sky130_fd_sc_hd__or2_1
XFILLER_41_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13413_ _13414_/B _13852_/B _14181_/B _13658_/A vssd1 vssd1 vccd1 vccd1 _13415_/A
+ sky130_fd_sc_hd__a22oi_1
X_10625_ _10970_/A _10786_/B _10528_/A _10526_/Y vssd1 vssd1 vccd1 vccd1 _10626_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_17181_ _17191_/A _17181_/B _17181_/C _17181_/D vssd1 vssd1 vccd1 vccd1 wire215/A
+ sky130_fd_sc_hd__nor4_1
X_14393_ _14393_/A _14393_/B _14393_/C vssd1 vssd1 vccd1 vccd1 _14394_/B sky130_fd_sc_hd__and3_1
X_16132_ _16133_/A _16133_/B vssd1 vssd1 vccd1 vccd1 _16241_/A sky130_fd_sc_hd__and2_1
XFILLER_127_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10556_ _10555_/A _10556_/B vssd1 vssd1 vccd1 vccd1 _10571_/B sky130_fd_sc_hd__and2b_1
X_13344_ _13462_/B _13344_/B vssd1 vssd1 vccd1 vccd1 _13346_/C sky130_fd_sc_hd__nand2_1
XFILLER_128_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16063_ _15955_/Y _16168_/C vssd1 vssd1 vccd1 vccd1 _16064_/B sky130_fd_sc_hd__and2b_1
XFILLER_127_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10487_ _10487_/A _10487_/B vssd1 vssd1 vccd1 vccd1 _10489_/B sky130_fd_sc_hd__xnor2_1
X_13275_ _12213_/X _12225_/X _13831_/S vssd1 vssd1 vccd1 vccd1 _13276_/B sky130_fd_sc_hd__mux2_1
XFILLER_108_571 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15014_ _14963_/X _14990_/X _15005_/X vssd1 vssd1 vccd1 vccd1 _15014_/Y sky130_fd_sc_hd__o21ai_1
X_12226_ _12222_/X _12225_/X _13833_/S vssd1 vssd1 vccd1 vccd1 _12226_/X sky130_fd_sc_hd__mux2_1
XFILLER_170_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12157_ _12787_/B _12320_/D _12158_/D _17413_/A vssd1 vssd1 vccd1 vccd1 _12161_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_78_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11108_ _11252_/A _11252_/B vssd1 vssd1 vccd1 vccd1 _11110_/B sky130_fd_sc_hd__nor2_1
XFILLER_78_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12088_ _17391_/A _17389_/A _12256_/D _12088_/D vssd1 vssd1 vccd1 vccd1 _12089_/B
+ sky130_fd_sc_hd__and4_1
X_16965_ _16974_/A _16965_/B _16965_/C vssd1 vssd1 vccd1 vccd1 _16966_/B sky130_fd_sc_hd__and3b_1
X_11039_ _11046_/A _11040_/B vssd1 vssd1 vccd1 vccd1 _11039_/Y sky130_fd_sc_hd__nand2b_1
X_15916_ _16129_/A _16743_/C _17043_/B _15918_/A vssd1 vssd1 vccd1 vccd1 _15916_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_83_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16896_ _16952_/B _16896_/B vssd1 vssd1 vccd1 vccd1 _16897_/C sky130_fd_sc_hd__and2_1
XFILLER_94_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15847_ _15846_/A _16355_/B _15846_/B vssd1 vssd1 vccd1 vccd1 _15848_/B sky130_fd_sc_hd__a21oi_1
XFILLER_64_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15778_ _15877_/B _15778_/B vssd1 vssd1 vccd1 vccd1 _15781_/A sky130_fd_sc_hd__or2_1
XFILLER_91_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17517_ fanout950/X _17517_/D vssd1 vssd1 vccd1 vccd1 _17517_/Q sky130_fd_sc_hd__dfxtp_4
X_14729_ _14729_/A _14729_/B vssd1 vssd1 vccd1 vccd1 _14731_/B sky130_fd_sc_hd__nor2_1
XFILLER_32_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17448_ fanout934/X _17448_/D vssd1 vssd1 vccd1 vccd1 _17448_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17379_ _17379_/A _17389_/B vssd1 vssd1 vccd1 vccd1 _17379_/X sky130_fd_sc_hd__or2_1
XFILLER_146_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_168 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09704_ _09835_/A _09835_/B vssd1 vssd1 vccd1 vccd1 _09718_/C sky130_fd_sc_hd__nand2_1
XFILLER_96_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09635_ _09639_/C _10072_/B _09517_/A _09515_/Y vssd1 vssd1 vccd1 vccd1 _09636_/B
+ sky130_fd_sc_hd__o2bb2a_1
Xwb_buttons_leds_959 vssd1 vssd1 vccd1 vccd1 wb_buttons_leds_959/HI led_enb[1] sky130_fd_sc_hd__conb_1
XFILLER_82_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09566_ _10254_/A _10014_/D vssd1 vssd1 vccd1 vccd1 _16982_/B sky130_fd_sc_hd__nand2_2
XFILLER_70_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09497_ _09497_/A _09504_/A _09497_/C vssd1 vssd1 vccd1 vccd1 _09498_/B sky130_fd_sc_hd__nor3_1
XFILLER_12_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_747 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10410_ _10315_/X _10408_/Y _10402_/Y _10402_/A vssd1 vssd1 vccd1 vccd1 _10410_/Y
+ sky130_fd_sc_hd__o211ai_1
XFILLER_20_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11390_ _11387_/C _11389_/X _11393_/B vssd1 vssd1 vccd1 vccd1 _11436_/B sky130_fd_sc_hd__o21ba_1
XFILLER_125_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10341_ _10352_/A _10340_/B _10337_/X vssd1 vssd1 vccd1 vccd1 _10342_/C sky130_fd_sc_hd__a21o_1
XFILLER_164_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13060_ _13060_/A _13060_/B vssd1 vssd1 vccd1 vccd1 _13061_/C sky130_fd_sc_hd__xnor2_1
X_10272_ _14784_/A _10142_/B _10270_/B _10142_/A vssd1 vssd1 vccd1 vccd1 _10272_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_152_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_850 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12011_ _09538_/A _09538_/B _09536_/A vssd1 vssd1 vccd1 vccd1 _12013_/B sky130_fd_sc_hd__a21oi_1
XFILLER_105_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_382 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout460 _14873_/B vssd1 vssd1 vccd1 vccd1 _16317_/A sky130_fd_sc_hd__buf_4
Xfanout471 _10904_/A vssd1 vssd1 vccd1 vccd1 _11006_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_59_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_970 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16750_ _16750_/A _16750_/B vssd1 vssd1 vccd1 vccd1 _16751_/C sky130_fd_sc_hd__xnor2_1
Xfanout482 _09873_/A vssd1 vssd1 vccd1 vccd1 _17385_/A sky130_fd_sc_hd__clkbuf_4
Xfanout493 _11095_/B vssd1 vssd1 vccd1 vccd1 _10963_/B sky130_fd_sc_hd__buf_2
X_13962_ _14047_/A _13962_/B vssd1 vssd1 vccd1 vccd1 _13964_/B sky130_fd_sc_hd__and2_1
XFILLER_46_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15701_ _11700_/A _11700_/C _11700_/B vssd1 vssd1 vccd1 vccd1 _15701_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12913_ _12913_/A _12913_/B vssd1 vssd1 vccd1 vccd1 _12915_/C sky130_fd_sc_hd__xnor2_1
X_16681_ _16681_/A _16827_/B _16681_/C _16681_/D vssd1 vssd1 vccd1 vccd1 _16682_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_73_130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13893_ _13893_/A _14426_/D vssd1 vssd1 vccd1 vccd1 _16864_/A sky130_fd_sc_hd__nand2_2
XFILLER_94_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15632_ _15628_/A _16219_/A1 _13142_/X _15626_/Y _15631_/X vssd1 vssd1 vccd1 vccd1
+ _15632_/X sky130_fd_sc_hd__o311a_1
XFILLER_46_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12844_ _12221_/X _12223_/X _17367_/A vssd1 vssd1 vccd1 vccd1 _12844_/X sky130_fd_sc_hd__mux2_1
XTAP_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15563_ _15564_/A _15564_/B vssd1 vssd1 vccd1 vccd1 _15563_/Y sky130_fd_sc_hd__nor2_1
X_12775_ _12775_/A _12775_/B vssd1 vssd1 vccd1 vccd1 _12776_/B sky130_fd_sc_hd__nor2_1
XTAP_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17302_ _17302_/A1 _17322_/A2 _17301_/X _17378_/C1 vssd1 vssd1 vccd1 vccd1 _17480_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14514_ _14514_/A _14514_/B vssd1 vssd1 vccd1 vccd1 _14515_/B sky130_fd_sc_hd__or2_1
X_11726_ _11726_/A _11726_/B vssd1 vssd1 vccd1 vccd1 _11727_/B sky130_fd_sc_hd__nand2_1
XTAP_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15494_ _15494_/A _15846_/B vssd1 vssd1 vccd1 vccd1 _15496_/A sky130_fd_sc_hd__and2_1
XFILLER_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17233_ _17445_/Q _17275_/A2 _17231_/X _17232_/X _17275_/C1 vssd1 vssd1 vccd1 vccd1
+ _17445_/D sky130_fd_sc_hd__o221a_1
X_14445_ _14445_/A _14445_/B _14445_/C vssd1 vssd1 vccd1 vccd1 _14446_/C sky130_fd_sc_hd__nand3_1
X_11657_ _11657_/A _11657_/B _11657_/C vssd1 vssd1 vccd1 vccd1 _11658_/D sky130_fd_sc_hd__or3_1
XFILLER_7_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10608_ _10699_/A _10607_/B _10607_/A vssd1 vssd1 vccd1 vccd1 _10610_/B sky130_fd_sc_hd__o21ba_1
X_17164_ _17164_/A _17164_/B _17164_/C _17164_/D vssd1 vssd1 vccd1 vccd1 _17164_/X
+ sky130_fd_sc_hd__or4_1
X_14376_ _14376_/A _14376_/B vssd1 vssd1 vccd1 vccd1 _14378_/C sky130_fd_sc_hd__xor2_1
X_11588_ _11579_/A _11579_/C _11579_/B vssd1 vssd1 vccd1 vccd1 _11614_/B sky130_fd_sc_hd__a21o_1
XFILLER_127_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16115_ _17140_/A _16115_/B _16115_/C vssd1 vssd1 vccd1 vccd1 _16122_/A sky130_fd_sc_hd__or3_1
XFILLER_143_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13327_ _13486_/A _13327_/B vssd1 vssd1 vccd1 vccd1 _13329_/C sky130_fd_sc_hd__nor2_1
X_10539_ _10540_/B _10540_/C _10540_/A vssd1 vssd1 vccd1 vccd1 _10550_/A sky130_fd_sc_hd__a21o_1
X_17095_ _17093_/Y _17095_/B vssd1 vssd1 vccd1 vccd1 _17096_/C sky130_fd_sc_hd__and2b_1
XFILLER_170_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16046_ _16046_/A _16046_/B vssd1 vssd1 vccd1 vccd1 _16048_/B sky130_fd_sc_hd__xnor2_1
XFILLER_115_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13258_ _13258_/A _13258_/B _13258_/C vssd1 vssd1 vccd1 vccd1 _13261_/B sky130_fd_sc_hd__or3_1
XFILLER_171_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12209_ _12374_/A _12018_/B _12375_/A vssd1 vssd1 vccd1 vccd1 _12210_/B sky130_fd_sc_hd__a21o_1
XFILLER_170_499 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13189_ _13189_/A _13189_/B _13189_/C vssd1 vssd1 vccd1 vccd1 _13189_/Y sky130_fd_sc_hd__nand3_1
XFILLER_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_767 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16948_ _16938_/A _09424_/X _15724_/X _16882_/A vssd1 vssd1 vccd1 vccd1 _16950_/B
+ sky130_fd_sc_hd__a31oi_1
XFILLER_38_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16879_ _16933_/A _15801_/A _17083_/A _16878_/X vssd1 vssd1 vccd1 vccd1 _16880_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_38_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09420_ _16983_/A _09415_/A _09415_/B vssd1 vssd1 vccd1 vccd1 _09423_/A sky130_fd_sc_hd__o21ba_1
XFILLER_93_995 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09351_ _09493_/A _12025_/B _14981_/A vssd1 vssd1 vccd1 vccd1 _09351_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_33_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09282_ _10126_/B _10897_/B vssd1 vssd1 vccd1 vccd1 _16990_/A sky130_fd_sc_hd__nand2_4
XFILLER_139_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08997_ _09325_/B _12439_/D _09350_/B _17373_/A vssd1 vssd1 vccd1 vccd1 _08999_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_29_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09618_ _09618_/A _09618_/B _09747_/A vssd1 vssd1 vccd1 vccd1 _09621_/B sky130_fd_sc_hd__nand3_1
X_10890_ _10891_/B _10891_/C _10891_/A vssd1 vssd1 vccd1 vccd1 _11148_/A sky130_fd_sc_hd__o21ai_1
XFILLER_55_185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09549_ _10236_/A _10236_/B _09843_/D _09838_/C vssd1 vssd1 vccd1 vccd1 _09552_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_93_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12560_ _12560_/A _12560_/B vssd1 vssd1 vccd1 vccd1 _12561_/C sky130_fd_sc_hd__xor2_1
XFILLER_70_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11511_ _11468_/Y _11471_/X _11469_/X vssd1 vssd1 vccd1 vccd1 _11512_/C sky130_fd_sc_hd__a21o_1
XFILLER_11_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12491_ _12491_/A _12642_/B vssd1 vssd1 vccd1 vccd1 _12492_/C sky130_fd_sc_hd__nor2_1
XFILLER_156_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14230_ _14230_/A _14230_/B vssd1 vssd1 vccd1 vccd1 _14232_/A sky130_fd_sc_hd__nor2_1
X_11442_ _11442_/A _11442_/B vssd1 vssd1 vccd1 vccd1 _11444_/B sky130_fd_sc_hd__xnor2_1
XFILLER_4_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11373_ _11370_/X _11373_/B vssd1 vssd1 vccd1 vccd1 _11529_/B sky130_fd_sc_hd__and2b_1
XFILLER_165_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14161_ _14161_/A _14161_/B vssd1 vssd1 vccd1 vccd1 _14237_/A sky130_fd_sc_hd__xor2_1
XFILLER_166_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_934 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13112_ _13112_/A _13112_/B vssd1 vssd1 vccd1 vccd1 _13114_/B sky130_fd_sc_hd__xnor2_1
X_10324_ _10445_/A _10324_/B vssd1 vssd1 vccd1 vccd1 _10325_/B sky130_fd_sc_hd__or2_1
XFILLER_124_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14092_ _14092_/A _14092_/B _14092_/C vssd1 vssd1 vccd1 vccd1 _14093_/B sky130_fd_sc_hd__and3_1
XFILLER_153_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13043_ _13043_/A _13043_/B _13043_/C vssd1 vssd1 vccd1 vccd1 _13044_/B sky130_fd_sc_hd__or3_1
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10255_ _10255_/A _10255_/B vssd1 vssd1 vccd1 vccd1 _10372_/A sky130_fd_sc_hd__nand2_1
XFILLER_106_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_691 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10186_ _10331_/A _10186_/B vssd1 vssd1 vccd1 vccd1 _10188_/C sky130_fd_sc_hd__and2_1
XFILLER_78_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16802_ _17143_/A1 _14421_/X _16801_/Y vssd1 vssd1 vccd1 vccd1 _16802_/X sky130_fd_sc_hd__o21a_1
XFILLER_121_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14994_ _15102_/A _14994_/B vssd1 vssd1 vccd1 vccd1 _14994_/Y sky130_fd_sc_hd__nand2_1
Xfanout290 _15056_/A vssd1 vssd1 vccd1 vccd1 _12212_/S sky130_fd_sc_hd__clkbuf_2
X_16733_ _16729_/B _17162_/A2 _16974_/B _16722_/A _16869_/C1 vssd1 vssd1 vccd1 vccd1
+ _16733_/X sky130_fd_sc_hd__a221o_1
X_13945_ _15457_/A _13943_/X _13944_/X vssd1 vssd1 vccd1 vccd1 _13945_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_75_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_984 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16664_ _16935_/B _16809_/C vssd1 vssd1 vccd1 vccd1 _16665_/B sky130_fd_sc_hd__nand2_1
X_13876_ _13977_/B _14213_/D _14141_/D _13977_/A vssd1 vssd1 vccd1 vccd1 _13878_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_62_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15615_ _15615_/A _16207_/B _15615_/C vssd1 vssd1 vccd1 vccd1 _15615_/X sky130_fd_sc_hd__or3_1
X_12827_ _12825_/A _12825_/B _12825_/C vssd1 vssd1 vccd1 vccd1 _12827_/Y sky130_fd_sc_hd__o21ai_1
X_16595_ _16595_/A _16595_/B _16503_/Y vssd1 vssd1 vccd1 vccd1 _16596_/B sky130_fd_sc_hd__or3b_1
XFILLER_34_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_583 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15546_ _16111_/A _15533_/Y _15545_/X _15528_/Y vssd1 vssd1 vccd1 vccd1 _15546_/X
+ sky130_fd_sc_hd__o211a_1
X_12758_ _12759_/A _12759_/B vssd1 vssd1 vccd1 vccd1 _12915_/B sky130_fd_sc_hd__nand2b_1
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11709_ _11465_/A _11464_/B _11708_/A vssd1 vssd1 vccd1 vccd1 _11709_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_129_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15477_ _16315_/B _15559_/A _16416_/A _15473_/X vssd1 vssd1 vccd1 vccd1 _15564_/A
+ sky130_fd_sc_hd__or4b_2
XFILLER_30_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12689_ _12689_/A _12689_/B _12689_/C vssd1 vssd1 vccd1 vccd1 _12691_/A sky130_fd_sc_hd__nor3_1
XFILLER_129_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17216_ _17581_/Q _17225_/A2 _17225_/B1 vssd1 vssd1 vccd1 vccd1 _17216_/X sky130_fd_sc_hd__a21o_1
XFILLER_129_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14428_ _14676_/A _14545_/D vssd1 vssd1 vccd1 vccd1 _14430_/B sky130_fd_sc_hd__nand2_1
XFILLER_128_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17147_ _17167_/B _16485_/A _17137_/X _17146_/X vssd1 vssd1 vccd1 vccd1 _17147_/X
+ sky130_fd_sc_hd__a31o_1
X_14359_ _14641_/B _16859_/A _14360_/D _14641_/A vssd1 vssd1 vccd1 vccd1 _14361_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_116_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17078_ _14826_/X _16485_/A _17069_/Y _17077_/X vssd1 vssd1 vccd1 vccd1 _17078_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_157_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16029_ _16315_/C _16662_/C _15917_/Y vssd1 vssd1 vccd1 vccd1 _16032_/A sky130_fd_sc_hd__o21a_1
X_08920_ _08947_/B _12258_/B _12256_/C _09078_/A vssd1 vssd1 vccd1 vccd1 _08922_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_115_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08851_ _08907_/A _08907_/B vssd1 vssd1 vccd1 vccd1 _08908_/A sky130_fd_sc_hd__and2_1
XFILLER_69_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08782_ _08783_/B _08783_/C _08783_/A vssd1 vssd1 vccd1 vccd1 _08801_/A sky130_fd_sc_hd__o21ai_4
XFILLER_85_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_951 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_848 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09403_ _09437_/A _09437_/B vssd1 vssd1 vccd1 vccd1 _09456_/A sky130_fd_sc_hd__nand2_1
XFILLER_164_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_358 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09334_ _09334_/A _09334_/B _09334_/C vssd1 vssd1 vccd1 vccd1 _09335_/A sky130_fd_sc_hd__and3_1
XFILLER_33_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09265_ _17403_/A _12068_/B _09265_/C _09409_/D vssd1 vssd1 vccd1 vccd1 _09268_/A
+ sky130_fd_sc_hd__and4_1
X_09196_ _09196_/A _09196_/B _09202_/A vssd1 vssd1 vccd1 vccd1 _09197_/B sky130_fd_sc_hd__or3_1
XFILLER_107_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10040_ _10045_/C _10311_/D _10034_/A _09900_/Y vssd1 vssd1 vccd1 vccd1 _10042_/C
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_103_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11991_ _12155_/A _11991_/B _11971_/X vssd1 vssd1 vccd1 vccd1 _12155_/B sky130_fd_sc_hd__nor3b_1
XFILLER_44_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13730_ _13514_/B _13935_/A _13728_/Y vssd1 vssd1 vccd1 vccd1 _13732_/B sky130_fd_sc_hd__o21ba_1
X_10942_ _10943_/A _10943_/B _10943_/C vssd1 vssd1 vccd1 vccd1 _10946_/A sky130_fd_sc_hd__a21o_1
XFILLER_28_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13661_ _13770_/A vssd1 vssd1 vccd1 vccd1 _13671_/A sky130_fd_sc_hd__inv_2
XFILLER_45_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10873_ _10874_/A _10874_/C vssd1 vssd1 vccd1 vccd1 _10879_/B sky130_fd_sc_hd__nor2_1
XFILLER_43_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15400_ _15481_/A _15400_/B vssd1 vssd1 vccd1 vccd1 _15424_/A sky130_fd_sc_hd__or2_1
XPHY_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12612_ _12612_/A _12612_/B _12612_/C vssd1 vssd1 vccd1 vccd1 _12612_/Y sky130_fd_sc_hd__nor3_4
XPHY_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16380_ _16381_/A _16381_/B vssd1 vssd1 vccd1 vccd1 _16563_/A sky130_fd_sc_hd__nand2_1
XPHY_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13592_ _13592_/A _13592_/B vssd1 vssd1 vccd1 vccd1 _13593_/B sky130_fd_sc_hd__and2_1
XFILLER_157_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15331_ _15331_/A _15331_/B vssd1 vssd1 vccd1 vccd1 _15334_/A sky130_fd_sc_hd__xor2_1
XFILLER_12_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12543_ _11832_/X _11838_/X _17367_/A vssd1 vssd1 vccd1 vccd1 _12543_/X sky130_fd_sc_hd__mux2_1
XFILLER_157_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15262_ _15262_/A _15262_/B _15262_/C _15262_/D vssd1 vssd1 vccd1 vccd1 _15262_/X
+ sky130_fd_sc_hd__or4_1
X_12474_ _12474_/A _12474_/B vssd1 vssd1 vccd1 vccd1 _12476_/C sky130_fd_sc_hd__xnor2_1
X_17001_ _17052_/B _17001_/B vssd1 vssd1 vccd1 vccd1 _17003_/C sky130_fd_sc_hd__or2_1
X_14213_ _14213_/A _14213_/B _14213_/C _14213_/D vssd1 vssd1 vccd1 vccd1 _14214_/B
+ sky130_fd_sc_hd__and4_1
X_11425_ _11380_/A _11380_/C _11380_/B vssd1 vssd1 vccd1 vccd1 _11426_/C sky130_fd_sc_hd__o21ai_1
XFILLER_126_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15193_ _14963_/X _16582_/B _15192_/X _14926_/X _15188_/Y vssd1 vssd1 vccd1 vccd1
+ _15193_/X sky130_fd_sc_hd__o221a_1
XANTENNA_7 _17516_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14144_ _14145_/A _14145_/B vssd1 vssd1 vccd1 vccd1 _14229_/B sky130_fd_sc_hd__nor2_1
X_11356_ _11357_/A _11357_/B vssd1 vssd1 vccd1 vccd1 _11416_/A sky130_fd_sc_hd__and2b_1
XFILLER_125_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10307_ _10307_/A _10307_/B vssd1 vssd1 vccd1 vccd1 _10314_/A sky130_fd_sc_hd__nor2_1
XFILLER_4_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14075_ _14165_/A _14075_/B vssd1 vssd1 vccd1 vccd1 _14077_/B sky130_fd_sc_hd__and2_1
X_11287_ _11291_/A _11256_/Y _11272_/Y _11311_/A vssd1 vssd1 vccd1 vccd1 _11288_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_140_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13026_ _13641_/A _13156_/B _13522_/D _14065_/B vssd1 vssd1 vccd1 vccd1 _13027_/B
+ sky130_fd_sc_hd__and4_1
X_10238_ _10366_/A _11027_/C vssd1 vssd1 vccd1 vccd1 _10370_/B sky130_fd_sc_hd__nand2_1
XFILLER_6_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10169_ _10170_/A _10170_/C vssd1 vssd1 vccd1 vccd1 _10174_/B sky130_fd_sc_hd__nor2_1
XFILLER_86_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14977_ _17131_/A _15028_/A _14977_/C vssd1 vssd1 vccd1 vccd1 _14977_/X sky130_fd_sc_hd__and3_1
XFILLER_35_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16716_ _16558_/B _16560_/A _16638_/B vssd1 vssd1 vccd1 vccd1 _16716_/Y sky130_fd_sc_hd__a21oi_2
X_13928_ _13929_/A _13929_/B vssd1 vssd1 vccd1 vccd1 _14030_/B sky130_fd_sc_hd__nand2b_1
XFILLER_47_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16647_ _16647_/A vssd1 vssd1 vccd1 vccd1 _16648_/C sky130_fd_sc_hd__inv_2
X_13859_ _13961_/B _13859_/B vssd1 vssd1 vccd1 vccd1 _13861_/C sky130_fd_sc_hd__or2_1
XFILLER_22_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_1042 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16578_ _16480_/A _16400_/B _16571_/A vssd1 vssd1 vccd1 vccd1 _16579_/C sky130_fd_sc_hd__a21oi_1
XFILLER_148_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15529_ _15472_/A _16209_/B _15541_/A vssd1 vssd1 vccd1 vccd1 _15529_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_148_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09050_ _09050_/A _09261_/A vssd1 vssd1 vccd1 vccd1 _09051_/C sky130_fd_sc_hd__nand2_1
XFILLER_129_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xmax_cap232 _14930_/Y vssd1 vssd1 vccd1 vccd1 fanout230/A sky130_fd_sc_hd__clkbuf_1
XFILLER_171_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09952_ _09952_/A _09952_/B vssd1 vssd1 vccd1 vccd1 _09953_/B sky130_fd_sc_hd__nor2_1
XFILLER_171_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08903_ _08903_/A _08903_/B vssd1 vssd1 vccd1 vccd1 _08905_/B sky130_fd_sc_hd__xnor2_1
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09883_ _09869_/X _09870_/Y _09877_/X _09881_/X vssd1 vssd1 vccd1 vccd1 _09885_/B
+ sky130_fd_sc_hd__a211o_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08834_ _08800_/X _08801_/Y _08832_/A _08832_/Y vssd1 vssd1 vccd1 vccd1 _08874_/B
+ sky130_fd_sc_hd__a211oi_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08765_ _08766_/A _08766_/B vssd1 vssd1 vccd1 vccd1 _11877_/B sky130_fd_sc_hd__nand2b_1
XFILLER_38_450 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_995 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09317_ _09317_/A _09323_/A _09317_/C vssd1 vssd1 vccd1 vccd1 _09318_/B sky130_fd_sc_hd__or3_1
XFILLER_166_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09248_ _09248_/A _09248_/B _09248_/C vssd1 vssd1 vccd1 vccd1 _09248_/Y sky130_fd_sc_hd__nand3_2
XFILLER_167_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09179_ _09179_/A _09179_/B vssd1 vssd1 vccd1 vccd1 _09345_/B sky130_fd_sc_hd__nor2_1
XFILLER_119_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11210_ _11719_/A _11208_/Y _11168_/A _11168_/Y vssd1 vssd1 vccd1 vccd1 _11211_/B
+ sky130_fd_sc_hd__a211o_1
X_12190_ _12190_/A _12190_/B vssd1 vssd1 vccd1 vccd1 _12192_/B sky130_fd_sc_hd__xnor2_1
XFILLER_134_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11141_ _11146_/A _11113_/Y _11128_/Y _11255_/A vssd1 vssd1 vccd1 vccd1 _11143_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_134_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput77 _17470_/Q vssd1 vssd1 vccd1 vccd1 leds[4] sky130_fd_sc_hd__clkbuf_1
X_11072_ _11072_/A _11072_/B _11072_/C vssd1 vssd1 vccd1 vccd1 _11075_/B sky130_fd_sc_hd__and3_1
Xoutput88 _17447_/Q vssd1 vssd1 vccd1 vccd1 o_wb_data[13] sky130_fd_sc_hd__clkbuf_1
Xoutput99 _17457_/Q vssd1 vssd1 vccd1 vccd1 o_wb_data[23] sky130_fd_sc_hd__clkbuf_1
XFILLER_1_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14900_ _17119_/A _16880_/A _15147_/C vssd1 vssd1 vccd1 vccd1 _14900_/X sky130_fd_sc_hd__o21a_1
XFILLER_49_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10023_ _10023_/A _10023_/B _10023_/C vssd1 vssd1 vccd1 vccd1 _10027_/B sky130_fd_sc_hd__nand3_1
XFILLER_76_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15880_ _15881_/A _15881_/B vssd1 vssd1 vccd1 vccd1 _15992_/B sky130_fd_sc_hd__nor2_1
XFILLER_48_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14831_ _17167_/A _17151_/A _17167_/B vssd1 vssd1 vccd1 vccd1 _14831_/Y sky130_fd_sc_hd__nand3_1
XFILLER_56_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17550_ fanout933/X _17550_/D vssd1 vssd1 vccd1 vccd1 _17550_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14762_ _14762_/A _14762_/B vssd1 vssd1 vccd1 vccd1 _14762_/Y sky130_fd_sc_hd__xnor2_1
X_11974_ _09234_/A _09236_/B _09234_/B vssd1 vssd1 vccd1 vccd1 _11984_/A sky130_fd_sc_hd__o21ba_1
X_16501_ _16609_/B _16501_/B vssd1 vssd1 vccd1 vccd1 _16507_/A sky130_fd_sc_hd__and2_1
XFILLER_147_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13713_ _13713_/A _13713_/B _13713_/C vssd1 vssd1 vccd1 vccd1 _13818_/A sky130_fd_sc_hd__or3_1
X_10925_ _10926_/A _10926_/B vssd1 vssd1 vccd1 vccd1 _11049_/B sky130_fd_sc_hd__and2_1
X_17481_ fanout942/X _17481_/D vssd1 vssd1 vccd1 vccd1 _17481_/Q sky130_fd_sc_hd__dfxtp_1
X_14693_ _14693_/A _14693_/B _14693_/C vssd1 vssd1 vccd1 vccd1 _14723_/B sky130_fd_sc_hd__and3_1
XFILLER_72_784 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16432_ _16760_/B _16809_/C _16432_/C vssd1 vssd1 vccd1 vccd1 _16511_/B sky130_fd_sc_hd__and3_1
X_13644_ _13644_/A _13644_/B vssd1 vssd1 vccd1 vccd1 _13645_/C sky130_fd_sc_hd__xnor2_1
XFILLER_72_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10856_ _10865_/A _10865_/B vssd1 vssd1 vccd1 vccd1 _10859_/C sky130_fd_sc_hd__nand2_1
XFILLER_31_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16363_ _16364_/B _16363_/B vssd1 vssd1 vccd1 vccd1 _16365_/A sky130_fd_sc_hd__and2b_1
XFILLER_157_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13575_ _13576_/A _13576_/B _13576_/C vssd1 vssd1 vccd1 vccd1 _13577_/A sky130_fd_sc_hd__a21oi_1
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10787_ _10991_/A _10932_/B _10991_/C vssd1 vssd1 vccd1 vccd1 _10787_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_40_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15314_ _15314_/A _15314_/B vssd1 vssd1 vccd1 vccd1 _15315_/C sky130_fd_sc_hd__nor2_1
X_12526_ _12526_/A _12526_/B _12526_/C vssd1 vssd1 vccd1 vccd1 _12528_/B sky130_fd_sc_hd__and3_1
X_16294_ _16294_/A _16294_/B vssd1 vssd1 vccd1 vccd1 _16295_/B sky130_fd_sc_hd__nor2_1
XFILLER_8_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15245_ _14983_/X _14986_/Y _15384_/S vssd1 vssd1 vccd1 vccd1 _15245_/X sky130_fd_sc_hd__mux2_1
X_12457_ _12458_/A _12458_/B _12626_/B _12458_/D vssd1 vssd1 vccd1 vccd1 _12457_/X
+ sky130_fd_sc_hd__a22o_1
X_11408_ _11408_/A _11408_/B _11408_/C vssd1 vssd1 vccd1 vccd1 _11458_/A sky130_fd_sc_hd__or3_1
XFILLER_67_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15176_ _15119_/A _15119_/B _15117_/A vssd1 vssd1 vccd1 vccd1 _15176_/Y sky130_fd_sc_hd__o21ai_1
X_12388_ _12384_/X _12387_/X _13840_/S vssd1 vssd1 vccd1 vccd1 _12388_/X sky130_fd_sc_hd__mux2_1
XFILLER_153_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_786 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14127_ _12226_/X _12230_/B _14356_/S vssd1 vssd1 vccd1 vccd1 _14127_/X sky130_fd_sc_hd__mux2_1
X_11339_ _11340_/B _11340_/A vssd1 vssd1 vccd1 vccd1 _11406_/A sky130_fd_sc_hd__nand2b_1
XFILLER_114_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14058_ _14058_/A _14058_/B vssd1 vssd1 vccd1 vccd1 _14060_/B sky130_fd_sc_hd__nand2_1
XFILLER_86_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13009_ _13010_/B _13268_/A vssd1 vssd1 vccd1 vccd1 _13009_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_79_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09102_ _09103_/B _09103_/A vssd1 vssd1 vccd1 vccd1 _09153_/A sky130_fd_sc_hd__and2b_1
XFILLER_148_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09033_ _09033_/A _09033_/B vssd1 vssd1 vccd1 vccd1 _09262_/B sky130_fd_sc_hd__xnor2_1
XFILLER_117_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout801 _10525_/D vssd1 vssd1 vccd1 vccd1 _14893_/B sky130_fd_sc_hd__clkbuf_4
X_09935_ _10075_/A _09935_/B vssd1 vssd1 vccd1 vccd1 _09936_/B sky130_fd_sc_hd__and2_1
Xfanout812 _10508_/D vssd1 vssd1 vccd1 vccd1 _10270_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_89_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout823 _09265_/C vssd1 vssd1 vccd1 vccd1 _10255_/B sky130_fd_sc_hd__buf_4
XFILLER_89_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout834 _09409_/D vssd1 vssd1 vccd1 vccd1 _12174_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_98_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout845 _12463_/D vssd1 vssd1 vccd1 vccd1 _12129_/B sky130_fd_sc_hd__buf_2
XFILLER_58_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout856 _12295_/D vssd1 vssd1 vccd1 vccd1 _09128_/B sky130_fd_sc_hd__clkbuf_4
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout867 fanout874/X vssd1 vssd1 vccd1 vccd1 _17306_/A1 sky130_fd_sc_hd__clkbuf_4
X_09866_ _09866_/A _09866_/B _09884_/B vssd1 vssd1 vccd1 vccd1 _09914_/B sky130_fd_sc_hd__and3_1
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout878 _17481_/Q vssd1 vssd1 vccd1 vccd1 _17304_/A1 sky130_fd_sc_hd__buf_2
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout889 _17480_/Q vssd1 vssd1 vccd1 vccd1 _17302_/A1 sky130_fd_sc_hd__buf_2
XFILLER_133_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08817_ _08831_/B _08831_/C _08831_/A vssd1 vssd1 vccd1 vccd1 _08832_/A sky130_fd_sc_hd__o21a_1
XFILLER_58_567 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09797_ _09797_/A _10111_/D _10062_/C vssd1 vssd1 vccd1 vccd1 _09801_/B sky130_fd_sc_hd__and3_1
XTAP_3227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08748_ _08748_/A _08748_/B vssd1 vssd1 vccd1 vccd1 _08750_/A sky130_fd_sc_hd__and2_1
XTAP_2515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10710_ _11180_/A _11180_/B vssd1 vssd1 vccd1 vccd1 _10729_/A sky130_fd_sc_hd__nand2_1
XTAP_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11690_ _11690_/A _11690_/B vssd1 vssd1 vccd1 vccd1 _11691_/B sky130_fd_sc_hd__xnor2_1
XFILLER_53_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10641_ _10641_/A _10724_/A vssd1 vssd1 vccd1 vccd1 _10649_/A sky130_fd_sc_hd__nor2_1
XFILLER_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13360_ _13360_/A _13360_/B vssd1 vssd1 vccd1 vccd1 _13363_/A sky130_fd_sc_hd__xor2_1
XFILLER_166_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10572_ _10572_/A _10572_/B _10586_/B vssd1 vssd1 vccd1 vccd1 _10572_/X sky130_fd_sc_hd__or3_1
XFILLER_166_163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12311_ _12311_/A _12311_/B vssd1 vssd1 vccd1 vccd1 _12312_/C sky130_fd_sc_hd__xor2_1
XFILLER_5_302 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13291_ _13292_/A _13292_/B vssd1 vssd1 vccd1 vccd1 _13411_/B sky130_fd_sc_hd__nand2_1
XFILLER_6_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15030_ _15030_/A _15089_/S _15093_/A _15030_/D vssd1 vssd1 vccd1 vccd1 _15093_/B
+ sky130_fd_sc_hd__nand4_1
X_12242_ _12722_/B _13450_/C _13334_/C _12722_/A vssd1 vssd1 vccd1 vccd1 _12244_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_135_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12173_ _17417_/A _12338_/D _12174_/D _17419_/A vssd1 vssd1 vccd1 vccd1 _12175_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_3_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11124_ _11125_/A _11123_/Y _11124_/C _14895_/B vssd1 vssd1 vccd1 vccd1 _11264_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_96_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16981_ _16974_/A _17170_/B1 _16980_/X vssd1 vssd1 vccd1 vccd1 _17569_/D sky130_fd_sc_hd__a21oi_1
XFILLER_111_929 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11055_ _11157_/B _11055_/B _11055_/C _11055_/D vssd1 vssd1 vccd1 vccd1 _11055_/X
+ sky130_fd_sc_hd__and4_1
X_15932_ _15932_/A _16138_/A _16681_/A _16827_/B vssd1 vssd1 vccd1 vccd1 _15933_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_110_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_480 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10006_ _09991_/Y _10005_/X _09865_/B _09975_/X vssd1 vssd1 vccd1 vccd1 _10028_/A
+ sky130_fd_sc_hd__o211a_1
X_15863_ _15863_/A _15863_/B vssd1 vssd1 vccd1 vccd1 _15864_/B sky130_fd_sc_hd__xnor2_1
XFILLER_37_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_504 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17602_ fanout933/X _17602_/D vssd1 vssd1 vccd1 vccd1 _17602_/Q sky130_fd_sc_hd__dfxtp_1
X_14814_ _14778_/X _14813_/X _08776_/C vssd1 vssd1 vccd1 vccd1 _16302_/C sky130_fd_sc_hd__a21o_1
XFILLER_91_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15794_ _16207_/B _15794_/B _15888_/B vssd1 vssd1 vccd1 vccd1 _15794_/X sky130_fd_sc_hd__or3b_2
XFILLER_91_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17533_ fanout945/X _17533_/D vssd1 vssd1 vccd1 vccd1 _17533_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14745_ _14745_/A _14745_/B vssd1 vssd1 vccd1 vccd1 _14747_/C sky130_fd_sc_hd__xnor2_1
X_11957_ _11957_/A _12163_/B vssd1 vssd1 vccd1 vccd1 _11958_/C sky130_fd_sc_hd__nor2_1
XFILLER_83_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10908_ _11005_/A _17468_/D vssd1 vssd1 vccd1 vccd1 _10909_/B sky130_fd_sc_hd__nand2_1
X_17464_ fanout951/X _17464_/D vssd1 vssd1 vccd1 vccd1 _17464_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_60_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14676_ _14676_/A _14738_/B vssd1 vssd1 vccd1 vccd1 _14677_/B sky130_fd_sc_hd__nand2_1
X_11888_ _11888_/A _11888_/B vssd1 vssd1 vccd1 vccd1 _11889_/B sky130_fd_sc_hd__or2_1
X_16415_ _16497_/A _16662_/C _17043_/B _16505_/A vssd1 vssd1 vccd1 vccd1 _16417_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_32_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13627_ _12702_/X _12704_/X _13627_/S vssd1 vssd1 vccd1 vccd1 _13627_/X sky130_fd_sc_hd__mux2_1
X_10839_ _10933_/A _11122_/B _10933_/D _10970_/B vssd1 vssd1 vccd1 vccd1 _10841_/A
+ sky130_fd_sc_hd__and4_1
X_17395_ _17395_/A _17425_/B vssd1 vssd1 vccd1 vccd1 _17395_/X sky130_fd_sc_hd__or2_1
XFILLER_32_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16346_ _16347_/A _16347_/B _16345_/X vssd1 vssd1 vccd1 vccd1 _16462_/A sky130_fd_sc_hd__o21ba_1
XFILLER_146_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13558_ _13558_/A _13558_/B _13558_/C vssd1 vssd1 vccd1 vccd1 _13559_/A sky130_fd_sc_hd__and3_1
XFILLER_158_675 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12509_ _12509_/A _12509_/B vssd1 vssd1 vccd1 vccd1 _12511_/A sky130_fd_sc_hd__nor2_1
XFILLER_9_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16277_ _16277_/A _16277_/B vssd1 vssd1 vccd1 vccd1 _16283_/A sky130_fd_sc_hd__nand2_1
X_13489_ _13486_/X _13487_/Y _13365_/Y _13369_/B vssd1 vssd1 vccd1 vccd1 _13490_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15228_ _15228_/A _15228_/B vssd1 vssd1 vccd1 vccd1 _15230_/B sky130_fd_sc_hd__xnor2_1
XFILLER_114_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15159_ _15159_/A _15159_/B vssd1 vssd1 vccd1 vccd1 _15161_/B sky130_fd_sc_hd__xnor2_1
XFILLER_141_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09720_ _09720_/A _09866_/A vssd1 vssd1 vccd1 vccd1 _09739_/B sky130_fd_sc_hd__nand2_1
XFILLER_110_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09651_ _11839_/S _14864_/A vssd1 vssd1 vccd1 vccd1 _09652_/C sky130_fd_sc_hd__and2_1
XFILLER_110_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09582_ _09730_/C _09446_/D _09447_/A _09445_/Y vssd1 vssd1 vccd1 vccd1 _09583_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_42_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09016_ _09016_/A _09016_/B _09016_/C vssd1 vssd1 vccd1 vccd1 _09016_/Y sky130_fd_sc_hd__nand3_1
XFILLER_117_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout620 _08967_/B vssd1 vssd1 vccd1 vccd1 _17153_/A sky130_fd_sc_hd__buf_2
Xfanout631 _17508_/Q vssd1 vssd1 vccd1 vccd1 _17139_/A sky130_fd_sc_hd__buf_4
XFILLER_99_990 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout642 _13035_/C vssd1 vssd1 vccd1 vccd1 _14008_/B sky130_fd_sc_hd__buf_2
X_09918_ _09912_/B _09912_/C _09912_/A vssd1 vssd1 vccd1 vccd1 _09922_/A sky130_fd_sc_hd__o21bai_1
XFILLER_144_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout653 _17028_/A vssd1 vssd1 vccd1 vccd1 _14593_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_58_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout664 _12025_/B vssd1 vssd1 vccd1 vccd1 _12445_/D sky130_fd_sc_hd__clkbuf_4
Xfanout675 _17502_/Q vssd1 vssd1 vccd1 vccd1 _12877_/C sky130_fd_sc_hd__clkbuf_2
Xfanout686 _12256_/C vssd1 vssd1 vccd1 vccd1 _11900_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_37_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout697 fanout699/X vssd1 vssd1 vccd1 vccd1 _14863_/B sky130_fd_sc_hd__clkbuf_4
X_09849_ _09976_/A _09976_/B vssd1 vssd1 vccd1 vccd1 _09863_/C sky130_fd_sc_hd__nand2_1
XTAP_3002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12860_ _12710_/A _15457_/C _16653_/A vssd1 vssd1 vccd1 vccd1 _12860_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_170_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11811_ _12025_/A _11932_/B vssd1 vssd1 vccd1 vccd1 _14979_/B sky130_fd_sc_hd__and2_1
XTAP_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12791_ _12791_/A _12947_/B vssd1 vssd1 vccd1 vccd1 _12792_/C sky130_fd_sc_hd__nor2_1
XTAP_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14530_ _14531_/A _14531_/B _14531_/C vssd1 vssd1 vccd1 vccd1 _14585_/A sky130_fd_sc_hd__o21ai_1
XTAP_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11742_ _11742_/A _11742_/B vssd1 vssd1 vccd1 vccd1 _11745_/A sky130_fd_sc_hd__or2_1
XFILLER_15_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14461_ _14382_/A _14395_/Y _14518_/B _14460_/X vssd1 vssd1 vccd1 vccd1 _14463_/B
+ sky130_fd_sc_hd__o211ai_2
XTAP_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11673_ _11673_/A _11673_/B vssd1 vssd1 vccd1 vccd1 _11674_/B sky130_fd_sc_hd__nor2_1
XTAP_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16200_ _16200_/A _16200_/B _16200_/C vssd1 vssd1 vccd1 vccd1 _16201_/B sky130_fd_sc_hd__and3_1
X_13412_ _13301_/A _13303_/B _13301_/B vssd1 vssd1 vccd1 vccd1 _13420_/A sky130_fd_sc_hd__o21ba_1
X_10624_ _10624_/A _10624_/B vssd1 vssd1 vccd1 vccd1 _10713_/A sky130_fd_sc_hd__xnor2_1
X_17180_ _17180_/A _17180_/B _17180_/C _17180_/D vssd1 vssd1 vccd1 vccd1 _17181_/D
+ sky130_fd_sc_hd__or4_1
XFILLER_168_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14392_ _14394_/A vssd1 vssd1 vccd1 vccd1 _14471_/A sky130_fd_sc_hd__inv_2
XFILLER_10_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16131_ _15913_/A _16023_/Y _16026_/B _16022_/X vssd1 vssd1 vccd1 vccd1 _16133_/B
+ sky130_fd_sc_hd__a2bb2o_1
X_13343_ _13903_/A _12871_/B _13342_/C vssd1 vssd1 vccd1 vccd1 _13344_/B sky130_fd_sc_hd__a21o_1
X_10555_ _10555_/A _10555_/B _10555_/C vssd1 vssd1 vccd1 vccd1 _10556_/B sky130_fd_sc_hd__or3_1
XFILLER_127_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16062_ _16695_/A _16589_/B _16062_/C vssd1 vssd1 vccd1 vccd1 _16064_/A sky130_fd_sc_hd__and3_1
X_13274_ _12710_/A _13273_/X _16653_/A vssd1 vssd1 vccd1 vccd1 _13274_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_108_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10486_ _10478_/A _10480_/B _10478_/B vssd1 vssd1 vccd1 vccd1 _10489_/A sky130_fd_sc_hd__o21ba_1
XFILLER_136_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15013_ _11655_/A _15804_/A2 _15007_/X _15012_/X vssd1 vssd1 vccd1 vccd1 _15013_/Y
+ sky130_fd_sc_hd__a211oi_2
XFILLER_5_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12225_ _12223_/X _12224_/X _17367_/A vssd1 vssd1 vccd1 vccd1 _12225_/X sky130_fd_sc_hd__mux2_1
XFILLER_108_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12156_ _12156_/A _12156_/B vssd1 vssd1 vccd1 vccd1 _12190_/A sky130_fd_sc_hd__nand2_1
XFILLER_69_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11107_ _11107_/A _11107_/B vssd1 vssd1 vccd1 vccd1 _11252_/B sky130_fd_sc_hd__or2_1
XFILLER_68_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_748 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12087_ _17389_/A _12256_/D _12088_/D _17391_/A vssd1 vssd1 vccd1 vccd1 _12089_/A
+ sky130_fd_sc_hd__a22oi_1
X_16964_ _16965_/C _16965_/B _16974_/A vssd1 vssd1 vccd1 vccd1 _16966_/A sky130_fd_sc_hd__a21boi_1
XFILLER_1_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11038_ _11038_/A _11038_/B vssd1 vssd1 vccd1 vccd1 _11040_/B sky130_fd_sc_hd__xnor2_1
X_15915_ _16028_/A _15915_/B vssd1 vssd1 vccd1 vccd1 _15923_/A sky130_fd_sc_hd__or2_1
XFILLER_49_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16895_ _16895_/A _16895_/B vssd1 vssd1 vccd1 vccd1 _16896_/B sky130_fd_sc_hd__nand2_1
XFILLER_37_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15846_ _15846_/A _15846_/B _16355_/B vssd1 vssd1 vccd1 vccd1 _15848_/A sky130_fd_sc_hd__and3_1
XFILLER_76_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12989_ _12819_/X _12824_/A _12987_/X _12988_/Y vssd1 vssd1 vccd1 vccd1 _12993_/A
+ sky130_fd_sc_hd__a211oi_2
X_15777_ _15877_/A _15776_/B _15776_/C vssd1 vssd1 vccd1 vccd1 _15778_/B sky130_fd_sc_hd__o21a_1
XTAP_3591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17516_ fanout942/X _17516_/D vssd1 vssd1 vccd1 vccd1 _17516_/Q sky130_fd_sc_hd__dfxtp_4
X_14728_ _14726_/X _14728_/B vssd1 vssd1 vccd1 vccd1 _14731_/A sky130_fd_sc_hd__nand2b_1
XTAP_2890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17447_ fanout934/X _17447_/D vssd1 vssd1 vccd1 vccd1 _17447_/Q sky130_fd_sc_hd__dfxtp_1
X_14659_ _14698_/A _14659_/B vssd1 vssd1 vccd1 vccd1 _14662_/A sky130_fd_sc_hd__and2_1
XFILLER_32_275 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17378_ input65/X _17377_/B _17377_/Y _17378_/C1 vssd1 vssd1 vccd1 vccd1 _17517_/D
+ sky130_fd_sc_hd__o211a_1
X_16329_ _16329_/A _16425_/B vssd1 vssd1 vccd1 vccd1 _16331_/A sky130_fd_sc_hd__nor2_1
XFILLER_145_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09703_ _09703_/A _09703_/B vssd1 vssd1 vccd1 vccd1 _09835_/B sky130_fd_sc_hd__xnor2_1
XFILLER_101_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09634_ _09634_/A _09634_/B vssd1 vssd1 vccd1 vccd1 _09645_/A sky130_fd_sc_hd__nor2_1
XFILLER_55_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09565_ _09565_/A _09565_/B vssd1 vssd1 vccd1 vccd1 _09573_/A sky130_fd_sc_hd__xnor2_1
XFILLER_83_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09496_ _09619_/B _09656_/A _09619_/A vssd1 vssd1 vccd1 vccd1 _09620_/A sky130_fd_sc_hd__o21ai_1
XFILLER_169_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_759 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_584 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10340_ _10337_/X _10340_/B vssd1 vssd1 vccd1 vccd1 _10352_/B sky130_fd_sc_hd__and2b_1
XFILLER_136_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10271_ _10271_/A _10743_/D vssd1 vssd1 vccd1 vccd1 _10391_/A sky130_fd_sc_hd__nand2_1
XFILLER_105_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_862 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12010_ _12010_/A _12010_/B vssd1 vssd1 vccd1 vccd1 _12013_/A sky130_fd_sc_hd__xnor2_1
XFILLER_151_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_394 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout450 _09412_/A vssd1 vssd1 vccd1 vccd1 _16021_/A sky130_fd_sc_hd__buf_2
XFILLER_48_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout461 _14873_/B vssd1 vssd1 vccd1 vccd1 _10254_/A sky130_fd_sc_hd__clkbuf_4
Xfanout472 _11790_/A vssd1 vssd1 vccd1 vccd1 _10904_/A sky130_fd_sc_hd__buf_2
X_13961_ _13961_/A _13961_/B _13961_/C vssd1 vssd1 vccd1 vccd1 _13962_/B sky130_fd_sc_hd__or3_1
XFILLER_59_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout483 _09873_/A vssd1 vssd1 vccd1 vccd1 _08913_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_93_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout494 _14784_/A vssd1 vssd1 vccd1 vccd1 _11095_/B sky130_fd_sc_hd__buf_2
XFILLER_87_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12912_ _12913_/A _12913_/B vssd1 vssd1 vccd1 vccd1 _13072_/A sky130_fd_sc_hd__and2_1
XFILLER_46_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15700_ _15700_/A _15700_/B vssd1 vssd1 vccd1 vccd1 _15700_/Y sky130_fd_sc_hd__xnor2_2
X_16680_ _16827_/B _16681_/C _16681_/D _16681_/A vssd1 vssd1 vccd1 vccd1 _16680_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_111_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13892_ _14013_/A _13892_/B vssd1 vssd1 vccd1 vccd1 _13912_/A sky130_fd_sc_hd__nand2_1
XFILLER_58_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_142 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12843_ _16922_/A _12843_/B vssd1 vssd1 vccd1 vccd1 _12856_/A sky130_fd_sc_hd__nand2_1
XTAP_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15631_ _16015_/A _15709_/B _15624_/Y _15628_/X _15630_/X vssd1 vssd1 vccd1 vccd1
+ _15631_/X sky130_fd_sc_hd__o32a_1
XTAP_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15562_ _15655_/A _15655_/B vssd1 vssd1 vccd1 vccd1 _15564_/B sky130_fd_sc_hd__xnor2_1
X_12774_ _12775_/A _12775_/B vssd1 vssd1 vccd1 vccd1 _12931_/A sky130_fd_sc_hd__and2_1
XTAP_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17301_ input58/X _17321_/B _17321_/C vssd1 vssd1 vccd1 vccd1 _17301_/X sky130_fd_sc_hd__or3_1
XTAP_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14513_ _14514_/A _14514_/B vssd1 vssd1 vccd1 vccd1 _14569_/B sky130_fd_sc_hd__nand2_1
XFILLER_159_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11725_ _11725_/A _11725_/B _11725_/C vssd1 vssd1 vccd1 vccd1 _11731_/B sky130_fd_sc_hd__and3_1
XFILLER_14_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15493_ _15493_/A _16747_/A vssd1 vssd1 vccd1 vccd1 _15846_/B sky130_fd_sc_hd__nor2_1
XFILLER_30_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17232_ _17554_/Q _17274_/B vssd1 vssd1 vccd1 vccd1 _17232_/X sky130_fd_sc_hd__and2_1
X_14444_ _14445_/A _14445_/B _14445_/C vssd1 vssd1 vccd1 vccd1 _14508_/A sky130_fd_sc_hd__a21o_1
X_11656_ _11657_/B _11657_/C _11657_/A vssd1 vssd1 vccd1 vccd1 _11681_/A sky130_fd_sc_hd__o21ai_2
XFILLER_156_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10607_ _10607_/A _10607_/B vssd1 vssd1 vccd1 vccd1 _10699_/B sky130_fd_sc_hd__nor2_1
X_17163_ _17151_/A _17163_/A2 _17162_/X vssd1 vssd1 vccd1 vccd1 _17163_/X sky130_fd_sc_hd__o21ba_1
XFILLER_155_420 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14375_ _14376_/B _14376_/A vssd1 vssd1 vccd1 vccd1 _14445_/B sky130_fd_sc_hd__nand2b_1
X_11587_ _11583_/A _11582_/C _11582_/A vssd1 vssd1 vccd1 vccd1 _11587_/X sky130_fd_sc_hd__a21o_1
XFILLER_128_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16114_ _16114_/A _16114_/B vssd1 vssd1 vccd1 vccd1 _16115_/C sky130_fd_sc_hd__nor2_1
X_13326_ _13326_/A _13326_/B _13326_/C vssd1 vssd1 vccd1 vccd1 _13327_/B sky130_fd_sc_hd__nor3_1
XFILLER_6_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17094_ _17093_/A _17093_/B _17093_/C vssd1 vssd1 vccd1 vccd1 _17095_/B sky130_fd_sc_hd__o21ai_1
X_10538_ _10540_/B _10540_/C _10540_/A vssd1 vssd1 vccd1 vccd1 _10538_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_127_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16045_ _16046_/A _16046_/B vssd1 vssd1 vccd1 vccd1 _16045_/X sky130_fd_sc_hd__and2b_1
XFILLER_127_199 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13257_ _13258_/A _13258_/B _13258_/C vssd1 vssd1 vccd1 vccd1 _13261_/A sky130_fd_sc_hd__o21ai_2
XFILLER_170_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10469_ _10469_/A _10469_/B _10469_/C vssd1 vssd1 vccd1 vccd1 _10470_/B sky130_fd_sc_hd__nor3_1
XFILLER_108_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12208_ _12375_/B _12208_/B vssd1 vssd1 vccd1 vccd1 _12374_/B sky130_fd_sc_hd__nor2_1
XFILLER_97_702 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13188_ _13189_/A _13189_/B _13189_/C vssd1 vssd1 vccd1 vccd1 _13188_/X sky130_fd_sc_hd__and3_1
XFILLER_151_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12139_ _12305_/A _12139_/B vssd1 vssd1 vccd1 vccd1 _12141_/B sky130_fd_sc_hd__and2_1
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16947_ _16947_/A _16947_/B vssd1 vssd1 vccd1 vccd1 _16950_/A sky130_fd_sc_hd__xnor2_1
X_16878_ _10126_/B _10014_/D _09711_/X vssd1 vssd1 vccd1 vccd1 _16878_/X sky130_fd_sc_hd__a21o_1
XFILLER_53_827 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15829_ _15932_/A _16827_/A _16514_/A _15734_/B vssd1 vssd1 vccd1 vccd1 _15829_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_52_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09350_ _09493_/A _09350_/B _14982_/B vssd1 vssd1 vccd1 vccd1 _09353_/A sky130_fd_sc_hd__and3_1
XFILLER_33_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09281_ _09281_/A _09281_/B vssd1 vssd1 vccd1 vccd1 _09289_/A sky130_fd_sc_hd__xnor2_1
XFILLER_21_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_328 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08996_ _08996_/A _08996_/B vssd1 vssd1 vccd1 vccd1 _09003_/A sky130_fd_sc_hd__nor2_1
XFILLER_125_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09617_ _09618_/B _09747_/A _09618_/A vssd1 vssd1 vccd1 vccd1 _09621_/A sky130_fd_sc_hd__a21o_1
XFILLER_141_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09548_ _09548_/A _09548_/B vssd1 vssd1 vccd1 vccd1 _09559_/A sky130_fd_sc_hd__nor2_1
XFILLER_71_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09479_ _09479_/A _09479_/B vssd1 vssd1 vccd1 vccd1 _09480_/C sky130_fd_sc_hd__xnor2_1
XFILLER_54_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11510_ _11553_/B _15042_/B _11509_/B _11506_/X vssd1 vssd1 vccd1 vccd1 _11512_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_157_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12490_ _12490_/A _12642_/A _12490_/C vssd1 vssd1 vccd1 vccd1 _12642_/B sky130_fd_sc_hd__nor3_1
XFILLER_133_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11441_ _11442_/B _11442_/A vssd1 vssd1 vccd1 vccd1 _11496_/A sky130_fd_sc_hd__nand2b_1
XFILLER_138_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14160_ _14064_/A _14066_/B _14064_/B vssd1 vssd1 vccd1 vccd1 _14161_/B sky130_fd_sc_hd__o21ba_1
X_11372_ _15373_/C _17467_/D _17466_/D _15396_/A vssd1 vssd1 vccd1 vccd1 _11373_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_138_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13111_ _13112_/A _13112_/B vssd1 vssd1 vccd1 vccd1 _13248_/A sky130_fd_sc_hd__and2b_1
XFILLER_152_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10323_ _10445_/A _10324_/B vssd1 vssd1 vccd1 vccd1 _10325_/A sky130_fd_sc_hd__nand2_1
X_14091_ _14092_/A _14092_/B _14092_/C vssd1 vssd1 vccd1 vccd1 _14200_/A sky130_fd_sc_hd__a21oi_1
XFILLER_152_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13042_ _13043_/A _13043_/B _13043_/C vssd1 vssd1 vccd1 vccd1 _13181_/B sky130_fd_sc_hd__o21ai_1
XFILLER_112_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10254_ _10254_/A _11790_/A _10920_/B _10799_/B vssd1 vssd1 vccd1 vccd1 _10257_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_133_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10185_ _10184_/A _10184_/B _10184_/C vssd1 vssd1 vccd1 vccd1 _10186_/B sky130_fd_sc_hd__o21ai_1
XFILLER_121_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16801_ _14925_/Y _15386_/B _16800_/X vssd1 vssd1 vccd1 vccd1 _16801_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_66_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout280 _08732_/X vssd1 vssd1 vccd1 vccd1 _16911_/A sky130_fd_sc_hd__buf_4
X_14993_ _15003_/B _10111_/D _09981_/D _09979_/C _09925_/A _14958_/A vssd1 vssd1 vccd1
+ vccd1 _14994_/B sky130_fd_sc_hd__mux4_1
XFILLER_75_930 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout291 _15036_/S vssd1 vssd1 vccd1 vccd1 _15056_/A sky130_fd_sc_hd__buf_4
XFILLER_75_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16732_ _14863_/B _16652_/B _16731_/Y vssd1 vssd1 vccd1 vccd1 _16732_/X sky130_fd_sc_hd__o21a_1
X_13944_ _11822_/X _14210_/B _14482_/B1 vssd1 vssd1 vccd1 vccd1 _13944_/X sky130_fd_sc_hd__o21a_1
XFILLER_47_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16663_ _16661_/X _16663_/B vssd1 vssd1 vccd1 vccd1 _16665_/A sky130_fd_sc_hd__nand2b_1
X_13875_ _13765_/A _13767_/B _13765_/B vssd1 vssd1 vccd1 vccd1 _13882_/A sky130_fd_sc_hd__o21ba_1
XFILLER_28_890 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15614_ _15614_/A _15614_/B vssd1 vssd1 vccd1 vccd1 _15615_/C sky130_fd_sc_hd__and2_1
X_12826_ _12826_/A vssd1 vssd1 vccd1 vccd1 _12826_/Y sky130_fd_sc_hd__inv_2
X_16594_ _16667_/A _16813_/B vssd1 vssd1 vccd1 vccd1 _16748_/C sky130_fd_sc_hd__nor2_1
XFILLER_61_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_90 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_988 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12757_ _12757_/A _12915_/A vssd1 vssd1 vccd1 vccd1 _12759_/B sky130_fd_sc_hd__and2_1
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15545_ _14924_/A _15457_/B _13012_/X _15536_/X _15544_/X vssd1 vssd1 vccd1 vccd1
+ _15545_/X sky130_fd_sc_hd__o311a_1
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_595 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11708_ _11708_/A _11708_/B vssd1 vssd1 vccd1 vccd1 _16105_/A sky130_fd_sc_hd__xor2_2
XFILLER_42_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15476_ _15559_/A vssd1 vssd1 vccd1 vccd1 _15476_/Y sky130_fd_sc_hd__inv_2
X_12688_ _12499_/B _12501_/B _12499_/A vssd1 vssd1 vccd1 vccd1 _12689_/C sky130_fd_sc_hd__o21ba_1
X_17215_ _17439_/Q _17245_/A2 _17213_/X _17214_/X _17275_/C1 vssd1 vssd1 vccd1 vccd1
+ _17439_/D sky130_fd_sc_hd__o221a_1
X_14427_ _14427_/A _14497_/A vssd1 vssd1 vccd1 vccd1 _14430_/A sky130_fd_sc_hd__or2_1
X_11639_ _11639_/A _11639_/B vssd1 vssd1 vccd1 vccd1 _11663_/B sky130_fd_sc_hd__xnor2_1
XFILLER_129_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14358_ _15457_/A _16735_/B _14357_/X vssd1 vssd1 vccd1 vccd1 _14358_/Y sky130_fd_sc_hd__a21oi_2
X_17146_ _16917_/A _17135_/Y _17136_/X _17145_/Y vssd1 vssd1 vccd1 vccd1 _17146_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_128_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13309_ _13309_/A _13309_/B vssd1 vssd1 vccd1 vccd1 _13312_/C sky130_fd_sc_hd__and2_1
X_17077_ _17077_/A _17077_/B _17077_/C _17076_/X vssd1 vssd1 vccd1 vccd1 _17077_/X
+ sky130_fd_sc_hd__or4b_1
X_14289_ _14708_/B _16789_/A _16722_/A _14290_/A vssd1 vssd1 vccd1 vccd1 _14291_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_171_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16028_ _16028_/A _16028_/B vssd1 vssd1 vccd1 vccd1 _16035_/A sky130_fd_sc_hd__xnor2_2
XFILLER_115_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08850_ _08996_/B _08850_/B vssd1 vssd1 vccd1 vccd1 _08907_/B sky130_fd_sc_hd__nor2_1
XFILLER_85_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08781_ _08802_/A _08802_/B vssd1 vssd1 vccd1 vccd1 _08783_/C sky130_fd_sc_hd__and2b_1
XFILLER_38_621 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09402_ _09292_/A _09291_/C _09291_/B vssd1 vssd1 vccd1 vccd1 _09437_/B sky130_fd_sc_hd__a21o_1
XFILLER_164_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09333_ _09333_/A _09333_/B vssd1 vssd1 vccd1 vccd1 _09334_/C sky130_fd_sc_hd__xnor2_1
X_09264_ _09269_/A _09269_/B vssd1 vssd1 vccd1 vccd1 _09275_/A sky130_fd_sc_hd__nor2_1
XFILLER_139_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09195_ _09196_/B _09202_/A _09196_/A vssd1 vssd1 vccd1 vccd1 _09227_/A sky130_fd_sc_hd__o21ai_1
XFILLER_147_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08979_ _17421_/A _11920_/D _08978_/C vssd1 vssd1 vccd1 vccd1 _08980_/B sky130_fd_sc_hd__a21oi_1
XFILLER_60_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11990_ _11990_/A _11990_/B _11990_/C vssd1 vssd1 vccd1 vccd1 _11991_/B sky130_fd_sc_hd__and3_1
XFILLER_28_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10941_ _10943_/A _10943_/B _10943_/C vssd1 vssd1 vccd1 vccd1 _10941_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_21_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13660_ _13662_/A _13662_/B _13662_/C vssd1 vssd1 vccd1 vccd1 _13770_/A sky130_fd_sc_hd__o21a_1
XFILLER_44_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10872_ _11124_/C _15624_/A _10854_/A _10852_/Y vssd1 vssd1 vccd1 vccd1 _10874_/C
+ sky130_fd_sc_hd__o2bb2a_1
XPHY_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12611_ _12612_/A _12612_/B _12612_/C vssd1 vssd1 vccd1 vccd1 _12611_/X sky130_fd_sc_hd__o21a_1
XFILLER_43_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13591_ _13592_/A _13592_/B vssd1 vssd1 vccd1 vccd1 _13688_/A sky130_fd_sc_hd__nor2_1
XPHY_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15330_ _15331_/A _15331_/B vssd1 vssd1 vccd1 vccd1 _15408_/A sky130_fd_sc_hd__nor2_1
X_12542_ _12372_/X _12380_/B _12696_/B _12541_/Y _15998_/A vssd1 vssd1 vccd1 vccd1
+ _12542_/Y sky130_fd_sc_hd__a311oi_2
XFILLER_61_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15261_ _16226_/C _15647_/A vssd1 vssd1 vccd1 vccd1 _15285_/A sky130_fd_sc_hd__nand2_1
XFILLER_157_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12473_ _12473_/A _12473_/B vssd1 vssd1 vccd1 vccd1 _12474_/B sky130_fd_sc_hd__xnor2_1
X_17000_ _17000_/A _17000_/B vssd1 vssd1 vccd1 vccd1 _17001_/B sky130_fd_sc_hd__nor2_1
X_14212_ _14050_/B _14213_/C _14213_/D _14213_/A vssd1 vssd1 vccd1 vccd1 _14214_/A
+ sky130_fd_sc_hd__a22oi_1
X_11424_ _11426_/B vssd1 vssd1 vccd1 vccd1 _11572_/A sky130_fd_sc_hd__inv_2
XFILLER_137_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15192_ _15901_/S _15805_/B _15190_/X vssd1 vssd1 vccd1 vccd1 _15192_/X sky130_fd_sc_hd__o21a_1
XFILLER_165_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_8 _17517_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14143_ _14676_/A _16722_/A vssd1 vssd1 vccd1 vccd1 _14145_/B sky130_fd_sc_hd__nand2_1
X_11355_ _11354_/A _11361_/A vssd1 vssd1 vccd1 vccd1 _11357_/B sky130_fd_sc_hd__nand2b_1
XFILLER_99_819 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10306_ _10182_/C _10309_/B _10183_/A _10181_/Y vssd1 vssd1 vccd1 vccd1 _10307_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_4_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14074_ _14074_/A _14074_/B vssd1 vssd1 vccd1 vccd1 _14075_/B sky130_fd_sc_hd__nand2_1
X_11286_ _11272_/Y _11311_/A _11291_/A _11256_/Y vssd1 vssd1 vccd1 vccd1 _11291_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_140_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13025_ _13156_/B _13522_/D _14065_/B _13641_/A vssd1 vssd1 vccd1 vccd1 _13027_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_112_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10237_ _10236_/B _11006_/C _11027_/D _10236_/A vssd1 vssd1 vccd1 vccd1 _10365_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_94_502 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10168_ _10045_/C _10543_/B _10162_/A _10044_/Y vssd1 vssd1 vccd1 vccd1 _10170_/C
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_120_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10099_ _10094_/A _10092_/X _09806_/A _09807_/Y vssd1 vssd1 vccd1 vccd1 _10348_/B
+ sky130_fd_sc_hd__o211a_1
X_14976_ _15846_/A _16127_/A _15278_/A _15726_/A vssd1 vssd1 vccd1 vccd1 _14977_/C
+ sky130_fd_sc_hd__a22o_1
X_16715_ _16853_/A _16853_/B vssd1 vssd1 vccd1 vccd1 _16715_/Y sky130_fd_sc_hd__nand2_1
XFILLER_35_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13927_ _13908_/A _13802_/B _13803_/A _13801_/A vssd1 vssd1 vccd1 vccd1 _13929_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_62_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16646_ _16572_/A _16574_/B _16643_/A _16644_/X vssd1 vssd1 vccd1 vccd1 _16647_/A
+ sky130_fd_sc_hd__a211o_1
X_13858_ _13858_/A _13858_/B vssd1 vssd1 vccd1 vccd1 _13859_/B sky130_fd_sc_hd__nor2_1
XFILLER_90_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12809_ _12809_/A _12809_/B vssd1 vssd1 vccd1 vccd1 _12812_/A sky130_fd_sc_hd__xnor2_1
XFILLER_62_498 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16577_ _16577_/A _16577_/B vssd1 vssd1 vccd1 vccd1 _16577_/X sky130_fd_sc_hd__xor2_1
XFILLER_31_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13789_ _14318_/A _14318_/B _14360_/D _16722_/A vssd1 vssd1 vccd1 vccd1 _13790_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_96_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15528_ _15525_/X _15526_/X _15527_/Y vssd1 vssd1 vccd1 vccd1 _15528_/Y sky130_fd_sc_hd__o21ai_1
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15459_ _11470_/A _14919_/X _15175_/A vssd1 vssd1 vccd1 vccd1 _15459_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_163_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17129_ _17130_/A _17130_/B vssd1 vssd1 vccd1 vccd1 _17131_/B sky130_fd_sc_hd__nand2_1
XFILLER_7_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_307 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09951_ _09951_/A _09951_/B _09951_/C vssd1 vssd1 vccd1 vccd1 _09952_/B sky130_fd_sc_hd__nor3_1
XFILLER_144_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08902_ _08903_/B _08903_/A vssd1 vssd1 vccd1 vccd1 _08910_/B sky130_fd_sc_hd__nand2b_1
XFILLER_106_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09882_ _09877_/X _09881_/X _09869_/X _09870_/Y vssd1 vssd1 vccd1 vccd1 _09885_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_106_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08833_ _08832_/A _08832_/Y _08800_/X _08801_/Y vssd1 vssd1 vccd1 vccd1 _08874_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_100_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08764_ _08764_/A _08764_/B vssd1 vssd1 vccd1 vccd1 _08766_/B sky130_fd_sc_hd__xor2_4
XFILLER_54_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09316_ _09316_/A _09316_/B _09316_/C vssd1 vssd1 vccd1 vccd1 _09316_/X sky130_fd_sc_hd__and3_1
XFILLER_51_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09247_ _11990_/B _09245_/Y _09152_/Y _09155_/A vssd1 vssd1 vccd1 vccd1 _09248_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_166_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09178_ _09178_/A _09178_/B _09178_/C vssd1 vssd1 vccd1 vccd1 _09179_/B sky130_fd_sc_hd__and3_1
XFILLER_119_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11140_ _11128_/Y _11255_/A _11146_/A _11113_/Y vssd1 vssd1 vccd1 vccd1 _11146_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_116_990 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput78 _17471_/Q vssd1 vssd1 vccd1 vccd1 leds[5] sky130_fd_sc_hd__clkbuf_1
X_11071_ _11065_/A _11065_/C _11065_/D _11065_/B vssd1 vssd1 vccd1 vccd1 _11071_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_0_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput89 _17448_/Q vssd1 vssd1 vccd1 vccd1 o_wb_data[14] sky130_fd_sc_hd__clkbuf_1
XFILLER_163_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10022_ _10136_/A _10136_/B vssd1 vssd1 vccd1 vccd1 _10023_/C sky130_fd_sc_hd__nand2_1
XFILLER_103_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14830_ _14597_/B _14828_/Y _14829_/X _17167_/A vssd1 vssd1 vccd1 vccd1 _17167_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_48_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11973_ _08993_/C _08992_/Y _08965_/Y vssd1 vssd1 vccd1 vccd1 _11986_/B sky130_fd_sc_hd__a21o_1
X_14761_ _14738_/A _14738_/B _14739_/Y _14748_/A _14760_/Y vssd1 vssd1 vccd1 vccd1
+ _14762_/B sky130_fd_sc_hd__a311o_1
XFILLER_91_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16500_ _16747_/A _16499_/B _16499_/C vssd1 vssd1 vccd1 vccd1 _16501_/B sky130_fd_sc_hd__o21ai_1
X_10924_ _10924_/A _10924_/B vssd1 vssd1 vccd1 vccd1 _10926_/B sky130_fd_sc_hd__xnor2_2
X_13712_ _13605_/A _13605_/B _13562_/A vssd1 vssd1 vccd1 vccd1 _13713_/C sky130_fd_sc_hd__a21oi_1
XFILLER_45_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17480_ fanout949/X _17480_/D vssd1 vssd1 vccd1 vccd1 _17480_/Q sky130_fd_sc_hd__dfxtp_4
X_14692_ _14723_/A _14692_/B vssd1 vssd1 vccd1 vccd1 _14693_/C sky130_fd_sc_hd__nor2_1
XFILLER_60_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16431_ _16431_/A _16511_/A vssd1 vssd1 vccd1 vccd1 _16432_/C sky130_fd_sc_hd__nor2_1
XFILLER_147_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_796 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10855_ _10855_/A _10855_/B vssd1 vssd1 vccd1 vccd1 _10865_/B sky130_fd_sc_hd__xnor2_1
X_13643_ _13643_/A _13852_/B vssd1 vssd1 vccd1 vccd1 _13644_/B sky130_fd_sc_hd__nand2_1
XFILLER_72_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16362_ _16362_/A _16362_/B vssd1 vssd1 vccd1 vccd1 _16364_/B sky130_fd_sc_hd__xnor2_1
X_13574_ _13702_/B _13574_/B vssd1 vssd1 vccd1 vccd1 _13576_/C sky130_fd_sc_hd__nand2_1
XFILLER_72_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10786_ _10991_/A _10786_/B _10991_/C vssd1 vssd1 vccd1 vccd1 _10901_/A sky130_fd_sc_hd__and3_1
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12525_ _12526_/A _12526_/B _12526_/C vssd1 vssd1 vccd1 vccd1 _12528_/A sky130_fd_sc_hd__a21oi_2
X_15313_ _12858_/Y _16011_/C _15312_/X _16011_/A vssd1 vssd1 vccd1 vccd1 _15313_/Y
+ sky130_fd_sc_hd__o22ai_2
XFILLER_157_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16293_ _16293_/A _16293_/B vssd1 vssd1 vccd1 vccd1 _16293_/Y sky130_fd_sc_hd__xnor2_4
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15244_ _15244_/A _15244_/B _15244_/C vssd1 vssd1 vccd1 vccd1 _15244_/X sky130_fd_sc_hd__or3_1
X_12456_ _12626_/A _12454_/Y _12280_/X _12284_/A vssd1 vssd1 vccd1 vccd1 _12458_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_8_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11407_ _11402_/A _11402_/B _11451_/A vssd1 vssd1 vccd1 vccd1 _11408_/C sky130_fd_sc_hd__o21ba_1
XFILLER_126_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15175_ _15175_/A _15175_/B _15450_/B vssd1 vssd1 vccd1 vccd1 _15175_/X sky130_fd_sc_hd__or3_1
XFILLER_126_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12387_ _12385_/X _12386_/X _12865_/S vssd1 vssd1 vccd1 vccd1 _12387_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_702 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14126_ _14763_/S _14124_/Y _14205_/B _14038_/Y vssd1 vssd1 vccd1 vccd1 _17593_/D
+ sky130_fd_sc_hd__a31o_1
X_11338_ _11386_/A _11337_/B _11337_/A vssd1 vssd1 vccd1 vccd1 _11340_/B sky130_fd_sc_hd__o21ba_1
XFILLER_126_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_595 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14057_ _14057_/A _14057_/B vssd1 vssd1 vccd1 vccd1 _14060_/A sky130_fd_sc_hd__xor2_1
XFILLER_113_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11269_ _11553_/A _11518_/C _15244_/A _11320_/A vssd1 vssd1 vccd1 vccd1 _11313_/A
+ sky130_fd_sc_hd__a31o_1
X_13008_ _11781_/B _12377_/Y _13005_/B _13005_/X _13007_/Y vssd1 vssd1 vccd1 vccd1
+ _13010_/B sky130_fd_sc_hd__a311o_2
XFILLER_97_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14959_ _14954_/A _14956_/Y _14958_/Y _15097_/A vssd1 vssd1 vccd1 vccd1 _14959_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_47_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16629_ _16630_/A _16630_/B _16630_/C vssd1 vssd1 vccd1 vccd1 _16711_/A sky130_fd_sc_hd__a21oi_1
XFILLER_35_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09101_ _09101_/A _09165_/A vssd1 vssd1 vccd1 vccd1 _09103_/B sky130_fd_sc_hd__nor2_1
XFILLER_149_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09032_ _17081_/A _09032_/B vssd1 vssd1 vccd1 vccd1 _09262_/A sky130_fd_sc_hd__xnor2_1
XFILLER_129_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_551 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_26 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout802 _10525_/D vssd1 vssd1 vccd1 vccd1 _10933_/D sky130_fd_sc_hd__buf_2
XFILLER_132_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09934_ _10075_/A _09935_/B vssd1 vssd1 vccd1 vccd1 _09936_/A sky130_fd_sc_hd__nor2_1
Xfanout813 _10508_/D vssd1 vssd1 vccd1 vccd1 _10970_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_120_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout824 _17487_/Q vssd1 vssd1 vccd1 vccd1 _09265_/C sky130_fd_sc_hd__buf_6
XFILLER_58_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout835 _09409_/D vssd1 vssd1 vccd1 vccd1 _09843_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_131_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout846 _17484_/Q vssd1 vssd1 vccd1 vccd1 _12463_/D sky130_fd_sc_hd__buf_4
X_09865_ _09865_/A _09865_/B vssd1 vssd1 vccd1 vccd1 _09884_/B sky130_fd_sc_hd__nand2_1
Xfanout857 _15238_/A vssd1 vssd1 vccd1 vccd1 _14906_/B sky130_fd_sc_hd__clkbuf_4
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout868 _15151_/B vssd1 vssd1 vccd1 vccd1 _15175_/B sky130_fd_sc_hd__buf_2
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout879 _15110_/A vssd1 vssd1 vccd1 vccd1 _15116_/B sky130_fd_sc_hd__buf_2
XFILLER_133_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08816_ _08876_/A _08876_/B vssd1 vssd1 vccd1 vccd1 _08831_/C sky130_fd_sc_hd__and2_1
XTAP_3206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09796_ _14770_/A _15003_/B vssd1 vssd1 vccd1 vccd1 _10062_/C sky130_fd_sc_hd__and2_1
XFILLER_100_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08747_ _08747_/A vssd1 vssd1 vccd1 vccd1 _08748_/B sky130_fd_sc_hd__clkinv_2
XFILLER_100_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10640_ _10641_/A _10639_/Y _11117_/C _10743_/D vssd1 vssd1 vccd1 vccd1 _10724_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_167_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10571_ _10571_/A _10571_/B vssd1 vssd1 vccd1 vccd1 _10586_/B sky130_fd_sc_hd__xnor2_1
XFILLER_139_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12310_ _12310_/A _12310_/B vssd1 vssd1 vccd1 vccd1 _12311_/B sky130_fd_sc_hd__nor2_1
XFILLER_10_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13290_ _13417_/B _13290_/B vssd1 vssd1 vccd1 vccd1 _13292_/B sky130_fd_sc_hd__nor2_1
XFILLER_10_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12241_ _12241_/A _12241_/B vssd1 vssd1 vccd1 vccd1 _12250_/A sky130_fd_sc_hd__xor2_1
XFILLER_108_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12172_ _12172_/A _12172_/B vssd1 vssd1 vccd1 vccd1 _12188_/A sky130_fd_sc_hd__xnor2_1
XFILLER_150_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11123_ _11122_/B _14850_/A _11518_/C _11122_/A vssd1 vssd1 vccd1 vccd1 _11123_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_123_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16980_ _17156_/B _16969_/Y _16979_/X _16963_/X vssd1 vssd1 vccd1 vccd1 _16980_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_1_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15931_ _16138_/A _16827_/B vssd1 vssd1 vccd1 vccd1 _16040_/A sky130_fd_sc_hd__nor2_1
X_11054_ _11041_/Y _11042_/X _11047_/Y _11050_/X vssd1 vssd1 vccd1 vccd1 _11055_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_49_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10005_ _10005_/A _10005_/B _10005_/C vssd1 vssd1 vccd1 vccd1 _10005_/X sky130_fd_sc_hd__and3_1
XFILLER_114_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15862_ _15863_/B _15863_/A vssd1 vssd1 vccd1 vccd1 _15980_/B sky130_fd_sc_hd__and2b_1
XFILLER_76_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17601_ fanout933/X _17601_/D vssd1 vssd1 vccd1 vccd1 _17601_/Q sky130_fd_sc_hd__dfxtp_1
X_14813_ _16112_/B _16112_/C _16315_/A vssd1 vssd1 vccd1 vccd1 _14813_/X sky130_fd_sc_hd__a21bo_1
XFILLER_18_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15793_ _15793_/A _15793_/B vssd1 vssd1 vccd1 vccd1 _15794_/B sky130_fd_sc_hd__nor2_1
XFILLER_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17532_ fanout944/X _17532_/D vssd1 vssd1 vccd1 vccd1 _17532_/Q sky130_fd_sc_hd__dfxtp_1
X_14744_ _14744_/A _14744_/B vssd1 vssd1 vccd1 vccd1 _14745_/B sky130_fd_sc_hd__nand2_1
X_11956_ _11956_/A _12163_/A _11956_/C vssd1 vssd1 vccd1 vccd1 _12163_/B sky130_fd_sc_hd__nor3_1
XFILLER_44_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10907_ _10907_/A _10907_/B vssd1 vssd1 vccd1 vccd1 _10909_/A sky130_fd_sc_hd__nor2_1
X_17463_ fanout953/X _17463_/D vssd1 vssd1 vccd1 vccd1 _17463_/Q sky130_fd_sc_hd__dfxtp_2
X_11887_ _11888_/A _11888_/B vssd1 vssd1 vccd1 vccd1 _12118_/B sky130_fd_sc_hd__nand2_1
XFILLER_72_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14675_ _14675_/A _17167_/A vssd1 vssd1 vccd1 vccd1 _14677_/A sky130_fd_sc_hd__xnor2_1
XFILLER_60_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16414_ _16414_/A _16414_/B vssd1 vssd1 vccd1 vccd1 _16422_/A sky130_fd_sc_hd__xor2_1
X_10838_ _11124_/C _10933_/C vssd1 vssd1 vccd1 vccd1 _10842_/A sky130_fd_sc_hd__nand2_1
X_13626_ _14421_/S _13626_/B vssd1 vssd1 vccd1 vccd1 _13841_/A sky130_fd_sc_hd__nand2_1
X_17394_ input42/X _17426_/A2 _17393_/X _17408_/C1 vssd1 vssd1 vccd1 vccd1 _17525_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_41_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16345_ _16345_/A _16345_/B vssd1 vssd1 vccd1 vccd1 _16345_/X sky130_fd_sc_hd__or2_1
XFILLER_157_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1046 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10769_ _10769_/A _10769_/B vssd1 vssd1 vccd1 vccd1 _10771_/C sky130_fd_sc_hd__and2_1
X_13557_ _13558_/A _13558_/B _13558_/C vssd1 vssd1 vccd1 vccd1 _13557_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_158_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12508_ _12508_/A _12508_/B _12508_/C vssd1 vssd1 vccd1 vccd1 _12509_/B sky130_fd_sc_hd__nor3_1
X_16276_ _16276_/A _16276_/B vssd1 vssd1 vccd1 vccd1 _16277_/B sky130_fd_sc_hd__nand2_1
X_13488_ _13365_/Y _13369_/B _13486_/X _13487_/Y vssd1 vssd1 vccd1 vccd1 _13490_/C
+ sky130_fd_sc_hd__a211oi_2
XFILLER_145_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12439_ _12592_/A _12592_/B _12592_/D _12439_/D vssd1 vssd1 vccd1 vccd1 _12616_/A
+ sky130_fd_sc_hd__and4_1
X_15227_ _15166_/A _15166_/B _15162_/A vssd1 vssd1 vccd1 vccd1 _15228_/B sky130_fd_sc_hd__o21a_1
XFILLER_154_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15158_ _15159_/A _15159_/B vssd1 vssd1 vccd1 vccd1 _15221_/A sky130_fd_sc_hd__nand2_1
XFILLER_99_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14109_ _14013_/A _14013_/B _14013_/C _14110_/B vssd1 vssd1 vccd1 vccd1 _14197_/B
+ sky130_fd_sc_hd__a211o_1
X_15089_ _16086_/A _15088_/Y _15089_/S vssd1 vssd1 vccd1 vccd1 _15091_/B sky130_fd_sc_hd__mux2_1
XFILLER_68_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09650_ _09654_/C _12025_/B _09619_/B _09494_/Y vssd1 vssd1 vccd1 vccd1 _09656_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_55_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09581_ _09581_/A _09581_/B _09581_/C vssd1 vssd1 vccd1 vccd1 _09581_/Y sky130_fd_sc_hd__nand3_1
XFILLER_83_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_805 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09015_ _09016_/A _09016_/B _09016_/C vssd1 vssd1 vccd1 vccd1 _09015_/X sky130_fd_sc_hd__and3_1
XFILLER_152_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout610 _17510_/Q vssd1 vssd1 vccd1 vccd1 _15058_/S0 sky130_fd_sc_hd__buf_2
XFILLER_59_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout621 _11932_/B vssd1 vssd1 vccd1 vccd1 _12592_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_120_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout632 _14094_/B vssd1 vssd1 vccd1 vccd1 _13846_/B sky130_fd_sc_hd__buf_2
X_09917_ _09915_/A _10059_/A _09770_/Y _09830_/X vssd1 vssd1 vccd1 vccd1 _09960_/A
+ sky130_fd_sc_hd__o211ai_4
Xfanout643 _14765_/B vssd1 vssd1 vccd1 vccd1 _13035_/C sky130_fd_sc_hd__buf_2
Xfanout654 _17505_/Q vssd1 vssd1 vccd1 vccd1 _17028_/A sky130_fd_sc_hd__clkbuf_4
Xfanout665 _17504_/Q vssd1 vssd1 vccd1 vccd1 _12025_/B sky130_fd_sc_hd__buf_4
Xfanout676 _16859_/A vssd1 vssd1 vccd1 vccd1 _14426_/D sky130_fd_sc_hd__clkbuf_4
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout687 fanout690/X vssd1 vssd1 vccd1 vccd1 _12256_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_85_140 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09848_ _09848_/A _09848_/B vssd1 vssd1 vccd1 vccd1 _09976_/B sky130_fd_sc_hd__xnor2_1
XFILLER_58_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout698 fanout699/X vssd1 vssd1 vccd1 vccd1 _10309_/B sky130_fd_sc_hd__buf_2
XTAP_3003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09779_ _09925_/A _14863_/A vssd1 vssd1 vccd1 vccd1 _14952_/A sky130_fd_sc_hd__and2_1
XTAP_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11810_ _11807_/Y _11809_/Y _12212_/S vssd1 vssd1 vccd1 vccd1 _11810_/X sky130_fd_sc_hd__mux2_1
XTAP_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12790_ _12790_/A _12947_/A _12790_/C vssd1 vssd1 vccd1 vccd1 _12947_/B sky130_fd_sc_hd__nor3_1
XTAP_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11741_ _10778_/A _10777_/C _10777_/A vssd1 vssd1 vccd1 vccd1 _11742_/B sky130_fd_sc_hd__o21a_1
XFILLER_57_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11672_ _11672_/A _11672_/B _11672_/C vssd1 vssd1 vccd1 vccd1 _11672_/Y sky130_fd_sc_hd__nand3_1
XTAP_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14460_ _14518_/A _14459_/B _14459_/C vssd1 vssd1 vccd1 vccd1 _14460_/X sky130_fd_sc_hd__a21o_1
XFILLER_144_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10623_ _10624_/B _10624_/A vssd1 vssd1 vccd1 vccd1 _10623_/X sky130_fd_sc_hd__and2b_1
X_13411_ _13411_/A _13411_/B _13411_/C vssd1 vssd1 vccd1 vccd1 _13423_/B sky130_fd_sc_hd__nand3_1
X_14391_ _14393_/A _14393_/B _14393_/C vssd1 vssd1 vccd1 vccd1 _14394_/A sky130_fd_sc_hd__a21oi_1
XFILLER_128_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16130_ _16130_/A _16130_/B vssd1 vssd1 vccd1 vccd1 _16133_/A sky130_fd_sc_hd__xor2_1
XFILLER_139_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13342_ _16723_/A _13564_/C _13342_/C vssd1 vssd1 vccd1 vccd1 _13462_/B sky130_fd_sc_hd__nand3_1
XFILLER_167_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10554_ _10406_/B _10474_/Y _10519_/A _10519_/Y vssd1 vssd1 vccd1 vccd1 _10555_/C
+ sky130_fd_sc_hd__a211oi_1
XFILLER_6_612 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16061_ _16352_/A _16061_/B vssd1 vssd1 vccd1 vccd1 _16168_/C sky130_fd_sc_hd__nand2_1
XFILLER_143_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13273_ _13831_/S _12222_/X _12229_/C _12858_/Y vssd1 vssd1 vccd1 vccd1 _13273_/X
+ sky130_fd_sc_hd__o22a_2
X_10485_ _10497_/A _10497_/B vssd1 vssd1 vccd1 vccd1 _10485_/X sky130_fd_sc_hd__or2_1
XFILLER_136_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15012_ _14796_/C _16008_/A2 _15009_/X _15011_/X _14944_/A vssd1 vssd1 vccd1 vccd1
+ _15012_/X sky130_fd_sc_hd__a2111o_1
XFILLER_6_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12224_ _11802_/Y _11842_/Y _12700_/B vssd1 vssd1 vccd1 vccd1 _12224_/X sky130_fd_sc_hd__mux2_1
XFILLER_136_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12155_ _12155_/A _12155_/B vssd1 vssd1 vccd1 vccd1 _12192_/A sky130_fd_sc_hd__nor2_1
XFILLER_151_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11106_ _11005_/A _17467_/D _17466_/D _10904_/A vssd1 vssd1 vccd1 vccd1 _11107_/B
+ sky130_fd_sc_hd__a22oi_1
XFILLER_151_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16963_ _16931_/X _16932_/X _16960_/X _16962_/Y vssd1 vssd1 vccd1 vccd1 _16963_/X
+ sky130_fd_sc_hd__a31o_2
X_12086_ _11882_/A _11884_/B _11882_/B vssd1 vssd1 vccd1 vccd1 _12096_/A sky130_fd_sc_hd__o21ba_1
X_11037_ _11038_/A _11038_/B vssd1 vssd1 vccd1 vccd1 _11181_/A sky130_fd_sc_hd__and2b_1
X_15914_ _16315_/B _15658_/Y _16813_/B _15820_/A vssd1 vssd1 vccd1 vccd1 _15915_/B
+ sky130_fd_sc_hd__o22a_1
X_16894_ _16895_/A _16895_/B vssd1 vssd1 vccd1 vccd1 _16952_/B sky130_fd_sc_hd__or2_1
XFILLER_37_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15845_ _16055_/A _16681_/D vssd1 vssd1 vccd1 vccd1 _16268_/A sky130_fd_sc_hd__or2_1
XFILLER_37_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_143 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15776_ _15877_/A _15776_/B _15776_/C vssd1 vssd1 vccd1 vccd1 _15877_/B sky130_fd_sc_hd__nor3_1
XTAP_3581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12988_ _13125_/B _12986_/Y _12825_/A _12826_/Y vssd1 vssd1 vccd1 vccd1 _12988_/Y
+ sky130_fd_sc_hd__a211oi_1
XFILLER_91_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17515_ fanout942/X _17515_/D vssd1 vssd1 vccd1 vccd1 _17515_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14727_ _14727_/A _14727_/B vssd1 vssd1 vccd1 vccd1 _14728_/B sky130_fd_sc_hd__or2_1
XFILLER_91_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11939_ _11939_/A _11939_/B vssd1 vssd1 vccd1 vccd1 _11941_/B sky130_fd_sc_hd__xor2_1
XTAP_2880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17446_ fanout940/X _17446_/D vssd1 vssd1 vccd1 vccd1 _17446_/Q sky130_fd_sc_hd__dfxtp_1
X_14658_ _14658_/A _14658_/B _14658_/C vssd1 vssd1 vccd1 vccd1 _14659_/B sky130_fd_sc_hd__or3_1
XFILLER_20_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13609_ _13718_/A _13607_/X _13486_/X _13490_/C vssd1 vssd1 vccd1 vccd1 _13609_/X
+ sky130_fd_sc_hd__a211o_1
X_17377_ _17377_/A _17377_/B vssd1 vssd1 vccd1 vccd1 _17377_/Y sky130_fd_sc_hd__nand2_1
XFILLER_158_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14589_ _13142_/X _13145_/B _14757_/S vssd1 vssd1 vccd1 vccd1 _14590_/B sky130_fd_sc_hd__mux2_1
XFILLER_174_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16328_ _16328_/A _16328_/B vssd1 vssd1 vccd1 vccd1 _16425_/B sky130_fd_sc_hd__nor2_1
XFILLER_146_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16259_ _16352_/A _16259_/B _16259_/C vssd1 vssd1 vccd1 vccd1 _16358_/A sky130_fd_sc_hd__and3_1
XFILLER_146_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_298 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09702_ _09702_/A _09706_/B vssd1 vssd1 vccd1 vccd1 _09835_/A sky130_fd_sc_hd__nor2_1
XFILLER_114_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09633_ _10560_/A _09843_/D _09520_/C vssd1 vssd1 vccd1 vccd1 _09634_/B sky130_fd_sc_hd__a21oi_1
XFILLER_110_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09564_ _09565_/A _09565_/B vssd1 vssd1 vccd1 vccd1 _09581_/A sky130_fd_sc_hd__nand2b_1
XFILLER_43_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09495_ _09619_/B _09494_/Y _09654_/C _12025_/B vssd1 vssd1 vccd1 vccd1 _09656_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_24_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1030 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10270_ _14784_/A _10270_/B vssd1 vssd1 vccd1 vccd1 _15622_/A sky130_fd_sc_hd__nand2_1
XFILLER_3_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout440 _12722_/B vssd1 vssd1 vccd1 vccd1 _13156_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_94_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout451 _09412_/A vssd1 vssd1 vccd1 vccd1 _16108_/C sky130_fd_sc_hd__buf_2
Xfanout462 _11006_/A vssd1 vssd1 vccd1 vccd1 _10954_/A sky130_fd_sc_hd__clkbuf_4
X_13960_ _13961_/A _13961_/B _13961_/C vssd1 vssd1 vccd1 vccd1 _14047_/A sky130_fd_sc_hd__o21ai_1
XFILLER_48_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout473 _17523_/Q vssd1 vssd1 vccd1 vccd1 _11790_/A sky130_fd_sc_hd__buf_4
XFILLER_19_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout484 _17521_/Q vssd1 vssd1 vccd1 vccd1 _09873_/A sky130_fd_sc_hd__buf_4
XFILLER_74_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout495 _15262_/B vssd1 vssd1 vccd1 vccd1 _14784_/A sky130_fd_sc_hd__buf_4
X_12911_ _13060_/A _12911_/B vssd1 vssd1 vccd1 vccd1 _12913_/B sky130_fd_sc_hd__and2_1
X_13891_ _13891_/A _13891_/B vssd1 vssd1 vccd1 vccd1 _13892_/B sky130_fd_sc_hd__or2_1
XTAP_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15630_ _15175_/A _15629_/X _15808_/A vssd1 vssd1 vccd1 vccd1 _15630_/X sky130_fd_sc_hd__a21o_1
X_12842_ _13003_/B _12842_/B vssd1 vssd1 vccd1 vccd1 _12843_/B sky130_fd_sc_hd__xnor2_1
XFILLER_73_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15561_ _15655_/A _15655_/B vssd1 vssd1 vccd1 vccd1 _15656_/A sky130_fd_sc_hd__nand2_1
X_12773_ _12773_/A _12773_/B vssd1 vssd1 vccd1 vccd1 _12775_/B sky130_fd_sc_hd__xnor2_1
XTAP_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17300_ _15003_/B _17322_/A2 _17299_/X _17378_/C1 vssd1 vssd1 vccd1 vccd1 _17479_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_70_850 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14512_ _14512_/A _14512_/B vssd1 vssd1 vccd1 vccd1 _14514_/B sky130_fd_sc_hd__nor2_1
XTAP_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11724_ _11217_/A _11215_/Y _11214_/Y vssd1 vssd1 vccd1 vccd1 _11725_/C sky130_fd_sc_hd__o21ai_1
XTAP_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15492_ _16315_/D _15492_/B vssd1 vssd1 vccd1 vccd1 _16334_/C sky130_fd_sc_hd__or2_1
XTAP_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17231_ _17586_/Q _17273_/A2 _17273_/B1 vssd1 vssd1 vccd1 vccd1 _17231_/X sky130_fd_sc_hd__a21o_1
X_11655_ _11655_/A _11676_/A vssd1 vssd1 vccd1 vccd1 _11657_/C sky130_fd_sc_hd__and2_1
X_14443_ _14443_/A _14443_/B vssd1 vssd1 vccd1 vccd1 _14445_/C sky130_fd_sc_hd__xor2_1
XFILLER_30_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10606_ _10904_/A _10703_/B _11005_/B _11006_/A vssd1 vssd1 vccd1 vccd1 _10607_/B
+ sky130_fd_sc_hd__a22oi_1
XFILLER_80_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17162_ _17151_/B _17162_/A2 _16974_/B _17153_/A _17162_/C1 vssd1 vssd1 vccd1 vccd1
+ _17162_/X sky130_fd_sc_hd__a221o_1
X_11586_ _11586_/A _11586_/B _11586_/C vssd1 vssd1 vccd1 vccd1 _11700_/A sky130_fd_sc_hd__nand3_1
XFILLER_11_983 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14374_ _14302_/A _14304_/B _14302_/B vssd1 vssd1 vccd1 vccd1 _14376_/B sky130_fd_sc_hd__o21ba_1
XFILLER_167_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16113_ _16315_/A _16112_/B _16112_/C vssd1 vssd1 vccd1 vccd1 _16113_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_155_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10537_ _10637_/A _10637_/B vssd1 vssd1 vccd1 vccd1 _10540_/C sky130_fd_sc_hd__nand2_1
X_13325_ _13326_/A _13326_/B _13326_/C vssd1 vssd1 vccd1 vccd1 _13486_/A sky130_fd_sc_hd__o21a_1
X_17093_ _17093_/A _17093_/B _17093_/C vssd1 vssd1 vccd1 vccd1 _17093_/Y sky130_fd_sc_hd__nor3_1
XFILLER_170_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16044_ _16044_/A _16044_/B vssd1 vssd1 vccd1 vccd1 _16046_/B sky130_fd_sc_hd__xor2_1
X_13256_ _13256_/A _13256_/B vssd1 vssd1 vccd1 vccd1 _13258_/C sky130_fd_sc_hd__and2_1
X_10468_ _10581_/A _10581_/B _10581_/C vssd1 vssd1 vccd1 vccd1 _11771_/A sky130_fd_sc_hd__o21ai_1
XFILLER_108_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12207_ _12371_/B _12206_/B _12206_/C vssd1 vssd1 vccd1 vccd1 _12208_/B sky130_fd_sc_hd__o21a_1
X_13187_ _13326_/B _13187_/B vssd1 vssd1 vccd1 vccd1 _13189_/C sky130_fd_sc_hd__nor2_1
XFILLER_9_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10399_ _10399_/A _10399_/B vssd1 vssd1 vccd1 vccd1 _10501_/B sky130_fd_sc_hd__nor2_1
X_12138_ _12138_/A _12138_/B _12138_/C vssd1 vssd1 vccd1 vccd1 _12139_/B sky130_fd_sc_hd__or3_1
XFILLER_69_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16946_ _16947_/A _16947_/B vssd1 vssd1 vccd1 vccd1 _17003_/A sky130_fd_sc_hd__nand2b_1
X_12069_ _12239_/A vssd1 vssd1 vccd1 vccd1 _12070_/D sky130_fd_sc_hd__inv_2
XFILLER_84_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16877_ _16931_/A _16931_/B _16851_/A vssd1 vssd1 vccd1 vccd1 _16910_/A sky130_fd_sc_hd__o21ai_1
XFILLER_49_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15828_ _15737_/A _15737_/B _15735_/B vssd1 vssd1 vccd1 vccd1 _15836_/A sky130_fd_sc_hd__o21ai_2
XFILLER_53_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15759_ _15759_/A _15759_/B vssd1 vssd1 vccd1 vccd1 _15760_/B sky130_fd_sc_hd__xnor2_1
XFILLER_127_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09280_ _09281_/A _09281_/B vssd1 vssd1 vccd1 vccd1 _09296_/A sky130_fd_sc_hd__nand2b_1
XFILLER_100_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17429_ input70/X _17429_/B _17429_/C vssd1 vssd1 vccd1 vccd1 _17433_/S sky130_fd_sc_hd__or3_4
XFILLER_159_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08995_ _09327_/C _11815_/B _08943_/A _08941_/B vssd1 vssd1 vccd1 vccd1 _09004_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_76_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09616_ _09618_/B _09747_/A _09618_/A vssd1 vssd1 vccd1 vccd1 _09616_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_44_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09547_ _10366_/A _09409_/D _09410_/A _09408_/Y vssd1 vssd1 vccd1 vccd1 _09548_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_43_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09478_ _09478_/A _09478_/B _09603_/A vssd1 vssd1 vccd1 vccd1 _09480_/B sky130_fd_sc_hd__nand3_1
XFILLER_34_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11440_ _11440_/A _11479_/A vssd1 vssd1 vccd1 vccd1 _11442_/B sky130_fd_sc_hd__nor2_1
XFILLER_149_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11371_ _11423_/B _11592_/B vssd1 vssd1 vccd1 vccd1 _11529_/A sky130_fd_sc_hd__nand2_1
XFILLER_125_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13110_ _13241_/A _13110_/B vssd1 vssd1 vccd1 vccd1 _13112_/B sky130_fd_sc_hd__and2_1
X_10322_ _10322_/A _10322_/B vssd1 vssd1 vccd1 vccd1 _10324_/B sky130_fd_sc_hd__xnor2_1
XFILLER_3_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14090_ _14090_/A _14090_/B vssd1 vssd1 vccd1 vccd1 _14092_/C sky130_fd_sc_hd__xnor2_1
XFILLER_166_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13041_ _13181_/A _13041_/B vssd1 vssd1 vccd1 vccd1 _13043_/C sky130_fd_sc_hd__and2_1
XFILLER_152_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10253_ _10253_/A _10253_/B vssd1 vssd1 vccd1 vccd1 _10260_/A sky130_fd_sc_hd__xnor2_1
XFILLER_121_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10184_ _10184_/A _10184_/B _10184_/C vssd1 vssd1 vccd1 vccd1 _10331_/A sky130_fd_sc_hd__or3_1
X_16800_ _12788_/A _14863_/A _17075_/A2 _16799_/X vssd1 vssd1 vccd1 vccd1 _16800_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_121_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14992_ _15102_/A _14992_/B vssd1 vssd1 vccd1 vccd1 _14992_/Y sky130_fd_sc_hd__nand2_1
XFILLER_47_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout270 _14940_/X vssd1 vssd1 vccd1 vccd1 _17153_/B sky130_fd_sc_hd__buf_2
Xfanout281 _11653_/B vssd1 vssd1 vccd1 vccd1 _11675_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_19_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_398 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout292 fanout299/X vssd1 vssd1 vccd1 vccd1 _17367_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_87_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16731_ _14863_/B _16652_/B _16731_/B1 vssd1 vssd1 vccd1 vccd1 _16731_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_47_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13943_ _11844_/X _11854_/X _14356_/S vssd1 vssd1 vccd1 vccd1 _13943_/X sky130_fd_sc_hd__mux2_1
XFILLER_75_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16662_ _16747_/A _16938_/B _16662_/C _16662_/D vssd1 vssd1 vccd1 vccd1 _16663_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_47_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13874_ _14018_/A _13874_/B vssd1 vssd1 vccd1 vccd1 _13918_/A sky130_fd_sc_hd__and2_1
XFILLER_34_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15613_ _15610_/Y _15611_/X _15612_/X vssd1 vssd1 vccd1 vccd1 _15613_/Y sky130_fd_sc_hd__a21boi_2
X_12825_ _12825_/A _12825_/B _12825_/C vssd1 vssd1 vccd1 vccd1 _12826_/A sky130_fd_sc_hd__or3_1
X_16593_ _16686_/B _16593_/B vssd1 vssd1 vccd1 vccd1 _16597_/A sky130_fd_sc_hd__nor2_1
XFILLER_15_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15544_ _16015_/A _15624_/B _15541_/Y _15543_/X _15540_/X vssd1 vssd1 vccd1 vccd1
+ _15544_/X sky130_fd_sc_hd__o311a_1
X_12756_ _12755_/A _12755_/B _12755_/C vssd1 vssd1 vccd1 vccd1 _12915_/A sky130_fd_sc_hd__o21ai_1
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11707_ _15997_/A _15997_/B vssd1 vssd1 vccd1 vccd1 _11707_/Y sky130_fd_sc_hd__nand2_1
XFILLER_30_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15475_ _15475_/A _16127_/A _16152_/A _16604_/B vssd1 vssd1 vccd1 vccd1 _15559_/A
+ sky130_fd_sc_hd__and4_1
X_12687_ _12684_/X _12685_/Y _12528_/A _12530_/A vssd1 vssd1 vccd1 vccd1 _12689_/B
+ sky130_fd_sc_hd__a211oi_1
X_17214_ _17548_/Q _17244_/B vssd1 vssd1 vccd1 vccd1 _17214_/X sky130_fd_sc_hd__and2_1
X_14426_ _14641_/A _14641_/B _14865_/B _14426_/D vssd1 vssd1 vccd1 vccd1 _14497_/A
+ sky130_fd_sc_hd__and4_1
X_11638_ _11659_/A _11659_/B vssd1 vssd1 vccd1 vccd1 _11663_/A sky130_fd_sc_hd__nand2_1
XFILLER_128_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17145_ _17070_/B _17138_/Y _17144_/X vssd1 vssd1 vccd1 vccd1 _17145_/Y sky130_fd_sc_hd__o21ai_1
X_14357_ _12703_/X _14210_/B _14482_/B1 vssd1 vssd1 vccd1 vccd1 _14357_/X sky130_fd_sc_hd__o21a_1
XFILLER_144_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11569_ _11557_/X _11603_/A _11526_/B _11552_/X vssd1 vssd1 vccd1 vccd1 _11576_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_156_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_424 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13308_ _13308_/A _13308_/B _13308_/C vssd1 vssd1 vccd1 vccd1 _13309_/B sky130_fd_sc_hd__nand3_1
XFILLER_6_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17076_ _17112_/A1 _17164_/C _15180_/X _16735_/A _14667_/B vssd1 vssd1 vccd1 vccd1
+ _17076_/X sky130_fd_sc_hd__o32a_1
XFILLER_144_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14288_ _14734_/A _16653_/B _14287_/X vssd1 vssd1 vccd1 vccd1 _14288_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_171_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16027_ _16028_/A _16028_/B vssd1 vssd1 vccd1 vccd1 _16027_/Y sky130_fd_sc_hd__nand2_1
X_13239_ _13366_/A _13239_/B vssd1 vssd1 vccd1 vccd1 _13241_/B sky130_fd_sc_hd__and2_1
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08780_ _08780_/A _08780_/B vssd1 vssd1 vccd1 vccd1 _08802_/B sky130_fd_sc_hd__xnor2_1
XFILLER_111_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16929_ _16304_/A _16918_/X _16919_/Y _16922_/Y _16928_/X vssd1 vssd1 vccd1 vccd1
+ _16929_/X sky130_fd_sc_hd__o311a_1
XFILLER_37_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09401_ _09401_/A _09401_/B vssd1 vssd1 vccd1 vccd1 _09483_/A sky130_fd_sc_hd__nor2_1
XFILLER_53_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09332_ _09332_/A _09332_/B _09463_/A vssd1 vssd1 vccd1 vccd1 _09334_/B sky130_fd_sc_hd__nand3_1
XFILLER_80_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09263_ _12070_/A _12338_/C _09026_/A _09024_/Y vssd1 vssd1 vccd1 vccd1 _09269_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_166_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09194_ _09196_/B _09194_/B _09639_/C _12338_/D vssd1 vssd1 vccd1 vccd1 _09202_/A
+ sky130_fd_sc_hd__and4b_1
XFILLER_147_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_796 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08978_ _17421_/A _11920_/D _08978_/C vssd1 vssd1 vccd1 vccd1 _09238_/B sky130_fd_sc_hd__and3_1
XFILLER_57_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10940_ _10940_/A _10940_/B vssd1 vssd1 vccd1 vccd1 _10943_/C sky130_fd_sc_hd__xnor2_1
XFILLER_28_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10871_ _14801_/A _11100_/B _10870_/A vssd1 vssd1 vccd1 vccd1 _10879_/A sky130_fd_sc_hd__a21oi_1
XPHY_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12610_ _12610_/A _12610_/B vssd1 vssd1 vccd1 vccd1 _12612_/C sky130_fd_sc_hd__xnor2_2
XPHY_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13590_ _13590_/A _13590_/B vssd1 vssd1 vccd1 vccd1 _13592_/B sky130_fd_sc_hd__nor2_1
XFILLER_43_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_382 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12541_ _12372_/X _12380_/B _12696_/B vssd1 vssd1 vccd1 vccd1 _12541_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_101_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15260_ _14906_/B _16494_/B1 _15259_/Y vssd1 vssd1 vccd1 vccd1 _17548_/D sky130_fd_sc_hd__a21oi_1
X_12472_ _12473_/A _12473_/B vssd1 vssd1 vccd1 vccd1 _12472_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_61_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_98 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14211_ _14734_/A _14209_/X _14210_/X _14758_/A vssd1 vssd1 vccd1 vccd1 _14211_/X
+ sky130_fd_sc_hd__a22o_1
X_11423_ _17517_/Q _11423_/B _17467_/D _17466_/D vssd1 vssd1 vccd1 vccd1 _11426_/B
+ sky130_fd_sc_hd__and4_1
X_15191_ _14916_/X _14959_/X _16011_/B vssd1 vssd1 vccd1 vccd1 _15805_/B sky130_fd_sc_hd__mux2_1
XFILLER_126_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_9 _15206_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11354_ _11354_/A _11354_/B _11354_/C vssd1 vssd1 vccd1 vccd1 _11361_/A sky130_fd_sc_hd__or3_1
XFILLER_125_424 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14142_ _14142_/A _14229_/A vssd1 vssd1 vccd1 vccd1 _14145_/A sky130_fd_sc_hd__or2_1
XFILLER_4_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10305_ _10305_/A _10305_/B _10305_/C vssd1 vssd1 vccd1 vccd1 _10315_/B sky130_fd_sc_hd__nand3_1
XFILLER_4_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11285_ _11285_/A _11285_/B _11285_/C vssd1 vssd1 vccd1 vccd1 _11311_/A sky130_fd_sc_hd__and3_1
X_14073_ _14074_/A _14074_/B vssd1 vssd1 vccd1 vccd1 _14165_/A sky130_fd_sc_hd__or2_1
XFILLER_152_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13024_ _13024_/A _13024_/B vssd1 vssd1 vccd1 vccd1 _13031_/A sky130_fd_sc_hd__xor2_1
X_10236_ _10236_/A _10236_/B _11006_/C _11027_/D vssd1 vssd1 vccd1 vccd1 _10236_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_117_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10167_ _10167_/A _10278_/A vssd1 vssd1 vccd1 vccd1 _10174_/A sky130_fd_sc_hd__nor2_1
XFILLER_94_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10098_ _10098_/A _10098_/B vssd1 vssd1 vccd1 vccd1 _17138_/A sky130_fd_sc_hd__and2_1
X_14975_ _15081_/A _15820_/A _16025_/A _15415_/A vssd1 vssd1 vccd1 vccd1 _15028_/A
+ sky130_fd_sc_hd__or4_1
X_16714_ _16714_/A _16714_/B vssd1 vssd1 vccd1 vccd1 _16853_/B sky130_fd_sc_hd__or2_1
XFILLER_75_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13926_ _14030_/A _13926_/B vssd1 vssd1 vccd1 vccd1 _13929_/A sky130_fd_sc_hd__nand2_1
XFILLER_47_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_90 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16645_ _16643_/A _16644_/X _16572_/A _16574_/B vssd1 vssd1 vccd1 vccd1 _16648_/B
+ sky130_fd_sc_hd__o211a_1
X_13857_ _13858_/A _13858_/B vssd1 vssd1 vccd1 vccd1 _13961_/B sky130_fd_sc_hd__and2_1
XFILLER_90_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12808_ _12809_/A _12809_/B vssd1 vssd1 vccd1 vccd1 _12972_/A sky130_fd_sc_hd__and2b_1
XFILLER_62_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16576_ _12869_/C _16576_/B vssd1 vssd1 vccd1 vccd1 _16577_/B sky130_fd_sc_hd__nand2b_1
X_13788_ _13893_/A _14360_/D _16722_/A _14318_/A vssd1 vssd1 vccd1 vccd1 _13790_/A
+ sky130_fd_sc_hd__a22oi_1
X_15527_ _15525_/X _15526_/X _16207_/B vssd1 vssd1 vccd1 vccd1 _15527_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_15_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12739_ _12739_/A _12739_/B vssd1 vssd1 vccd1 vccd1 _12741_/B sky130_fd_sc_hd__xnor2_1
XFILLER_31_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15458_ _15901_/S _15458_/B vssd1 vssd1 vccd1 vccd1 _15458_/Y sky130_fd_sc_hd__nor2_1
XFILLER_129_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14409_ _14409_/A _14473_/A _14409_/C vssd1 vssd1 vccd1 vccd1 _14473_/B sky130_fd_sc_hd__nand3_1
XFILLER_117_914 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15389_ _14889_/C _16219_/A1 _12852_/X _15377_/Y _15388_/X vssd1 vssd1 vccd1 vccd1
+ _15390_/B sky130_fd_sc_hd__o311a_1
XFILLER_144_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17128_ _17128_/A _17128_/B vssd1 vssd1 vccd1 vccd1 _17130_/B sky130_fd_sc_hd__and2_1
XFILLER_7_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_906 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17059_ _17037_/B _17009_/B _17014_/B _17014_/C vssd1 vssd1 vccd1 vccd1 _17060_/B
+ sky130_fd_sc_hd__o22ai_1
XFILLER_131_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xmax_cap267 _15147_/Y vssd1 vssd1 vccd1 vccd1 fanout266/A sky130_fd_sc_hd__clkbuf_1
X_09950_ _09951_/B _09951_/C _09951_/A vssd1 vssd1 vccd1 vccd1 _09952_/A sky130_fd_sc_hd__o21a_1
XFILLER_89_319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08901_ _09037_/A _08900_/B _08900_/A vssd1 vssd1 vccd1 vccd1 _08903_/B sky130_fd_sc_hd__o21ba_1
XFILLER_131_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09881_ _10007_/A _10007_/B vssd1 vssd1 vccd1 vccd1 _09881_/X sky130_fd_sc_hd__and2_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08832_ _08832_/A _08832_/B _08832_/C vssd1 vssd1 vccd1 vccd1 _08832_/Y sky130_fd_sc_hd__nor3_4
XFILLER_44_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1029 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08763_ _17393_/A _13208_/C vssd1 vssd1 vccd1 vccd1 _08764_/B sky130_fd_sc_hd__nand2_2
XFILLER_39_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_831 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09315_ _09316_/A _09316_/B _09316_/C vssd1 vssd1 vccd1 vccd1 _09344_/A sky130_fd_sc_hd__a21oi_2
XFILLER_139_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09246_ _09152_/Y _09155_/A _11990_/B _09245_/Y vssd1 vssd1 vccd1 vccd1 _09248_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_166_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09177_ _09357_/A _09364_/A _09357_/C vssd1 vssd1 vccd1 vccd1 _09358_/A sky130_fd_sc_hd__o21a_1
XFILLER_31_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11070_ _11069_/B _11069_/C _11069_/A vssd1 vssd1 vccd1 vccd1 _11070_/Y sky130_fd_sc_hd__o21ai_1
Xoutput79 _17472_/Q vssd1 vssd1 vccd1 vccd1 leds[6] sky130_fd_sc_hd__clkbuf_1
XFILLER_150_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10021_ _10021_/A _10021_/B vssd1 vssd1 vccd1 vccd1 _10136_/B sky130_fd_sc_hd__nor2_1
XFILLER_89_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14760_ _14745_/A _14745_/B _14743_/A vssd1 vssd1 vccd1 vccd1 _14760_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_91_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11972_ _09240_/A _09240_/B _09239_/A vssd1 vssd1 vccd1 vccd1 _11988_/A sky130_fd_sc_hd__a21o_1
XFILLER_16_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13711_ _13814_/A _13710_/B _13817_/A _13710_/D vssd1 vssd1 vccd1 vccd1 _13713_/B
+ sky130_fd_sc_hd__o22a_1
X_10923_ _10799_/Y _14805_/A _10922_/X vssd1 vssd1 vccd1 vccd1 _10924_/B sky130_fd_sc_hd__o21a_1
X_14691_ _14691_/A _14691_/B vssd1 vssd1 vccd1 vccd1 _14692_/B sky130_fd_sc_hd__and2_1
X_16430_ _16604_/B _16589_/B _16758_/B _16814_/B vssd1 vssd1 vccd1 vccd1 _16511_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_44_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13642_ _13642_/A _13642_/B vssd1 vssd1 vccd1 vccd1 _13644_/A sky130_fd_sc_hd__nor2_1
XFILLER_60_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10854_ _10854_/A _10874_/A vssd1 vssd1 vccd1 vccd1 _10865_/A sky130_fd_sc_hd__or2_1
XFILLER_44_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16361_ _16361_/A _16361_/B vssd1 vssd1 vccd1 vccd1 _16362_/B sky130_fd_sc_hd__xnor2_1
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13573_ _14176_/A _13464_/B _13572_/C vssd1 vssd1 vccd1 vccd1 _13574_/B sky130_fd_sc_hd__a21o_1
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10785_ _11132_/B _10899_/D vssd1 vssd1 vccd1 vccd1 _10991_/C sky130_fd_sc_hd__and2_2
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15312_ _15034_/Y _15037_/X _15312_/S vssd1 vssd1 vccd1 vccd1 _15312_/X sky130_fd_sc_hd__mux2_1
XFILLER_169_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12524_ _12524_/A _12524_/B vssd1 vssd1 vccd1 vccd1 _12526_/C sky130_fd_sc_hd__nand2_1
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16292_ _16382_/A _16292_/B vssd1 vssd1 vccd1 vccd1 _16293_/B sky130_fd_sc_hd__nor2_2
XFILLER_13_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15243_ _15244_/A _15244_/B _15244_/C vssd1 vssd1 vccd1 vccd1 _15243_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_9_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12455_ _12280_/X _12284_/A _12626_/A _12454_/Y vssd1 vssd1 vccd1 vccd1 _12626_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_173_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_571 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11406_ _11406_/A _11406_/B vssd1 vssd1 vccd1 vccd1 _11408_/B sky130_fd_sc_hd__xnor2_1
XFILLER_67_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15174_ _15175_/A _15450_/B _15175_/B vssd1 vssd1 vccd1 vccd1 _15174_/Y sky130_fd_sc_hd__o21ai_1
X_12386_ _12020_/Y _12055_/Y _15095_/B vssd1 vssd1 vccd1 vccd1 _12386_/X sky130_fd_sc_hd__mux2_1
X_14125_ _14278_/A _14125_/B vssd1 vssd1 vccd1 vccd1 _14205_/B sky130_fd_sc_hd__or2_1
XFILLER_99_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11337_ _11337_/A _11337_/B vssd1 vssd1 vccd1 vccd1 _11386_/B sky130_fd_sc_hd__nor2_1
XFILLER_141_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14056_ _14057_/A _14057_/B vssd1 vssd1 vccd1 vccd1 _14150_/B sky130_fd_sc_hd__and2b_1
XFILLER_113_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11268_ _11553_/B _11387_/B _11268_/C _11268_/D vssd1 vssd1 vccd1 vccd1 _11320_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_106_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13007_ _12695_/X _13004_/B _13006_/Y vssd1 vssd1 vccd1 vccd1 _13007_/Y sky130_fd_sc_hd__o21bai_1
X_10219_ _10219_/A _10219_/B _10219_/C vssd1 vssd1 vccd1 vccd1 _10342_/A sky130_fd_sc_hd__or3_1
X_11199_ _11201_/A _11201_/B vssd1 vssd1 vccd1 vccd1 _11199_/X sky130_fd_sc_hd__and2b_1
XFILLER_121_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14958_ _14958_/A _15056_/B vssd1 vssd1 vccd1 vccd1 _14958_/Y sky130_fd_sc_hd__nor2_1
XFILLER_47_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13909_ _13908_/A _13908_/B _13908_/C vssd1 vssd1 vccd1 vccd1 _13910_/B sky130_fd_sc_hd__a21oi_1
XFILLER_35_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14889_ _15305_/C _14924_/A _14889_/C _15025_/B vssd1 vssd1 vccd1 vccd1 _14889_/X
+ sky130_fd_sc_hd__or4_2
XFILLER_36_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16628_ _16628_/A _16628_/B vssd1 vssd1 vccd1 vccd1 _16630_/C sky130_fd_sc_hd__xnor2_1
XFILLER_23_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16559_ _16558_/B _16558_/C _16558_/A vssd1 vssd1 vccd1 vccd1 _16560_/B sky130_fd_sc_hd__a21o_1
XFILLER_22_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09100_ _09101_/A _09099_/Y _09654_/C _11815_/B vssd1 vssd1 vccd1 vccd1 _09165_/A
+ sky130_fd_sc_hd__and4bb_1
X_09031_ _09031_/A _09031_/B vssd1 vssd1 vccd1 vccd1 _09032_/B sky130_fd_sc_hd__nor2_1
XFILLER_50_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_880 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1025 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_563 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09933_ _09933_/A _09933_/B vssd1 vssd1 vccd1 vccd1 _09935_/B sky130_fd_sc_hd__nand2_1
Xfanout803 _10525_/D vssd1 vssd1 vccd1 vccd1 _10142_/B sky130_fd_sc_hd__clkbuf_4
Xfanout814 _11281_/B vssd1 vssd1 vccd1 vccd1 _10508_/D sky130_fd_sc_hd__buf_4
XFILLER_113_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout825 _09267_/D vssd1 vssd1 vccd1 vccd1 _12338_/D sky130_fd_sc_hd__buf_2
Xfanout836 _12618_/D vssd1 vssd1 vccd1 vccd1 _09409_/D sky130_fd_sc_hd__buf_2
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09864_ _09865_/A _09864_/B _09864_/C vssd1 vssd1 vccd1 vccd1 _09865_/B sky130_fd_sc_hd__nand3_1
XFILLER_98_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout847 _14849_/A vssd1 vssd1 vccd1 vccd1 _15314_/A sky130_fd_sc_hd__buf_4
Xfanout858 _15238_/A vssd1 vssd1 vccd1 vccd1 _11561_/C sky130_fd_sc_hd__clkbuf_4
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout869 fanout874/X vssd1 vssd1 vccd1 vccd1 _15151_/B sky130_fd_sc_hd__buf_2
X_08815_ _08815_/A _08815_/B vssd1 vssd1 vccd1 vccd1 _08876_/B sky130_fd_sc_hd__xnor2_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09795_ _09795_/A _09795_/B vssd1 vssd1 vccd1 vccd1 _09801_/A sky130_fd_sc_hd__nor2_1
XTAP_3207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08746_ _12068_/A _12068_/B _11861_/B _09030_/C vssd1 vssd1 vccd1 vccd1 _08747_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_45_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_45 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10570_ _10572_/A _10572_/B vssd1 vssd1 vccd1 vccd1 _10586_/A sky130_fd_sc_hd__nor2_1
XFILLER_22_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09229_ _12171_/A _09229_/B vssd1 vssd1 vccd1 vccd1 _09230_/B sky130_fd_sc_hd__nand2_1
XFILLER_154_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12240_ _12241_/B _12241_/A vssd1 vssd1 vccd1 vccd1 _12421_/A sky130_fd_sc_hd__nand2b_1
XFILLER_5_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_777 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12171_ _12171_/A _12328_/B vssd1 vssd1 vccd1 vccd1 _12172_/B sky130_fd_sc_hd__nand2_1
X_11122_ _11122_/A _11122_/B _14850_/A _11518_/C vssd1 vssd1 vccd1 vccd1 _11125_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_150_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_555 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11053_ _11055_/C vssd1 vssd1 vccd1 vccd1 _11053_/Y sky130_fd_sc_hd__inv_2
X_15930_ _15397_/A _16604_/B _16758_/B _16136_/B vssd1 vssd1 vccd1 vccd1 _15933_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_67_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10004_ _10004_/A _10004_/B _10004_/C vssd1 vssd1 vccd1 vccd1 _10005_/C sky130_fd_sc_hd__nand3_1
XFILLER_114_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15861_ _15861_/A _15861_/B vssd1 vssd1 vccd1 vccd1 _15863_/B sky130_fd_sc_hd__xnor2_1
XFILLER_77_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17600_ fanout935/X _17600_/D vssd1 vssd1 vccd1 vccd1 _17600_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14812_ _16005_/B _16005_/C _17119_/B vssd1 vssd1 vccd1 vccd1 _16112_/C sky130_fd_sc_hd__a21bo_1
X_15792_ _15788_/Y _15790_/X _15791_/Y vssd1 vssd1 vccd1 vccd1 _15792_/X sky130_fd_sc_hd__a21o_1
XFILLER_29_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17531_ fanout945/X _17531_/D vssd1 vssd1 vccd1 vccd1 _17531_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_45_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14743_ _14743_/A _14743_/B vssd1 vssd1 vccd1 vccd1 _14745_/A sky130_fd_sc_hd__nand2_1
XFILLER_17_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11955_ _11956_/A _12163_/A _11956_/C vssd1 vssd1 vccd1 vccd1 _11957_/A sky130_fd_sc_hd__o21a_1
XFILLER_18_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10906_ _11006_/B _10954_/D _10905_/D _10954_/A vssd1 vssd1 vccd1 vccd1 _10907_/B
+ sky130_fd_sc_hd__a22oi_1
X_17462_ fanout934/X _17462_/D vssd1 vssd1 vccd1 vccd1 _17462_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_32_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14674_ _14675_/A _17167_/A vssd1 vssd1 vccd1 vccd1 _14674_/X sky130_fd_sc_hd__or2_1
X_11886_ _11886_/A _11886_/B vssd1 vssd1 vccd1 vccd1 _11888_/B sky130_fd_sc_hd__xor2_1
XFILLER_33_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16413_ _16414_/A _16414_/B vssd1 vssd1 vccd1 vccd1 _16509_/A sky130_fd_sc_hd__nand2_1
X_13625_ _13625_/A _13625_/B vssd1 vssd1 vccd1 vccd1 _13625_/Y sky130_fd_sc_hd__nor2_1
X_10837_ _10803_/A _10802_/B _10802_/A vssd1 vssd1 vccd1 vccd1 _10844_/A sky130_fd_sc_hd__o21ba_1
X_17393_ _17393_/A _17425_/B vssd1 vssd1 vccd1 vccd1 _17393_/X sky130_fd_sc_hd__or2_1
XFILLER_41_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16344_ _16344_/A _16344_/B vssd1 vssd1 vccd1 vccd1 _16345_/B sky130_fd_sc_hd__nor2_1
X_13556_ _13680_/B _13556_/B vssd1 vssd1 vccd1 vccd1 _13558_/C sky130_fd_sc_hd__nor2_1
XFILLER_158_655 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10768_ _10655_/A _10655_/B _10669_/B _10669_/A vssd1 vssd1 vccd1 vccd1 _10769_/B
+ sky130_fd_sc_hd__o31ai_1
XFILLER_12_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12507_ _12508_/A _12508_/B _12508_/C vssd1 vssd1 vccd1 vccd1 _12509_/A sky130_fd_sc_hd__o21a_1
XFILLER_173_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16275_ _16276_/A _16276_/B vssd1 vssd1 vccd1 vccd1 _16277_/A sky130_fd_sc_hd__or2_1
XFILLER_121_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13487_ _13603_/B _13486_/C _13486_/A vssd1 vssd1 vccd1 vccd1 _13487_/Y sky130_fd_sc_hd__a21oi_1
X_10699_ _10699_/A _10699_/B vssd1 vssd1 vccd1 vccd1 _10701_/B sky130_fd_sc_hd__xnor2_2
X_15226_ _15226_/A _15226_/B vssd1 vssd1 vccd1 vccd1 _15228_/A sky130_fd_sc_hd__xnor2_1
X_12438_ _12592_/B _12592_/D _12439_/D _12592_/A vssd1 vssd1 vccd1 vccd1 _12440_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_8_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_563 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15157_ _15157_/A _15157_/B vssd1 vssd1 vccd1 vccd1 _15159_/B sky130_fd_sc_hd__xnor2_1
X_12369_ _12170_/B _12172_/B _12170_/A vssd1 vssd1 vccd1 vccd1 _12370_/B sky130_fd_sc_hd__o21ba_1
XFILLER_153_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14108_ _14108_/A _14108_/B vssd1 vssd1 vccd1 vccd1 _14110_/B sky130_fd_sc_hd__xor2_1
X_15088_ _16127_/A _15088_/B vssd1 vssd1 vccd1 vccd1 _15088_/Y sky130_fd_sc_hd__nand2_1
XFILLER_114_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14039_ _13950_/A _14181_/B _13951_/A _13949_/B vssd1 vssd1 vccd1 vccd1 _14043_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_67_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09580_ _09581_/A _09581_/B _09581_/C vssd1 vssd1 vccd1 vccd1 _09580_/X sky130_fd_sc_hd__a21o_1
XFILLER_63_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_817 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09014_ _09014_/A _09014_/B vssd1 vssd1 vccd1 vccd1 _09016_/C sky130_fd_sc_hd__xnor2_1
XFILLER_163_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout600 _11630_/A vssd1 vssd1 vccd1 vccd1 _11520_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_137_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout611 _17510_/Q vssd1 vssd1 vccd1 vccd1 _11651_/A sky130_fd_sc_hd__clkbuf_4
Xfanout622 _08967_/B vssd1 vssd1 vccd1 vccd1 _11932_/B sky130_fd_sc_hd__buf_4
X_09916_ _09973_/A _09973_/B vssd1 vssd1 vccd1 vccd1 _10059_/A sky130_fd_sc_hd__nor2_2
Xfanout633 _13037_/B vssd1 vssd1 vccd1 vccd1 _14094_/B sky130_fd_sc_hd__clkbuf_4
Xfanout644 _17065_/A vssd1 vssd1 vccd1 vccd1 _14433_/B sky130_fd_sc_hd__buf_4
Xfanout655 _12445_/C vssd1 vssd1 vccd1 vccd1 _11895_/C sky130_fd_sc_hd__clkbuf_4
Xfanout666 _17503_/Q vssd1 vssd1 vccd1 vccd1 _13522_/D sky130_fd_sc_hd__clkbuf_4
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout677 _17502_/Q vssd1 vssd1 vccd1 vccd1 _16859_/A sky130_fd_sc_hd__buf_4
X_09847_ _09847_/A _09847_/B vssd1 vssd1 vccd1 vccd1 _09976_/A sky130_fd_sc_hd__xnor2_1
XFILLER_101_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout688 fanout690/X vssd1 vssd1 vccd1 vccd1 _14863_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_100_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout699 _17500_/Q vssd1 vssd1 vccd1 vccd1 fanout699/X sky130_fd_sc_hd__buf_8
XTAP_3004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09778_ _14954_/A _11808_/B _09655_/A _09653_/Y vssd1 vssd1 vccd1 vccd1 _09784_/B
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_3037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08729_ input28/X vssd1 vssd1 vccd1 vccd1 _17362_/A sky130_fd_sc_hd__inv_2
XTAP_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11740_ _11737_/Y _11753_/A _11732_/Y _11733_/X vssd1 vssd1 vccd1 vccd1 _11758_/A
+ sky130_fd_sc_hd__a211oi_2
XTAP_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11671_ _15524_/C _11671_/B vssd1 vssd1 vccd1 vccd1 _11672_/C sky130_fd_sc_hd__or2_1
XFILLER_30_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13410_ _13411_/A _13411_/B _13411_/C vssd1 vssd1 vccd1 vccd1 _13545_/A sky130_fd_sc_hd__a21o_1
X_10622_ _10716_/A _10621_/B _10621_/A vssd1 vssd1 vccd1 vccd1 _10624_/B sky130_fd_sc_hd__o21ba_1
XFILLER_41_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14390_ _14456_/A _14456_/B vssd1 vssd1 vccd1 vccd1 _14393_/C sky130_fd_sc_hd__xnor2_1
XFILLER_10_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13341_ _13341_/A _13462_/A vssd1 vssd1 vccd1 vccd1 _13342_/C sky130_fd_sc_hd__and2_1
X_10553_ _10566_/B _10553_/B vssd1 vssd1 vccd1 vccd1 _10555_/B sky130_fd_sc_hd__nand2_1
XFILLER_6_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_647 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16060_ _16060_/A _16060_/B vssd1 vssd1 vccd1 vccd1 _16070_/A sky130_fd_sc_hd__xor2_1
XFILLER_155_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13272_ _14756_/A1 _13270_/Y _13386_/B _13143_/Y _13146_/X vssd1 vssd1 vccd1 vccd1
+ _17585_/D sky130_fd_sc_hd__a32o_1
XFILLER_108_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10484_ _10484_/A _10484_/B vssd1 vssd1 vccd1 vccd1 _10497_/B sky130_fd_sc_hd__xor2_1
XFILLER_6_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_134 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15011_ _15011_/A _16389_/A _15011_/C vssd1 vssd1 vccd1 vccd1 _15011_/X sky130_fd_sc_hd__and3_1
X_12223_ _11837_/Y _11840_/Y _17365_/A vssd1 vssd1 vccd1 vccd1 _12223_/X sky130_fd_sc_hd__mux2_1
XFILLER_135_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12154_ _12316_/B _12152_/X _11917_/X _11947_/X vssd1 vssd1 vccd1 vccd1 _12193_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_78_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11105_ _11112_/B _11105_/B vssd1 vssd1 vccd1 vccd1 _11252_/A sky130_fd_sc_hd__nand2_1
XFILLER_150_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16962_ _17131_/A _17014_/A vssd1 vssd1 vccd1 vccd1 _16962_/Y sky130_fd_sc_hd__nand2_1
X_12085_ _12085_/A _12085_/B _12085_/C vssd1 vssd1 vccd1 vccd1 _12098_/B sky130_fd_sc_hd__nand3_1
XFILLER_110_216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11036_ _11036_/A _11036_/B vssd1 vssd1 vccd1 vccd1 _11038_/B sky130_fd_sc_hd__xnor2_1
X_15913_ _15913_/A _16939_/B vssd1 vssd1 vccd1 vccd1 _16028_/A sky130_fd_sc_hd__nor2_1
XFILLER_110_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16893_ _16893_/A _16893_/B vssd1 vssd1 vccd1 vccd1 _16895_/B sky130_fd_sc_hd__xnor2_1
XFILLER_49_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15844_ _16807_/A _16054_/B vssd1 vssd1 vccd1 vccd1 _16681_/D sky130_fd_sc_hd__nand2_2
XFILLER_77_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15775_ _15775_/A _15775_/B vssd1 vssd1 vccd1 vccd1 _15776_/C sky130_fd_sc_hd__xor2_1
XTAP_3560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12987_ _12825_/A _12826_/Y _13125_/B _12986_/Y vssd1 vssd1 vccd1 vccd1 _12987_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17514_ fanout950/X _17514_/D vssd1 vssd1 vccd1 vccd1 _17514_/Q sky130_fd_sc_hd__dfxtp_2
X_14726_ _14727_/A _14750_/A _14726_/C vssd1 vssd1 vccd1 vccd1 _14726_/X sky130_fd_sc_hd__and3_1
X_11938_ _09004_/A _09004_/B _09002_/X vssd1 vssd1 vccd1 vccd1 _11939_/B sky130_fd_sc_hd__a21oi_1
XTAP_2870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17445_ fanout940/X _17445_/D vssd1 vssd1 vccd1 vccd1 _17445_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14657_ _14658_/A _14658_/B _14658_/C vssd1 vssd1 vccd1 vccd1 _14698_/A sky130_fd_sc_hd__o21ai_1
X_11869_ _17393_/A _12077_/C vssd1 vssd1 vccd1 vccd1 _11871_/B sky130_fd_sc_hd__nand2_1
XFILLER_33_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13608_ _13486_/X _13490_/C _13718_/A _13607_/X vssd1 vssd1 vccd1 vccd1 _13718_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_159_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17376_ input64/X _17424_/A2 _17375_/X _17388_/C1 vssd1 vssd1 vccd1 vccd1 _17516_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_158_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14588_ _14763_/S _14586_/X _14587_/Y _14541_/X _14543_/Y vssd1 vssd1 vccd1 vccd1
+ _17600_/D sky130_fd_sc_hd__a32o_1
XFILLER_158_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16327_ _16328_/A _16328_/B vssd1 vssd1 vccd1 vccd1 _16329_/A sky130_fd_sc_hd__and2_1
XFILLER_158_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13539_ _13643_/A _13846_/B _13408_/A _13406_/B vssd1 vssd1 vccd1 vccd1 _13541_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_158_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16258_ _16174_/A _16174_/B _16175_/B _16175_/A vssd1 vssd1 vccd1 vccd1 _16272_/A
+ sky130_fd_sc_hd__a22oi_2
XFILLER_145_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15209_ _15203_/X _15208_/X _14906_/B vssd1 vssd1 vccd1 vccd1 _15397_/A sky130_fd_sc_hd__a21boi_4
XFILLER_173_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16189_ _16189_/A _16189_/B vssd1 vssd1 vccd1 vccd1 _16191_/A sky130_fd_sc_hd__nor2_1
XFILLER_114_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09701_ _10244_/A _10508_/D _09701_/C vssd1 vssd1 vccd1 vccd1 _09706_/B sky130_fd_sc_hd__and3_1
XFILLER_83_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09632_ _09632_/A _09632_/B vssd1 vssd1 vccd1 vccd1 _09665_/A sky130_fd_sc_hd__xnor2_1
XFILLER_28_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09563_ _16990_/B _09563_/B vssd1 vssd1 vccd1 vccd1 _09565_/B sky130_fd_sc_hd__xnor2_4
XFILLER_71_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09494_ _09493_/A _11808_/B _14948_/B vssd1 vssd1 vccd1 vccd1 _09494_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_130_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1042 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout430 _13641_/A vssd1 vssd1 vccd1 vccd1 _13852_/A sky130_fd_sc_hd__buf_2
Xfanout441 _16209_/C vssd1 vssd1 vccd1 vccd1 _12722_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_87_940 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout452 _10244_/A vssd1 vssd1 vccd1 vccd1 _11027_/B sky130_fd_sc_hd__buf_4
Xfanout463 _14873_/B vssd1 vssd1 vccd1 vccd1 _11006_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_58_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout474 _17522_/Q vssd1 vssd1 vccd1 vccd1 _17387_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_47_815 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_761 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout485 _11095_/A vssd1 vssd1 vccd1 vccd1 _10963_/A sky130_fd_sc_hd__buf_2
XFILLER_86_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12910_ _12910_/A _12910_/B _12910_/C vssd1 vssd1 vccd1 vccd1 _12911_/B sky130_fd_sc_hd__or3_1
Xfanout496 _09299_/B vssd1 vssd1 vccd1 vccd1 _15262_/B sky130_fd_sc_hd__buf_4
XFILLER_19_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_1016 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13890_ _13891_/A _13891_/B vssd1 vssd1 vccd1 vccd1 _14013_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12841_ _13003_/A _12698_/B _12693_/X vssd1 vssd1 vccd1 vccd1 _12842_/B sky130_fd_sc_hd__o21ai_1
XTAP_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15560_ _15558_/Y _15675_/A vssd1 vssd1 vccd1 vccd1 _15655_/B sky130_fd_sc_hd__and2b_1
XTAP_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12772_ _17421_/A _13067_/D vssd1 vssd1 vccd1 vccd1 _12773_/B sky130_fd_sc_hd__nand2_1
XTAP_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14511_ _14509_/A _14509_/B _14509_/C vssd1 vssd1 vccd1 vccd1 _14512_/B sky130_fd_sc_hd__o21a_1
XTAP_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11723_ _10766_/C _10766_/B _10764_/X vssd1 vssd1 vccd1 vccd1 _11725_/B sky130_fd_sc_hd__a21bo_1
XTAP_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15491_ _16315_/D _15492_/B vssd1 vssd1 vccd1 vccd1 _16061_/B sky130_fd_sc_hd__nor2_2
XTAP_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17230_ _17444_/Q _17275_/A2 _17228_/X _17229_/X _17364_/C1 vssd1 vssd1 vccd1 vccd1
+ _17444_/D sky130_fd_sc_hd__o221a_1
XFILLER_70_1000 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14442_ _14367_/A _17023_/A _14370_/A vssd1 vssd1 vccd1 vccd1 _14443_/B sky130_fd_sc_hd__o21ba_1
X_11654_ _14796_/A _11675_/C _11650_/X vssd1 vssd1 vccd1 vccd1 _11676_/A sky130_fd_sc_hd__o21a_1
X_10605_ _15393_/A _10963_/C vssd1 vssd1 vccd1 vccd1 _10699_/A sky130_fd_sc_hd__nand2_1
X_17161_ _11932_/B _17140_/B _17160_/Y vssd1 vssd1 vccd1 vccd1 _17166_/B sky130_fd_sc_hd__o21ai_1
X_14373_ _14445_/A _14373_/B vssd1 vssd1 vccd1 vccd1 _14376_/A sky130_fd_sc_hd__and2_1
X_11585_ _11543_/A _11543_/B _11542_/X vssd1 vssd1 vccd1 vccd1 _11586_/C sky130_fd_sc_hd__o21bai_1
XFILLER_127_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16112_ _16315_/A _16112_/B _16112_/C vssd1 vssd1 vccd1 vccd1 _16112_/X sky130_fd_sc_hd__and3_1
XFILLER_167_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13324_ _13324_/A _13324_/B vssd1 vssd1 vccd1 vccd1 _13326_/C sky130_fd_sc_hd__xnor2_1
XFILLER_6_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10536_ _10536_/A _10536_/B vssd1 vssd1 vccd1 vccd1 _10637_/B sky130_fd_sc_hd__xnor2_1
XFILLER_128_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17092_ _17118_/A _17092_/B vssd1 vssd1 vccd1 vccd1 _17093_/C sky130_fd_sc_hd__xnor2_1
XFILLER_127_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_466 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16043_ _16043_/A _16043_/B vssd1 vssd1 vccd1 vccd1 _16044_/B sky130_fd_sc_hd__and2_1
XFILLER_115_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13255_ _13252_/A _13253_/Y _13118_/A _13119_/Y vssd1 vssd1 vccd1 vccd1 _13256_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_108_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10467_ _10467_/A _10470_/A vssd1 vssd1 vccd1 vccd1 _10581_/C sky130_fd_sc_hd__nor2_1
XFILLER_109_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_842 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12206_ _12371_/B _12206_/B _12206_/C vssd1 vssd1 vccd1 vccd1 _12375_/B sky130_fd_sc_hd__nor3_1
XFILLER_142_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13186_ _13186_/A _13186_/B vssd1 vssd1 vccd1 vccd1 _13187_/B sky130_fd_sc_hd__and2_1
X_10398_ _14788_/A _10647_/D _10293_/A _10291_/Y vssd1 vssd1 vccd1 vccd1 _10399_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_69_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12137_ _12138_/A _12138_/B _12138_/C vssd1 vssd1 vccd1 vccd1 _12305_/A sky130_fd_sc_hd__o21ai_1
XFILLER_111_514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16945_ _16065_/B _15658_/Y _17119_/C _16883_/C _16887_/A vssd1 vssd1 vccd1 vccd1
+ _16947_/B sky130_fd_sc_hd__a41o_1
X_12068_ _12068_/A _12068_/B _13208_/D _12942_/D vssd1 vssd1 vccd1 vccd1 _12239_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_96_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11019_ _11020_/A _11020_/B vssd1 vssd1 vccd1 vccd1 _11019_/X sky130_fd_sc_hd__and2_1
XFILLER_64_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16876_ _16859_/A _17170_/B1 _16857_/Y _16875_/X vssd1 vssd1 vccd1 vccd1 _17567_/D
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_37_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15827_ _15827_/A _15827_/B vssd1 vssd1 vccd1 vccd1 _15837_/A sky130_fd_sc_hd__xor2_2
XFILLER_53_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15758_ _15759_/A _15759_/B vssd1 vssd1 vccd1 vccd1 _15758_/X sky130_fd_sc_hd__or2_1
XFILLER_92_497 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_339 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14709_ _14677_/A _14677_/B _14674_/X vssd1 vssd1 vccd1 vccd1 _14744_/A sky130_fd_sc_hd__o21ai_1
XFILLER_61_873 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15689_ _15782_/B _15689_/B vssd1 vssd1 vccd1 vccd1 _15690_/C sky130_fd_sc_hd__nand2_1
XFILLER_166_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17428_ input68/X _17428_/B _17428_/C _17428_/D vssd1 vssd1 vccd1 vccd1 _17542_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_159_761 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17359_ input60/X _17359_/B _17359_/C vssd1 vssd1 vccd1 vccd1 _17359_/X sky130_fd_sc_hd__or3_1
XFILLER_147_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08994_ _08994_/A _08994_/B vssd1 vssd1 vccd1 vccd1 _09009_/A sky130_fd_sc_hd__xnor2_1
XFILLER_87_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09615_ _09746_/A _09754_/A _09746_/C vssd1 vssd1 vccd1 vccd1 _09747_/A sky130_fd_sc_hd__o21ai_2
XFILLER_141_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_987 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09546_ _09546_/A _09546_/B vssd1 vssd1 vccd1 vccd1 _09574_/A sky130_fd_sc_hd__xor2_1
XFILLER_52_840 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09477_ _09478_/B _09603_/A _09478_/A vssd1 vssd1 vccd1 vccd1 _09480_/A sky130_fd_sc_hd__a21o_1
XFILLER_51_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xwire116 wire116/A vssd1 vssd1 vccd1 vccd1 wire116/X sky130_fd_sc_hd__clkbuf_2
XFILLER_165_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11370_ _11370_/A _15373_/C _17467_/D _17466_/D vssd1 vssd1 vccd1 vccd1 _11370_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_153_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10321_ _10321_/A _10321_/B _15003_/B _17478_/Q vssd1 vssd1 vccd1 vccd1 _10445_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_4_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13040_ _13040_/A _13040_/B _13040_/C vssd1 vssd1 vccd1 vccd1 _13041_/B sky130_fd_sc_hd__or3_1
XFILLER_3_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10252_ _10253_/A _10253_/B vssd1 vssd1 vccd1 vccd1 _10267_/A sky130_fd_sc_hd__nand2b_1
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10183_ _10183_/A _10307_/A vssd1 vssd1 vccd1 vccd1 _10184_/C sky130_fd_sc_hd__nor2_1
XFILLER_105_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_759 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14991_ _10072_/B _09937_/B _09843_/D _09843_/C _09925_/A _14958_/A vssd1 vssd1 vccd1
+ vccd1 _14992_/B sky130_fd_sc_hd__mux4_1
Xfanout260 _17429_/C vssd1 vssd1 vccd1 vccd1 _17321_/C sky130_fd_sc_hd__buf_2
XFILLER_120_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout271 _17134_/C vssd1 vssd1 vccd1 vccd1 _16965_/B sky130_fd_sc_hd__buf_2
Xfanout282 _17363_/A vssd1 vssd1 vccd1 vccd1 _12025_/A sky130_fd_sc_hd__buf_2
XFILLER_93_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13942_ _17070_/B _13940_/X _14032_/B _13842_/X vssd1 vssd1 vccd1 vccd1 _17591_/D
+ sky130_fd_sc_hd__o31ai_1
X_16730_ _16730_/A _16730_/B vssd1 vssd1 vccd1 vccd1 _16730_/Y sky130_fd_sc_hd__xnor2_1
Xfanout293 fanout299/X vssd1 vssd1 vccd1 vccd1 _12848_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_101_580 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_442 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16661_ _16938_/B _16662_/C _16662_/D _16747_/A vssd1 vssd1 vccd1 vccd1 _16661_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_19_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13873_ _13873_/A _13873_/B vssd1 vssd1 vccd1 vccd1 _13874_/B sky130_fd_sc_hd__or2_1
X_15612_ _15610_/Y _15611_/X _16911_/A vssd1 vssd1 vccd1 vccd1 _15612_/X sky130_fd_sc_hd__o21a_1
X_12824_ _12824_/A _12824_/B vssd1 vssd1 vccd1 vccd1 _12825_/C sky130_fd_sc_hd__nand2_1
XFILLER_62_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16592_ _16814_/B _16935_/B _16591_/C vssd1 vssd1 vccd1 vccd1 _16593_/B sky130_fd_sc_hd__a21oi_1
XFILLER_27_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15543_ _10716_/A _17163_/A2 _15542_/X vssd1 vssd1 vccd1 vccd1 _15543_/X sky130_fd_sc_hd__o21ba_1
X_12755_ _12755_/A _12755_/B _12755_/C vssd1 vssd1 vccd1 vccd1 _12757_/A sky130_fd_sc_hd__or3_1
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11706_ _15793_/A _15793_/B _15889_/A _11705_/Y _11704_/B vssd1 vssd1 vccd1 vccd1
+ _15997_/B sky130_fd_sc_hd__a32o_1
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15474_ _14899_/X _14968_/X _16827_/A _11675_/B vssd1 vssd1 vccd1 vccd1 _15645_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_42_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12686_ _12528_/A _12530_/A _12684_/X _12685_/Y vssd1 vssd1 vccd1 vccd1 _12689_/A
+ sky130_fd_sc_hd__o211a_1
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17213_ _17580_/Q _17225_/A2 _17225_/B1 vssd1 vssd1 vccd1 vccd1 _17213_/X sky130_fd_sc_hd__a21o_1
X_14425_ _14641_/B _14865_/B _14426_/D _14641_/A vssd1 vssd1 vccd1 vccd1 _14427_/A
+ sky130_fd_sc_hd__a22oi_1
X_11637_ _11637_/A _11637_/B vssd1 vssd1 vccd1 vccd1 _11659_/B sky130_fd_sc_hd__nor2_1
XFILLER_30_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17144_ _17164_/C _16011_/X _17140_/X _17143_/X vssd1 vssd1 vccd1 vccd1 _17144_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_128_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14356_ _12706_/X _12710_/B _14356_/S vssd1 vssd1 vccd1 vccd1 _16735_/B sky130_fd_sc_hd__mux2_1
X_11568_ _11568_/A _11568_/B _11568_/C vssd1 vssd1 vccd1 vccd1 _11603_/A sky130_fd_sc_hd__and3_1
XFILLER_129_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13307_ _13308_/A _13308_/B _13308_/C vssd1 vssd1 vccd1 vccd1 _13309_/A sky130_fd_sc_hd__a21o_1
XFILLER_6_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10519_ _10519_/A _10519_/B _10519_/C vssd1 vssd1 vccd1 vccd1 _10519_/Y sky130_fd_sc_hd__nor3_2
XFILLER_7_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17075_ _14434_/Y _17075_/A2 _17074_/X vssd1 vssd1 vccd1 vccd1 _17077_/C sky130_fd_sc_hd__a21o_1
X_14287_ _12549_/X _14210_/B _14482_/B1 vssd1 vssd1 vccd1 vccd1 _14287_/X sky130_fd_sc_hd__o21a_1
XFILLER_170_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11499_ _11499_/A _11499_/B _11499_/C vssd1 vssd1 vccd1 vccd1 _11539_/A sky130_fd_sc_hd__nor3_2
XFILLER_143_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16026_ _16026_/A _16026_/B vssd1 vssd1 vccd1 vccd1 _16028_/B sky130_fd_sc_hd__xnor2_2
X_13238_ _13238_/A _13238_/B vssd1 vssd1 vccd1 vccd1 _13239_/B sky130_fd_sc_hd__nand2_1
XFILLER_152_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13169_ _13658_/A _13414_/B _14094_/B _14008_/B vssd1 vssd1 vccd1 vccd1 _13170_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16928_ _14734_/A _14543_/B _16924_/Y _16927_/X vssd1 vssd1 vccd1 vccd1 _16928_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_37_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16859_ _16859_/A _17153_/B vssd1 vssd1 vccd1 vccd1 _16859_/Y sky130_fd_sc_hd__nor2_1
XFILLER_92_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09400_ _09311_/A _09316_/B _09311_/C vssd1 vssd1 vccd1 vccd1 _09401_/B sky130_fd_sc_hd__a21oi_1
XFILLER_19_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09331_ _09332_/B _09463_/A _09332_/A vssd1 vssd1 vccd1 vccd1 _09334_/A sky130_fd_sc_hd__a21o_1
XFILLER_40_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09262_ _09262_/A _09262_/B vssd1 vssd1 vccd1 vccd1 _09290_/A sky130_fd_sc_hd__xnor2_1
XFILLER_166_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09193_ _09194_/B vssd1 vssd1 vccd1 vccd1 _09193_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_174_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_926 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_970 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08977_ _08977_/A _09238_/A vssd1 vssd1 vccd1 vccd1 _08978_/C sky130_fd_sc_hd__nor2_1
XFILLER_29_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_976 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10870_ _10870_/A _10870_/B vssd1 vssd1 vccd1 vccd1 _11100_/B sky130_fd_sc_hd__nor2_1
XFILLER_71_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_851 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09529_ _09391_/C _09399_/Y _09458_/X _09628_/A vssd1 vssd1 vccd1 vccd1 _09530_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12540_ _12540_/A _12540_/B vssd1 vssd1 vccd1 vccd1 _12696_/B sky130_fd_sc_hd__xnor2_1
XFILLER_169_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12471_ _12471_/A _12592_/C _12471_/C vssd1 vssd1 vccd1 vccd1 _12473_/B sky130_fd_sc_hd__and3_1
XFILLER_12_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_898 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14210_ _14210_/A _14210_/B vssd1 vssd1 vccd1 vccd1 _14210_/X sky130_fd_sc_hd__or2_1
X_11422_ _11395_/B _11383_/C _11383_/B vssd1 vssd1 vccd1 vccd1 _11435_/B sky130_fd_sc_hd__a21o_1
X_15190_ _10180_/A _14918_/Y _15189_/Y _15805_/A vssd1 vssd1 vccd1 vccd1 _15190_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_165_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14141_ _14290_/A _14708_/B _16651_/A _14141_/D vssd1 vssd1 vccd1 vccd1 _14229_/A
+ sky130_fd_sc_hd__and4_1
X_11353_ _11351_/A _11351_/C _11402_/A vssd1 vssd1 vccd1 vccd1 _11354_/C sky130_fd_sc_hd__a21oi_1
XFILLER_4_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10304_ _10305_/B _10305_/C _10305_/A vssd1 vssd1 vccd1 vccd1 _10315_/A sky130_fd_sc_hd__a21o_1
X_14072_ _14072_/A _14072_/B vssd1 vssd1 vccd1 vccd1 _14074_/B sky130_fd_sc_hd__nor2_1
X_11284_ _11352_/A _11284_/B vssd1 vssd1 vccd1 vccd1 _11285_/C sky130_fd_sc_hd__and2_1
XFILLER_98_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13023_ _13024_/A _13024_/B vssd1 vssd1 vccd1 vccd1 _13165_/A sky130_fd_sc_hd__nand2_1
XFILLER_117_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10235_ _10236_/B _11027_/D vssd1 vssd1 vccd1 vccd1 _10709_/A sky130_fd_sc_hd__nand2_2
XFILLER_79_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10166_ _10167_/A _10165_/Y _14788_/A _10993_/D vssd1 vssd1 vccd1 vccd1 _10278_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_67_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_943 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10097_ _10097_/A _10097_/B vssd1 vssd1 vccd1 vccd1 _10098_/B sky130_fd_sc_hd__nand2_1
X_14974_ _15750_/A vssd1 vssd1 vccd1 vccd1 _15415_/A sky130_fd_sc_hd__inv_2
X_16713_ _16714_/A _16714_/B vssd1 vssd1 vccd1 vccd1 _16853_/A sky130_fd_sc_hd__nand2_1
X_13925_ _13925_/A _13925_/B _13925_/C vssd1 vssd1 vccd1 vccd1 _13926_/B sky130_fd_sc_hd__nand3_1
XFILLER_48_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13856_ _13856_/A _13856_/B vssd1 vssd1 vccd1 vccd1 _13858_/B sky130_fd_sc_hd__xnor2_1
X_16644_ _16651_/A _16644_/B _16644_/C vssd1 vssd1 vccd1 vccd1 _16644_/X sky130_fd_sc_hd__and3b_1
XFILLER_74_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12807_ _12807_/A _12807_/B vssd1 vssd1 vccd1 vccd1 _12809_/B sky130_fd_sc_hd__xnor2_1
XFILLER_22_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13787_ _13787_/A _13787_/B vssd1 vssd1 vccd1 vccd1 _13805_/A sky130_fd_sc_hd__xnor2_1
X_16575_ _16481_/A _16482_/Y _16572_/Y _16574_/Y vssd1 vssd1 vccd1 vccd1 _16575_/X
+ sky130_fd_sc_hd__a31o_1
X_10999_ _10999_/A _10999_/B _10999_/C vssd1 vssd1 vccd1 vccd1 _10999_/X sky130_fd_sc_hd__and3_1
XFILLER_62_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15526_ _15524_/B _11671_/B _15447_/A vssd1 vssd1 vccd1 vccd1 _15526_/X sky130_fd_sc_hd__a21o_1
XFILLER_15_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12738_ _12739_/A _12739_/B vssd1 vssd1 vccd1 vccd1 _12903_/A sky130_fd_sc_hd__and2b_1
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15457_ _15457_/A _15457_/B _15457_/C vssd1 vssd1 vccd1 vccd1 _15467_/C sky130_fd_sc_hd__or3_1
X_12669_ _12816_/A _12669_/B vssd1 vssd1 vccd1 vccd1 _12670_/B sky130_fd_sc_hd__and2_1
XFILLER_129_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14408_ _14424_/B _14406_/Y _14340_/B _14342_/A vssd1 vssd1 vccd1 vccd1 _14409_/C
+ sky130_fd_sc_hd__o211ai_1
XFILLER_163_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_550 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15388_ _16582_/A _15380_/X _15387_/X _15379_/X vssd1 vssd1 vccd1 vccd1 _15388_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_144_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17127_ _17127_/A _17127_/B vssd1 vssd1 vccd1 vccd1 _17128_/B sky130_fd_sc_hd__nand2_1
X_14339_ _14336_/X _14337_/Y _14222_/A _14265_/B vssd1 vssd1 vccd1 vccd1 _14340_/C
+ sky130_fd_sc_hd__o211ai_1
XFILLER_143_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17058_ _17096_/A _17058_/B vssd1 vssd1 vccd1 vccd1 _17062_/A sky130_fd_sc_hd__nor2_1
XFILLER_132_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08900_ _08900_/A _08900_/B vssd1 vssd1 vccd1 vccd1 _09037_/B sky130_fd_sc_hd__nor2_1
XFILLER_103_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16009_ _17119_/B _14931_/X _16008_/X vssd1 vssd1 vccd1 vccd1 _16017_/A sky130_fd_sc_hd__o21ba_1
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09880_ _09880_/A _09880_/B vssd1 vssd1 vccd1 vccd1 _10007_/B sky130_fd_sc_hd__nor2_1
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08831_ _08831_/A _08831_/B _08831_/C vssd1 vssd1 vccd1 vccd1 _08832_/C sky130_fd_sc_hd__nor3_2
XFILLER_112_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08762_ _08760_/Y _16302_/A _08758_/X vssd1 vssd1 vccd1 vccd1 _08764_/A sky130_fd_sc_hd__o21ai_4
XFILLER_39_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09314_ _09314_/A _09314_/B vssd1 vssd1 vccd1 vccd1 _09316_/C sky130_fd_sc_hd__xnor2_1
XFILLER_80_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_854 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_528 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_876 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09245_ _09245_/A _09245_/B _09245_/C vssd1 vssd1 vccd1 vccd1 _09245_/Y sky130_fd_sc_hd__nand3_1
X_09176_ _09176_/A _09176_/B vssd1 vssd1 vccd1 vccd1 _09357_/C sky130_fd_sc_hd__xnor2_1
XFILLER_108_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10020_ _09894_/C _10299_/D _09895_/A _09893_/Y vssd1 vssd1 vccd1 vccd1 _10021_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_163_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11971_ _11971_/A _11971_/B vssd1 vssd1 vccd1 vccd1 _11971_/X sky130_fd_sc_hd__and2_1
XFILLER_57_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13710_ _13814_/A _13710_/B _13817_/A _13710_/D vssd1 vssd1 vccd1 vccd1 wire118/A
+ sky130_fd_sc_hd__nor4_1
X_10922_ _14787_/A _10920_/B _10799_/B _14786_/A vssd1 vssd1 vccd1 vccd1 _10922_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_16_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14690_ _14691_/A _14691_/B vssd1 vssd1 vccd1 vccd1 _14723_/A sky130_fd_sc_hd__nor2_1
XFILLER_44_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13641_ _13641_/A _13745_/B _13844_/C _13846_/B vssd1 vssd1 vccd1 vccd1 _13642_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_16_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10853_ _10854_/A _10852_/Y _11124_/C _10970_/B vssd1 vssd1 vccd1 vccd1 _10874_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_32_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16360_ _16361_/A _16361_/B vssd1 vssd1 vccd1 vccd1 _16443_/B sky130_fd_sc_hd__nand2b_1
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13572_ _13903_/A _16789_/A _13572_/C vssd1 vssd1 vccd1 vccd1 _13702_/B sky130_fd_sc_hd__nand3_1
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10784_ _10784_/A _10784_/B vssd1 vssd1 vccd1 vccd1 _16866_/A sky130_fd_sc_hd__xnor2_2
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15311_ _15456_/B _15311_/B _14801_/X vssd1 vssd1 vccd1 vccd1 _15321_/B sky130_fd_sc_hd__or3b_1
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12523_ _12522_/A _12522_/B _12522_/C vssd1 vssd1 vccd1 vccd1 _12524_/B sky130_fd_sc_hd__o21ai_1
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16291_ _16382_/B _16562_/C vssd1 vssd1 vccd1 vccd1 _16293_/A sky130_fd_sc_hd__nand2b_2
XFILLER_13_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15242_ _15454_/A _15242_/B _15242_/C vssd1 vssd1 vccd1 vccd1 _15257_/A sky130_fd_sc_hd__and3_1
X_12454_ _12454_/A _12454_/B _12454_/C vssd1 vssd1 vccd1 vccd1 _12454_/Y sky130_fd_sc_hd__nand3_1
XFILLER_126_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11405_ _11405_/A vssd1 vssd1 vccd1 vccd1 _11419_/A sky130_fd_sc_hd__inv_2
XFILLER_138_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15173_ _15235_/C _15173_/B vssd1 vssd1 vccd1 vccd1 _15173_/Y sky130_fd_sc_hd__nand2_1
XFILLER_153_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12385_ _12051_/Y _12053_/Y _14948_/A vssd1 vssd1 vccd1 vccd1 _12385_/X sky130_fd_sc_hd__mux2_1
XFILLER_165_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14124_ _14278_/A _14125_/B vssd1 vssd1 vccd1 vccd1 _14124_/Y sky130_fd_sc_hd__nand2_1
X_11336_ _11518_/B _15617_/A _14851_/A _11561_/A vssd1 vssd1 vccd1 vccd1 _11337_/B
+ sky130_fd_sc_hd__a22oi_1
XFILLER_140_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14055_ _14158_/B _14055_/B vssd1 vssd1 vccd1 vccd1 _14057_/B sky130_fd_sc_hd__nor2_1
X_11267_ _11553_/A _11437_/D _11561_/C _11427_/A vssd1 vssd1 vccd1 vccd1 _11268_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_97_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13006_ _12693_/X _12840_/B _12838_/Y vssd1 vssd1 vccd1 vccd1 _13006_/Y sky130_fd_sc_hd__a21oi_1
X_10218_ _10216_/A _10216_/B _10216_/C vssd1 vssd1 vccd1 vccd1 _10219_/C sky130_fd_sc_hd__a21oi_1
XFILLER_122_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11198_ _11198_/A _11198_/B vssd1 vssd1 vccd1 vccd1 _11201_/B sky130_fd_sc_hd__xnor2_1
XFILLER_94_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10149_ _10149_/A _10149_/B vssd1 vssd1 vccd1 vccd1 _10265_/A sky130_fd_sc_hd__nor2_1
XFILLER_48_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14957_ _12054_/A _10993_/D _10657_/C vssd1 vssd1 vccd1 vccd1 _15056_/B sky130_fd_sc_hd__a21o_1
XFILLER_36_946 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13908_ _13908_/A _13908_/B _13908_/C vssd1 vssd1 vccd1 vccd1 _14027_/B sky130_fd_sc_hd__and3_1
X_14888_ _14888_/A _14888_/B _14888_/C _14888_/D vssd1 vssd1 vccd1 vccd1 _15025_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_51_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16627_ _16627_/A _16627_/B vssd1 vssd1 vccd1 vccd1 _16628_/B sky130_fd_sc_hd__xnor2_1
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13839_ _14841_/B _14840_/B _14733_/S vssd1 vssd1 vccd1 vccd1 _13839_/X sky130_fd_sc_hd__mux2_1
XFILLER_62_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16558_ _16558_/A _16558_/B _16558_/C vssd1 vssd1 vccd1 vccd1 _16560_/A sky130_fd_sc_hd__nand3_1
XFILLER_31_640 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15509_ _15510_/A _15510_/B vssd1 vssd1 vccd1 vccd1 _15509_/Y sky130_fd_sc_hd__nor2_1
XFILLER_148_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16489_ _14775_/X _16799_/A2 _16580_/B1 _16480_/A _17162_/C1 vssd1 vssd1 vccd1 vccd1
+ _16489_/X sky130_fd_sc_hd__a221o_1
XFILLER_30_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09030_ _17397_/A _17395_/A _09030_/C _11961_/B vssd1 vssd1 vccd1 vccd1 _09031_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_129_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_918 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09932_ _09932_/A _09932_/B vssd1 vssd1 vccd1 vccd1 _09933_/B sky130_fd_sc_hd__nand2_1
XFILLER_89_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout804 fanout805/X vssd1 vssd1 vccd1 vccd1 _10525_/D sky130_fd_sc_hd__clkbuf_4
Xfanout815 _17488_/Q vssd1 vssd1 vccd1 vccd1 _11281_/B sky130_fd_sc_hd__buf_4
Xfanout826 _12770_/D vssd1 vssd1 vccd1 vccd1 _09267_/D sky130_fd_sc_hd__clkbuf_4
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout837 _17485_/Q vssd1 vssd1 vccd1 vccd1 _12618_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_86_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09863_ _09863_/A _09863_/B _09863_/C vssd1 vssd1 vccd1 vccd1 _09864_/C sky130_fd_sc_hd__nand3_1
Xfanout848 _11437_/D vssd1 vssd1 vccd1 vccd1 _11518_/C sky130_fd_sc_hd__buf_2
XFILLER_100_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_984 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout859 _12295_/D vssd1 vssd1 vccd1 vccd1 _15238_/A sky130_fd_sc_hd__clkbuf_4
X_08814_ _08814_/A _08814_/B vssd1 vssd1 vccd1 vccd1 _08876_/A sky130_fd_sc_hd__xnor2_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09794_ _09639_/C _10203_/B _09640_/A _09638_/Y vssd1 vssd1 vccd1 vccd1 _09795_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_100_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_879 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08745_ _12068_/B _11861_/B _09030_/C _12068_/A vssd1 vssd1 vccd1 vccd1 _08748_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_38_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_935 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09228_ _09228_/A _09228_/B vssd1 vssd1 vccd1 vccd1 _09230_/A sky130_fd_sc_hd__nor2_1
XFILLER_155_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09159_ _11839_/S _11813_/B vssd1 vssd1 vccd1 vccd1 _14948_/B sky130_fd_sc_hd__and2_1
XFILLER_108_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12170_ _12170_/A _12170_/B vssd1 vssd1 vccd1 vccd1 _12172_/A sky130_fd_sc_hd__nor2_1
XFILLER_101_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11121_ _11121_/A _11126_/A _11121_/C vssd1 vssd1 vccd1 vccd1 _11130_/B sky130_fd_sc_hd__or3_1
XFILLER_123_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_567 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11052_ _11047_/Y _11050_/X _11041_/Y _11042_/X vssd1 vssd1 vccd1 vccd1 _11055_/C
+ sky130_fd_sc_hd__o211ai_2
XFILLER_150_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_1044 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_846 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10003_ _10003_/A _10003_/B vssd1 vssd1 vccd1 vccd1 _10005_/B sky130_fd_sc_hd__xnor2_1
X_15860_ _15861_/A _15861_/B vssd1 vssd1 vccd1 vccd1 _15980_/A sky130_fd_sc_hd__and2_1
XFILLER_49_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14811_ _15895_/B _15895_/C _09424_/X vssd1 vssd1 vccd1 vccd1 _16005_/C sky130_fd_sc_hd__a21o_1
XFILLER_76_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15791_ _15788_/Y _15790_/X _16911_/A vssd1 vssd1 vccd1 vccd1 _15791_/Y sky130_fd_sc_hd__o21ai_1
X_17530_ fanout945/X _17530_/D vssd1 vssd1 vccd1 vccd1 _17530_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_91_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11954_ _17409_/A _12320_/D vssd1 vssd1 vccd1 vccd1 _11956_/C sky130_fd_sc_hd__nand2_1
X_14742_ _14742_/A _14742_/B vssd1 vssd1 vccd1 vccd1 _14743_/B sky130_fd_sc_hd__nand2_1
XFILLER_45_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10905_ _10954_/A _11006_/B _10954_/D _10905_/D vssd1 vssd1 vccd1 vccd1 _10907_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_44_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17461_ fanout933/X _17461_/D vssd1 vssd1 vccd1 vccd1 _17461_/Q sky130_fd_sc_hd__dfxtp_2
X_14673_ _17134_/A _14829_/B vssd1 vssd1 vccd1 vccd1 _17167_/A sky130_fd_sc_hd__nand2_4
X_11885_ _11886_/A _11886_/B vssd1 vssd1 vccd1 vccd1 _12118_/A sky130_fd_sc_hd__nand2_1
XFILLER_33_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16412_ _16318_/A _16504_/B _16316_/B vssd1 vssd1 vccd1 vccd1 _16414_/B sky130_fd_sc_hd__o21ai_1
XFILLER_44_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13624_ _14421_/S _13624_/B vssd1 vssd1 vccd1 vccd1 _13624_/X sky130_fd_sc_hd__or2_1
X_10836_ _10836_/A _10850_/A vssd1 vssd1 vccd1 vccd1 _10846_/A sky130_fd_sc_hd__or2_1
XFILLER_60_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17392_ input41/X _17426_/A2 _17391_/X _17426_/C1 vssd1 vssd1 vccd1 vccd1 _17524_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_13_640 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16343_ _16344_/A _16344_/B vssd1 vssd1 vccd1 vccd1 _16345_/A sky130_fd_sc_hd__and2_1
X_13555_ _13555_/A _13555_/B vssd1 vssd1 vccd1 vccd1 _13556_/B sky130_fd_sc_hd__and2_1
XFILLER_13_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10767_ _10766_/C _11725_/A _10667_/Y _10692_/X vssd1 vssd1 vccd1 vccd1 _10774_/A
+ sky130_fd_sc_hd__a211oi_2
XFILLER_34_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_8 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12506_ _12506_/A _12506_/B vssd1 vssd1 vccd1 vccd1 _12508_/C sky130_fd_sc_hd__xnor2_1
XFILLER_12_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16274_ _16181_/A _16279_/C _16180_/B _16160_/X vssd1 vssd1 vccd1 vccd1 _16276_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_145_306 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13486_ _13486_/A _13603_/B _13486_/C vssd1 vssd1 vccd1 vccd1 _13486_/X sky130_fd_sc_hd__and3_1
X_10698_ _11027_/B _11006_/C _10697_/B _10694_/X vssd1 vssd1 vccd1 vccd1 _10701_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_139_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15225_ _15225_/A _15225_/B vssd1 vssd1 vccd1 vccd1 _15226_/B sky130_fd_sc_hd__xnor2_1
X_12437_ _12437_/A _12437_/B _12437_/C vssd1 vssd1 vccd1 vccd1 _12458_/B sky130_fd_sc_hd__nand3_1
XFILLER_126_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15156_ _15157_/A _15157_/B vssd1 vssd1 vccd1 vccd1 _15222_/B sky130_fd_sc_hd__nand2b_1
X_12368_ _12368_/A _12368_/B vssd1 vssd1 vccd1 vccd1 _12370_/A sky130_fd_sc_hd__xnor2_2
XFILLER_126_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14107_ _14108_/A _14108_/B vssd1 vssd1 vccd1 vccd1 _14197_/A sky130_fd_sc_hd__nand2b_1
X_11319_ _11553_/B _11387_/B _11268_/C _11268_/D vssd1 vssd1 vccd1 vccd1 _11320_/C
+ sky130_fd_sc_hd__a22oi_1
XFILLER_5_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15087_ _15161_/A _15087_/B vssd1 vssd1 vccd1 vccd1 _15091_/A sky130_fd_sc_hd__nand2_1
X_12299_ _12299_/A _12299_/B vssd1 vssd1 vccd1 vccd1 _12300_/B sky130_fd_sc_hd__and2_1
XFILLER_99_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14038_ _15457_/A _14036_/X _14037_/X vssd1 vssd1 vccd1 vccd1 _14038_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_68_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_879 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15989_ _15989_/A _15989_/B _15987_/X vssd1 vssd1 vccd1 vccd1 _15990_/B sky130_fd_sc_hd__or3b_1
XFILLER_94_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09013_ _09013_/A _09013_/B vssd1 vssd1 vccd1 vccd1 _09014_/B sky130_fd_sc_hd__nor2_1
XFILLER_129_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1025 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout601 _11630_/A vssd1 vssd1 vccd1 vccd1 _11281_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout612 _17510_/Q vssd1 vssd1 vccd1 vccd1 _10430_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_77_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09915_ _09915_/A _09915_/B vssd1 vssd1 vccd1 vccd1 _09973_/B sky130_fd_sc_hd__or2_1
XFILLER_144_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout623 _17509_/Q vssd1 vssd1 vccd1 vccd1 _08967_/B sky130_fd_sc_hd__buf_4
Xfanout634 _15033_/A3 vssd1 vssd1 vccd1 vccd1 _13037_/B sky130_fd_sc_hd__clkbuf_2
Xfanout645 _17065_/A vssd1 vssd1 vccd1 vccd1 _14641_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_98_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout656 _11813_/B vssd1 vssd1 vccd1 vccd1 _12445_/C sky130_fd_sc_hd__clkbuf_4
Xfanout667 _17503_/Q vssd1 vssd1 vccd1 vccd1 _13704_/B sky130_fd_sc_hd__buf_2
X_09846_ _10244_/A _10255_/B vssd1 vssd1 vccd1 vccd1 _09847_/B sky130_fd_sc_hd__nand2_1
XFILLER_98_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout678 _08860_/B vssd1 vssd1 vccd1 vccd1 _12258_/B sky130_fd_sc_hd__clkbuf_4
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout689 fanout690/X vssd1 vssd1 vccd1 vccd1 _10180_/B sky130_fd_sc_hd__buf_2
XFILLER_100_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09777_ _09777_/A _09777_/B vssd1 vssd1 vccd1 vccd1 _09811_/A sky130_fd_sc_hd__nor2_1
XFILLER_85_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08728_ _15008_/B vssd1 vssd1 vccd1 vccd1 _15553_/A sky130_fd_sc_hd__clkinv_4
XFILLER_2_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_275 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_12 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1018 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11670_ _15524_/C _11690_/A _11670_/C vssd1 vssd1 vccd1 vccd1 _11671_/B sky130_fd_sc_hd__and3b_1
XFILLER_42_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10621_ _10621_/A _10621_/B vssd1 vssd1 vccd1 vccd1 _10716_/B sky130_fd_sc_hd__nor2_1
XFILLER_139_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13340_ _13339_/A _13339_/B _13339_/C vssd1 vssd1 vccd1 vccd1 _13462_/A sky130_fd_sc_hd__o21ai_1
XFILLER_139_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10552_ _10566_/A _10523_/Y _10538_/Y _10550_/X vssd1 vssd1 vccd1 vccd1 _10553_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_155_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13271_ _13271_/A _13271_/B vssd1 vssd1 vccd1 vccd1 _13386_/B sky130_fd_sc_hd__or2_1
XFILLER_155_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10483_ _10597_/A _10597_/B vssd1 vssd1 vccd1 vccd1 _10497_/A sky130_fd_sc_hd__nand2_1
XFILLER_136_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15010_ _11651_/A _15008_/A _15008_/B _14794_/A vssd1 vssd1 vccd1 vccd1 _15011_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_108_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12222_ _12220_/X _12221_/X _17367_/A vssd1 vssd1 vccd1 vccd1 _12222_/X sky130_fd_sc_hd__mux2_1
XFILLER_170_618 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12153_ _11917_/X _11947_/X _12316_/B _12152_/X vssd1 vssd1 vccd1 vccd1 _12360_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_64_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1019 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11104_ _11104_/A _11104_/B _11104_/C vssd1 vssd1 vccd1 vccd1 _11105_/B sky130_fd_sc_hd__nand3_1
XFILLER_2_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16961_ _16931_/X _16932_/X _16960_/X vssd1 vssd1 vccd1 vccd1 _17014_/A sky130_fd_sc_hd__a21o_1
X_12084_ _12085_/A _12085_/B _12085_/C vssd1 vssd1 vccd1 vccd1 _12268_/A sky130_fd_sc_hd__a21o_1
XFILLER_111_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_386 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11035_ _11035_/A _11035_/B vssd1 vssd1 vccd1 vccd1 _11038_/A sky130_fd_sc_hd__xor2_1
X_15912_ _16809_/C _16129_/B vssd1 vssd1 vccd1 vccd1 _16939_/B sky130_fd_sc_hd__nand2_2
XFILLER_49_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16892_ _16827_/A _16827_/C _16758_/B _16935_/A vssd1 vssd1 vccd1 vccd1 _16893_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_49_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15843_ _16807_/A _16054_/B vssd1 vssd1 vccd1 vccd1 _16355_/B sky130_fd_sc_hd__and2_2
XFILLER_77_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12986_ _12985_/A _12985_/B _12985_/C vssd1 vssd1 vccd1 vccd1 _12986_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_94_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15774_ _16281_/A _16065_/B vssd1 vssd1 vccd1 vccd1 _15775_/B sky130_fd_sc_hd__nand2_1
XTAP_3561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17513_ fanout949/X _17513_/D vssd1 vssd1 vccd1 vccd1 _17513_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14725_ _14727_/B vssd1 vssd1 vccd1 vccd1 _14725_/Y sky130_fd_sc_hd__inv_2
XTAP_3594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11937_ _11937_/A _11937_/B vssd1 vssd1 vccd1 vccd1 _11939_/A sky130_fd_sc_hd__xnor2_1
XTAP_2860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17444_ fanout938/X _17444_/D vssd1 vssd1 vccd1 vccd1 _17444_/Q sky130_fd_sc_hd__dfxtp_1
X_11868_ _11868_/A _12093_/A vssd1 vssd1 vccd1 vccd1 _11871_/A sky130_fd_sc_hd__nor2_1
X_14656_ _14691_/A _14656_/B vssd1 vssd1 vccd1 vccd1 _14658_/C sky130_fd_sc_hd__and2_1
XFILLER_32_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10819_ _11095_/A _11095_/B _17468_/D _11240_/C vssd1 vssd1 vccd1 vccd1 _10822_/A
+ sky130_fd_sc_hd__and4_1
X_13607_ _13607_/A _13607_/B _13607_/C vssd1 vssd1 vccd1 vccd1 _13607_/X sky130_fd_sc_hd__or3_1
XFILLER_60_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17375_ _17375_/A _17389_/B vssd1 vssd1 vccd1 vccd1 _17375_/X sky130_fd_sc_hd__or2_1
X_14587_ _14629_/C _14587_/B vssd1 vssd1 vccd1 vccd1 _14587_/Y sky130_fd_sc_hd__nand2_1
X_11799_ _14888_/C _11799_/B vssd1 vssd1 vccd1 vccd1 _11800_/D sky130_fd_sc_hd__or2_1
XFILLER_159_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16326_ _16326_/A _16326_/B vssd1 vssd1 vccd1 vccd1 _16328_/B sky130_fd_sc_hd__xor2_1
X_13538_ _13538_/A _13538_/B vssd1 vssd1 vccd1 vccd1 _13543_/A sky130_fd_sc_hd__xnor2_1
XFILLER_146_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16257_ _16257_/A _16257_/B vssd1 vssd1 vccd1 vccd1 _16273_/A sky130_fd_sc_hd__xor2_1
X_13469_ _13469_/A _13469_/B vssd1 vssd1 vccd1 vccd1 _13471_/A sky130_fd_sc_hd__nor2_1
XFILLER_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15208_ _15208_/A _15262_/C _15208_/C _15208_/D vssd1 vssd1 vccd1 vccd1 _15208_/X
+ sky130_fd_sc_hd__or4_2
XFILLER_160_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16188_ _16188_/A _16188_/B _16188_/C vssd1 vssd1 vccd1 vccd1 _16189_/B sky130_fd_sc_hd__nor3_1
XFILLER_127_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15139_ _15147_/A _17614_/Q _15147_/C vssd1 vssd1 vccd1 vccd1 _15270_/B sky130_fd_sc_hd__nor3_2
XFILLER_88_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09700_ _10244_/A _10508_/D _09701_/C vssd1 vssd1 vccd1 vccd1 _09702_/A sky130_fd_sc_hd__a21oi_1
XFILLER_96_952 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09631_ _09632_/B _09632_/A vssd1 vssd1 vccd1 vccd1 _09631_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_95_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_635 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09562_ _09556_/A _09558_/B _09556_/B vssd1 vssd1 vccd1 vccd1 _09565_/A sky130_fd_sc_hd__o21ba_1
XFILLER_82_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09493_ _09493_/A _11813_/B _14949_/A vssd1 vssd1 vccd1 vccd1 _09619_/B sky130_fd_sc_hd__and3_1
XFILLER_24_724 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_607 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_919 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout420 _17529_/Q vssd1 vssd1 vccd1 vccd1 _10111_/C sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout431 _12722_/A vssd1 vssd1 vccd1 vccd1 _13641_/A sky130_fd_sc_hd__buf_2
XFILLER_120_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout442 _10242_/A1 vssd1 vssd1 vccd1 vccd1 _16209_/C sky130_fd_sc_hd__clkbuf_4
Xfanout453 _09412_/A vssd1 vssd1 vccd1 vccd1 _10244_/A sky130_fd_sc_hd__clkbuf_4
Xfanout464 _17524_/Q vssd1 vssd1 vccd1 vccd1 _14873_/B sky130_fd_sc_hd__buf_4
Xfanout475 _17522_/Q vssd1 vssd1 vccd1 vccd1 _13302_/A sky130_fd_sc_hd__buf_6
Xfanout486 _10142_/A vssd1 vssd1 vccd1 vccd1 _11095_/A sky130_fd_sc_hd__buf_2
XFILLER_171_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout497 _17520_/Q vssd1 vssd1 vccd1 vccd1 _09299_/B sky130_fd_sc_hd__buf_6
X_09829_ _09813_/A _09813_/C _09813_/B vssd1 vssd1 vccd1 vccd1 _09829_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_86_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12840_ _12838_/Y _12840_/B vssd1 vssd1 vccd1 vccd1 _13003_/B sky130_fd_sc_hd__nand2b_1
XFILLER_62_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_668 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12771_ _12771_/A _12771_/B vssd1 vssd1 vccd1 vccd1 _12773_/A sky130_fd_sc_hd__nor2_1
XTAP_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11722_ _11722_/A _11722_/B vssd1 vssd1 vccd1 vccd1 _11731_/A sky130_fd_sc_hd__nor2_1
X_14510_ _14512_/A vssd1 vssd1 vccd1 vccd1 _14579_/A sky130_fd_sc_hd__inv_2
XTAP_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15490_ _08731_/A _15208_/C _15208_/A vssd1 vssd1 vccd1 vccd1 _15492_/B sky130_fd_sc_hd__a21bo_1
XTAP_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_885 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11653_ _15056_/A _11653_/B vssd1 vssd1 vccd1 vccd1 _11655_/A sky130_fd_sc_hd__nor2_2
XTAP_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14441_ _14441_/A _14441_/B vssd1 vssd1 vccd1 vccd1 _14443_/A sky130_fd_sc_hd__nor2_1
XTAP_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10604_ _11006_/A _10904_/A _10703_/B _11005_/B vssd1 vssd1 vccd1 vccd1 _10607_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_70_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14372_ _14372_/A _14372_/B _14372_/C vssd1 vssd1 vccd1 vccd1 _14373_/B sky130_fd_sc_hd__or3_1
X_17160_ _11932_/B _17140_/B _17140_/A vssd1 vssd1 vccd1 vccd1 _17160_/Y sky130_fd_sc_hd__a21oi_1
X_11584_ _11584_/A _11584_/B _11583_/Y vssd1 vssd1 vccd1 vccd1 _11586_/B sky130_fd_sc_hd__nor3b_1
XFILLER_7_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13323_ _14215_/A _13551_/D vssd1 vssd1 vccd1 vccd1 _13324_/B sky130_fd_sc_hd__nand2_1
X_16111_ _16111_/A _16111_/B _16111_/C vssd1 vssd1 vccd1 vccd1 _16111_/X sky130_fd_sc_hd__or3_1
X_10535_ _10535_/A _10644_/A vssd1 vssd1 vccd1 vccd1 _10637_/A sky130_fd_sc_hd__or2_1
X_17091_ _17091_/A _17118_/B vssd1 vssd1 vccd1 vccd1 _17092_/B sky130_fd_sc_hd__or2_1
XFILLER_156_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_978 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_478 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16042_ _16667_/A _16041_/B _16041_/C vssd1 vssd1 vccd1 vccd1 _16043_/B sky130_fd_sc_hd__o21ai_1
XFILLER_129_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13254_ _13118_/A _13119_/Y _13252_/A _13253_/Y vssd1 vssd1 vccd1 vccd1 _13256_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_170_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10466_ _10469_/A _10469_/B _10469_/C vssd1 vssd1 vccd1 vccd1 _10470_/A sky130_fd_sc_hd__o21a_1
XFILLER_136_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12205_ _12010_/A _12010_/B _12006_/X vssd1 vssd1 vccd1 vccd1 _12206_/C sky130_fd_sc_hd__a21oi_1
XFILLER_89_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13185_ _13186_/A _13186_/B vssd1 vssd1 vccd1 vccd1 _13326_/B sky130_fd_sc_hd__nor2_1
XFILLER_151_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10397_ _10397_/A _10397_/B vssd1 vssd1 vccd1 vccd1 _10501_/A sky130_fd_sc_hd__xnor2_1
XFILLER_43_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12136_ _12136_/A _12136_/B vssd1 vssd1 vccd1 vccd1 _12138_/C sky130_fd_sc_hd__nor2_1
XFILLER_69_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16944_ _16994_/B _16944_/B vssd1 vssd1 vccd1 vccd1 _16947_/A sky130_fd_sc_hd__nand2_1
X_12067_ _12068_/B _13208_/D _12942_/D _12068_/A vssd1 vssd1 vccd1 vccd1 _12070_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_49_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11018_ _11018_/A _11018_/B vssd1 vssd1 vccd1 vccd1 _11020_/B sky130_fd_sc_hd__nor2_1
X_16875_ _16917_/A _16862_/X _16863_/Y _16874_/X vssd1 vssd1 vccd1 vccd1 _16875_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_92_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15826_ _15827_/A _15827_/B vssd1 vssd1 vccd1 vccd1 _15826_/Y sky130_fd_sc_hd__nor2_1
XFILLER_93_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15757_ _15668_/A _15668_/B _15665_/Y vssd1 vssd1 vccd1 vccd1 _15759_/B sky130_fd_sc_hd__o21a_1
XTAP_3391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12969_ _12805_/A _12807_/B _12805_/B vssd1 vssd1 vccd1 vccd1 _12971_/B sky130_fd_sc_hd__o21ba_1
XFILLER_61_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14708_ _14738_/A _14708_/B _14738_/B _14708_/D vssd1 vssd1 vccd1 vccd1 _14713_/B
+ sky130_fd_sc_hd__nand4_1
XTAP_2690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15688_ _16281_/A _16589_/B _15686_/Y vssd1 vssd1 vccd1 vccd1 _15689_/B sky130_fd_sc_hd__a21o_1
XFILLER_61_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17427_ input28/X input29/X wire215/X vssd1 vssd1 vccd1 vccd1 _17428_/D sky130_fd_sc_hd__a21boi_1
XFILLER_60_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14639_ _14641_/B _14641_/C _14641_/D _14641_/A vssd1 vssd1 vccd1 vccd1 _14642_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_159_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17358_ _12592_/D _17360_/A2 _17357_/X _17358_/C1 vssd1 vssd1 vccd1 vccd1 _17508_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_158_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16309_ _17143_/A1 _13943_/X _14926_/X _14990_/X vssd1 vssd1 vccd1 vccd1 _16310_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_9_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17289_ _17573_/Q _17289_/B vssd1 vssd1 vccd1 vccd1 _17289_/X sky130_fd_sc_hd__and2_1
XFILLER_162_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1025 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_824 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08993_ _09493_/A _11932_/B _08993_/C vssd1 vssd1 vccd1 vccd1 _08994_/B sky130_fd_sc_hd__and3_1
XFILLER_88_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09614_ _09614_/A _09614_/B vssd1 vssd1 vccd1 vccd1 _09746_/C sky130_fd_sc_hd__xnor2_1
XFILLER_28_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09545_ _09577_/A _09577_/B vssd1 vssd1 vccd1 vccd1 _09596_/A sky130_fd_sc_hd__nand2_1
XFILLER_43_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09476_ _09478_/B _09603_/A _09478_/A vssd1 vssd1 vccd1 vccd1 _09476_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_24_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_935 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10320_ _10319_/A _10319_/Y _10193_/B _10229_/X vssd1 vssd1 vccd1 vccd1 _10336_/A
+ sky130_fd_sc_hd__a211oi_2
XFILLER_109_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10251_ _10251_/A _10251_/B vssd1 vssd1 vccd1 vccd1 _10253_/B sky130_fd_sc_hd__xnor2_1
XFILLER_117_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10182_ _10183_/A _10181_/Y _10182_/C _10309_/B vssd1 vssd1 vccd1 vccd1 _10307_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_120_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_708 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14990_ _15537_/B _14989_/X _15901_/S vssd1 vssd1 vccd1 vccd1 _14990_/X sky130_fd_sc_hd__mux2_1
Xfanout250 _14836_/Y vssd1 vssd1 vccd1 vccd1 _15456_/B sky130_fd_sc_hd__buf_2
Xfanout261 _17355_/C vssd1 vssd1 vccd1 vccd1 _17353_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_87_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout272 _14939_/X vssd1 vssd1 vccd1 vccd1 _17134_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_13941_ _14122_/A wire116/X vssd1 vssd1 vccd1 vccd1 _14032_/B sky130_fd_sc_hd__nor2_1
Xfanout283 _17363_/A vssd1 vssd1 vccd1 vccd1 _12054_/A sky130_fd_sc_hd__clkbuf_4
Xfanout294 fanout299/X vssd1 vssd1 vccd1 vccd1 _12865_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_74_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16660_ _16651_/A _16806_/A2 _16659_/X vssd1 vssd1 vccd1 vccd1 _17564_/D sky130_fd_sc_hd__a21oi_1
X_13872_ _13873_/A _13873_/B vssd1 vssd1 vccd1 vccd1 _14018_/A sky130_fd_sc_hd__nand2_1
XFILLER_74_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15611_ _15522_/A _15521_/B _15519_/X vssd1 vssd1 vccd1 vccd1 _15611_/X sky130_fd_sc_hd__a21o_1
XFILLER_28_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12823_ _12822_/B _12823_/B vssd1 vssd1 vccd1 vccd1 _12824_/B sky130_fd_sc_hd__nand2b_1
XFILLER_74_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16591_ _16814_/B _16591_/B _16591_/C vssd1 vssd1 vccd1 vccd1 _16686_/B sky130_fd_sc_hd__and3_1
XFILLER_61_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15542_ _14785_/X _16008_/A2 _15713_/B1 _15541_/A _16869_/C1 vssd1 vssd1 vccd1 vccd1
+ _15542_/X sky130_fd_sc_hd__a221o_1
X_12754_ _12754_/A _12754_/B vssd1 vssd1 vccd1 vccd1 _12755_/C sky130_fd_sc_hd__xnor2_1
XFILLER_43_863 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11705_ _11705_/A _15888_/A vssd1 vssd1 vccd1 vccd1 _11705_/Y sky130_fd_sc_hd__nand2_1
XFILLER_30_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15473_ _16127_/A _16152_/A _16604_/B _15475_/A vssd1 vssd1 vccd1 vccd1 _15473_/X
+ sky130_fd_sc_hd__a22o_1
X_12685_ _12685_/A _12685_/B vssd1 vssd1 vccd1 vccd1 _12685_/Y sky130_fd_sc_hd__nand2_1
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17212_ _17438_/Q _17275_/A2 _17210_/X _17211_/X _17364_/C1 vssd1 vssd1 vccd1 vccd1
+ _17438_/D sky130_fd_sc_hd__o221a_1
X_11636_ _15116_/A _11653_/B _15553_/A _15175_/A vssd1 vssd1 vccd1 vccd1 _11637_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_30_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14424_ _14424_/A _14424_/B vssd1 vssd1 vccd1 vccd1 _14469_/A sky130_fd_sc_hd__nor2_1
XFILLER_168_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17143_ _17143_/A1 _14734_/B _17142_/X vssd1 vssd1 vccd1 vccd1 _17143_/X sky130_fd_sc_hd__o21a_1
XFILLER_156_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11567_ _11558_/A _11558_/C _11558_/B vssd1 vssd1 vccd1 vccd1 _11568_/C sky130_fd_sc_hd__a21o_1
X_14355_ _14763_/S _14353_/Y _14354_/X _14288_/Y vssd1 vssd1 vccd1 vccd1 _17596_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_10_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10518_ _10384_/X _10475_/Y _10485_/X _10499_/A vssd1 vssd1 vccd1 vccd1 _10519_/C
+ sky130_fd_sc_hd__o211a_1
X_13306_ _13306_/A _13306_/B vssd1 vssd1 vccd1 vccd1 _13308_/C sky130_fd_sc_hd__xnor2_1
X_14286_ _12545_/X _12553_/B _14356_/S vssd1 vssd1 vccd1 vccd1 _16653_/B sky130_fd_sc_hd__mux2_1
X_17074_ _14765_/X _17162_/A2 _16974_/B _17065_/A _17162_/C1 vssd1 vssd1 vccd1 vccd1
+ _17074_/X sky130_fd_sc_hd__a221o_1
X_11498_ _11495_/A _11495_/B _11532_/A vssd1 vssd1 vccd1 vccd1 _11499_/C sky130_fd_sc_hd__o21ba_1
XFILLER_144_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16025_ _16025_/A _16813_/B vssd1 vssd1 vccd1 vccd1 _16026_/B sky130_fd_sc_hd__nor2_1
X_13237_ _13238_/A _13238_/B vssd1 vssd1 vccd1 vccd1 _13366_/A sky130_fd_sc_hd__or2_1
X_10449_ _10563_/A _10563_/B vssd1 vssd1 vccd1 vccd1 _10564_/A sky130_fd_sc_hd__nand2_1
XFILLER_124_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13168_ _13414_/B _13846_/B _14008_/B _13658_/A vssd1 vssd1 vccd1 vccd1 _13170_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_152_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12119_ _11905_/X _11909_/A _12309_/A _12118_/Y vssd1 vssd1 vccd1 vccd1 _12309_/B
+ sky130_fd_sc_hd__o211ai_4
X_13099_ _13099_/A _13099_/B vssd1 vssd1 vccd1 vccd1 _13101_/A sky130_fd_sc_hd__nor2_1
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16927_ _17164_/C _15537_/X _16926_/Y vssd1 vssd1 vccd1 vccd1 _16927_/X sky130_fd_sc_hd__o21a_1
XFILLER_66_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16858_ _14383_/A _16965_/B _16859_/A vssd1 vssd1 vccd1 vccd1 _16858_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_37_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15809_ _15805_/Y _15806_/Y _15808_/Y vssd1 vssd1 vccd1 vccd1 _15809_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_37_189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16789_ _16789_/A _17153_/B vssd1 vssd1 vccd1 vccd1 _16789_/Y sky130_fd_sc_hd__nor2_1
XFILLER_92_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09330_ _09462_/A _09468_/A _09462_/C vssd1 vssd1 vccd1 vccd1 _09463_/A sky130_fd_sc_hd__o21ai_1
XFILLER_21_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09261_ _09261_/A _09261_/B vssd1 vssd1 vccd1 vccd1 _09310_/A sky130_fd_sc_hd__nand2_1
XFILLER_21_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09192_ _09514_/B _12174_/D _12129_/B _09942_/A vssd1 vssd1 vccd1 vccd1 _09194_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_119_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_982 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_610 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08976_ _12770_/A _17423_/A _09362_/D _09172_/B vssd1 vssd1 vccd1 vccd1 _09238_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_152_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_774 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09528_ _09391_/C _09399_/Y _09458_/X _09628_/A vssd1 vssd1 vccd1 vccd1 _09528_/Y
+ sky130_fd_sc_hd__a211oi_1
XFILLER_169_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09459_ _09334_/A _09334_/B _09334_/C vssd1 vssd1 vccd1 vccd1 _09459_/Y sky130_fd_sc_hd__a21oi_1
XPHY_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12470_ _12303_/A _12470_/B vssd1 vssd1 vccd1 vccd1 _12471_/C sky130_fd_sc_hd__nand2b_1
XFILLER_8_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_732 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11421_ _11396_/A _11396_/C _11396_/B vssd1 vssd1 vccd1 vccd1 _11421_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_137_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14140_ _14708_/B _16651_/A _14141_/D _14290_/A vssd1 vssd1 vccd1 vccd1 _14142_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_165_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11352_ _11352_/A _11352_/B vssd1 vssd1 vccd1 vccd1 _11354_/B sky130_fd_sc_hd__xnor2_1
XFILLER_4_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_595 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10303_ _10305_/B _10305_/C _10305_/A vssd1 vssd1 vccd1 vccd1 _10303_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_3_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14071_ _14071_/A _14071_/B vssd1 vssd1 vccd1 vccd1 _14074_/A sky130_fd_sc_hd__xor2_1
X_11283_ _11283_/A _11283_/B _11333_/A vssd1 vssd1 vccd1 vccd1 _11284_/B sky130_fd_sc_hd__or3_1
X_13022_ _13846_/A _12871_/B _12872_/A _12870_/B vssd1 vssd1 vccd1 vccd1 _13024_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_3_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10234_ _10234_/A _10234_/B vssd1 vssd1 vccd1 vccd1 _10246_/A sky130_fd_sc_hd__nor2_1
XFILLER_10_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_60 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10165_ _14787_/A _10647_/D _10745_/D _14786_/A vssd1 vssd1 vccd1 vccd1 _10165_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_120_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14973_ _14886_/X _14972_/X _15056_/A vssd1 vssd1 vccd1 vccd1 _14973_/Y sky130_fd_sc_hd__a21oi_1
X_10096_ _09968_/B _09970_/A _09968_/A vssd1 vssd1 vccd1 vccd1 _11778_/B sky130_fd_sc_hd__o21ai_1
XFILLER_59_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16712_ _16786_/A _16712_/B vssd1 vssd1 vccd1 vccd1 _16714_/B sky130_fd_sc_hd__and2_1
X_13924_ _13925_/A _13925_/B _13925_/C vssd1 vssd1 vccd1 vccd1 _14030_/A sky130_fd_sc_hd__a21o_1
XFILLER_47_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_903 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16643_ _16643_/A vssd1 vssd1 vccd1 vccd1 _16643_/Y sky130_fd_sc_hd__inv_2
X_13855_ _13856_/A _13856_/B vssd1 vssd1 vccd1 vccd1 _13961_/A sky130_fd_sc_hd__and2b_1
XFILLER_34_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12806_ _17415_/A _13434_/D vssd1 vssd1 vccd1 vccd1 _12807_/B sky130_fd_sc_hd__nand2_1
X_16574_ _16917_/A _16574_/B vssd1 vssd1 vccd1 vccd1 _16574_/Y sky130_fd_sc_hd__nand2_1
X_10998_ _11159_/A _10998_/B vssd1 vssd1 vccd1 vccd1 _10999_/C sky130_fd_sc_hd__and2_1
X_13786_ _13787_/A _13787_/B vssd1 vssd1 vccd1 vccd1 _13915_/A sky130_fd_sc_hd__and2b_1
XFILLER_163_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15525_ _15525_/A _15525_/B vssd1 vssd1 vccd1 vccd1 _15525_/X sky130_fd_sc_hd__and2_1
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12737_ _12737_/A _12737_/B vssd1 vssd1 vccd1 vccd1 _12739_/B sky130_fd_sc_hd__xnor2_1
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15456_ _15456_/A _15456_/B _15455_/X vssd1 vssd1 vccd1 vccd1 _15467_/B sky130_fd_sc_hd__or3b_1
XFILLER_124_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12668_ _12668_/A _12668_/B vssd1 vssd1 vccd1 vccd1 _12669_/B sky130_fd_sc_hd__nand2_1
XFILLER_30_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14407_ _14340_/B _14342_/A _14424_/B _14406_/Y vssd1 vssd1 vccd1 vccd1 _14473_/A
+ sky130_fd_sc_hd__a211o_1
X_11619_ _11584_/A _11584_/B _11583_/Y vssd1 vssd1 vccd1 vccd1 _11620_/C sky130_fd_sc_hd__o21ba_1
XFILLER_128_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15387_ _16015_/A _15463_/B _15381_/Y _15383_/X _15386_/Y vssd1 vssd1 vccd1 vccd1
+ _15387_/X sky130_fd_sc_hd__o311a_1
XFILLER_117_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12599_ _12599_/A _12599_/B vssd1 vssd1 vccd1 vccd1 _12755_/B sky130_fd_sc_hd__and2_1
XFILLER_156_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17126_ _17127_/A _17127_/B vssd1 vssd1 vccd1 vccd1 _17128_/A sky130_fd_sc_hd__or2_1
XFILLER_116_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14338_ _14222_/A _14265_/B _14336_/X _14337_/Y vssd1 vssd1 vccd1 vccd1 _14340_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_116_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17057_ _17056_/B _17057_/B vssd1 vssd1 vccd1 vccd1 _17058_/B sky130_fd_sc_hd__and2b_1
X_14269_ _14270_/A _14270_/B _14270_/C vssd1 vssd1 vccd1 vccd1 _14350_/A sky130_fd_sc_hd__a21oi_1
X_16008_ _16005_/B _16008_/A2 _16008_/B1 _16014_/A _16494_/B1 vssd1 vssd1 vccd1 vccd1
+ _16008_/X sky130_fd_sc_hd__a221o_1
XFILLER_83_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08830_ _08830_/A _08869_/B vssd1 vssd1 vccd1 vccd1 _08832_/B sky130_fd_sc_hd__nand2_1
XFILLER_111_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08761_ _12077_/A _13208_/D vssd1 vssd1 vccd1 vccd1 _16302_/A sky130_fd_sc_hd__nand2_4
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09313_ _09338_/A _09338_/B vssd1 vssd1 vccd1 vccd1 _09391_/B sky130_fd_sc_hd__or2_1
XFILLER_40_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09244_ _09245_/A _09245_/B _09245_/C vssd1 vssd1 vccd1 vccd1 _11990_/B sky130_fd_sc_hd__a21o_1
XFILLER_22_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_354 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09175_ _09357_/A _09174_/Y _09502_/A _10067_/B vssd1 vssd1 vccd1 vccd1 _09364_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_119_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08959_ _08959_/A _08959_/B vssd1 vssd1 vccd1 vccd1 _09077_/B sky130_fd_sc_hd__xnor2_1
XFILLER_102_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11970_ _11970_/A _11970_/B vssd1 vssd1 vccd1 vccd1 _11971_/B sky130_fd_sc_hd__nand2_1
XFILLER_56_67 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10921_ _14786_/A _15463_/A vssd1 vssd1 vccd1 vccd1 _14805_/A sky130_fd_sc_hd__nand2_1
X_10852_ _10851_/B _10971_/B _14895_/B _10933_/A vssd1 vssd1 vccd1 vccd1 _10852_/Y
+ sky130_fd_sc_hd__a22oi_1
X_13640_ _13745_/B _13844_/C _13846_/B _13641_/A vssd1 vssd1 vccd1 vccd1 _13642_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_72_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13571_ _13571_/A _13702_/A vssd1 vssd1 vccd1 vccd1 _13572_/C sky130_fd_sc_hd__and2_1
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10783_ _10784_/A _10784_/B _11768_/B vssd1 vssd1 vccd1 vccd1 _11767_/B sky130_fd_sc_hd__o21ba_1
XFILLER_24_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15310_ _14801_/A _14801_/B _14801_/C vssd1 vssd1 vccd1 vccd1 _15311_/B sky130_fd_sc_hd__o21a_1
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12522_ _12522_/A _12522_/B _12522_/C vssd1 vssd1 vccd1 vccd1 _12524_/A sky130_fd_sc_hd__or3_1
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16290_ _16290_/A _16290_/B _16290_/C vssd1 vssd1 vccd1 vccd1 _16562_/C sky130_fd_sc_hd__or3_1
XFILLER_8_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15241_ _15241_/A _15241_/B _15241_/C vssd1 vssd1 vccd1 vccd1 _15242_/C sky130_fd_sc_hd__nand3_1
X_12453_ _12454_/A _12454_/B _12454_/C vssd1 vssd1 vccd1 vccd1 _12626_/A sky130_fd_sc_hd__a21o_1
X_11404_ _11406_/A _11406_/B vssd1 vssd1 vccd1 vccd1 _11405_/A sky130_fd_sc_hd__or2_1
XFILLER_166_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15172_ _15106_/A _11683_/B _15998_/A vssd1 vssd1 vccd1 vccd1 _15173_/B sky130_fd_sc_hd__a21oi_1
X_12384_ _12382_/X _12383_/X _12865_/S vssd1 vssd1 vccd1 vccd1 _12384_/X sky130_fd_sc_hd__mux2_1
XFILLER_126_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11335_ _11520_/C _15208_/A vssd1 vssd1 vccd1 vccd1 _11386_/A sky130_fd_sc_hd__nand2_1
XFILLER_125_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14123_ _13939_/Y _14281_/A _14121_/X vssd1 vssd1 vccd1 vccd1 _14125_/B sky130_fd_sc_hd__a21oi_1
XFILLER_21_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1028 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11266_ _11427_/A _11553_/A _11437_/D _11561_/C vssd1 vssd1 vccd1 vccd1 _11268_/C
+ sky130_fd_sc_hd__nand4_1
X_14054_ _14054_/A _14054_/B vssd1 vssd1 vccd1 vccd1 _14055_/B sky130_fd_sc_hd__and2_1
XFILLER_141_749 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13005_ _13005_/A _13005_/B vssd1 vssd1 vccd1 vccd1 _13005_/X sky130_fd_sc_hd__and2_1
XFILLER_79_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10217_ _10209_/A _10210_/A _10209_/B _10211_/Y vssd1 vssd1 vccd1 vccd1 _10219_/B
+ sky130_fd_sc_hd__o31a_1
X_11197_ _11198_/B _11198_/A vssd1 vssd1 vccd1 vccd1 _11229_/A sky130_fd_sc_hd__and2b_1
XFILLER_67_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10148_ _10148_/A _10148_/B _10148_/C vssd1 vssd1 vccd1 vccd1 _10149_/B sky130_fd_sc_hd__nor3_1
XFILLER_48_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10079_ _10080_/A _10080_/B vssd1 vssd1 vccd1 vccd1 _10081_/A sky130_fd_sc_hd__nand2_1
X_14956_ _14956_/A _14956_/B vssd1 vssd1 vccd1 vccd1 _14956_/Y sky130_fd_sc_hd__nor2_1
XFILLER_36_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13907_ _14027_/A _13907_/B vssd1 vssd1 vccd1 vccd1 _13908_/C sky130_fd_sc_hd__nor2_1
XFILLER_35_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14887_ _14888_/A _14887_/B vssd1 vssd1 vccd1 vccd1 _14887_/Y sky130_fd_sc_hd__nor2_1
X_16626_ _16624_/X _16626_/B vssd1 vssd1 vccd1 vccd1 _16627_/B sky130_fd_sc_hd__and2b_1
XFILLER_35_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13838_ _12857_/X _12861_/X _17369_/A vssd1 vssd1 vccd1 vccd1 _14840_/B sky130_fd_sc_hd__mux2_1
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16557_ _16557_/A _16557_/B _16557_/C vssd1 vssd1 vccd1 vccd1 _16558_/C sky130_fd_sc_hd__or3_1
X_13769_ _13770_/A _13770_/B _13770_/C vssd1 vssd1 vccd1 vccd1 _13921_/A sky130_fd_sc_hd__o21ai_1
XFILLER_43_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15508_ _15687_/A _15755_/B vssd1 vssd1 vccd1 vccd1 _15510_/B sky130_fd_sc_hd__or2_1
X_16488_ _16480_/A _16400_/B _16487_/Y vssd1 vssd1 vccd1 vccd1 _16492_/A sky130_fd_sc_hd__o21ai_1
XFILLER_31_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15439_ _15439_/A _15439_/B vssd1 vssd1 vccd1 vccd1 _15442_/A sky130_fd_sc_hd__xor2_1
XFILLER_163_307 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17109_ _17140_/A _17139_/B _17109_/C vssd1 vssd1 vccd1 vccd1 _17113_/A sky130_fd_sc_hd__or3_1
XFILLER_116_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09931_ _10074_/A _10074_/B vssd1 vssd1 vccd1 vccd1 _10075_/A sky130_fd_sc_hd__or2_1
XFILLER_104_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout805 _17489_/Q vssd1 vssd1 vccd1 vccd1 fanout805/X sky130_fd_sc_hd__clkbuf_4
Xfanout816 _12338_/C vssd1 vssd1 vccd1 vccd1 _09555_/D sky130_fd_sc_hd__buf_4
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout827 _12770_/D vssd1 vssd1 vccd1 vccd1 _09843_/C sky130_fd_sc_hd__clkbuf_4
X_09862_ _09862_/A _09862_/B vssd1 vssd1 vccd1 vccd1 _09864_/B sky130_fd_sc_hd__xnor2_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout838 _14850_/A vssd1 vssd1 vccd1 vccd1 _15381_/A sky130_fd_sc_hd__buf_4
Xfanout849 _14849_/A vssd1 vssd1 vccd1 vccd1 _11437_/D sky130_fd_sc_hd__buf_2
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08813_ _17393_/A _10297_/D vssd1 vssd1 vccd1 vccd1 _08814_/B sky130_fd_sc_hd__nand2_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09793_ _09793_/A _09793_/B vssd1 vssd1 vccd1 vccd1 _09805_/A sky130_fd_sc_hd__nor2_1
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08744_ _15071_/A _08743_/A _08743_/Y vssd1 vssd1 vccd1 vccd1 _17611_/D sky130_fd_sc_hd__a21o_1
XFILLER_38_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_796 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_1044 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_112 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09227_ _09227_/A _09227_/B _09227_/C vssd1 vssd1 vccd1 vccd1 _09228_/B sky130_fd_sc_hd__and3_1
XFILLER_166_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09158_ _09165_/A _09165_/B vssd1 vssd1 vccd1 vccd1 _09168_/A sky130_fd_sc_hd__nor2_1
XFILLER_163_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09089_ _09317_/A _09323_/A _09317_/C vssd1 vssd1 vccd1 vccd1 _09318_/A sky130_fd_sc_hd__o21ai_1
XFILLER_162_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11120_ _11121_/A _11121_/C vssd1 vssd1 vccd1 vccd1 _11126_/B sky130_fd_sc_hd__nor2_1
XFILLER_107_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11051_ _11051_/A _11051_/B _11051_/C vssd1 vssd1 vccd1 vccd1 _11061_/A sky130_fd_sc_hd__nand3_1
XFILLER_67_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10002_ _10003_/B _10003_/A vssd1 vssd1 vccd1 vccd1 _10009_/B sky130_fd_sc_hd__nand2b_1
XFILLER_88_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14810_ _15801_/B _15802_/A _16809_/B vssd1 vssd1 vccd1 vccd1 _15895_/C sky130_fd_sc_hd__a21o_1
X_15790_ _15610_/Y _15611_/X _15700_/A _15789_/X vssd1 vssd1 vccd1 vccd1 _15790_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_45_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_571 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14741_ _14742_/A _14742_/B vssd1 vssd1 vccd1 vccd1 _14743_/A sky130_fd_sc_hd__or2_1
X_11953_ _17413_/A _17411_/A _12158_/D _12923_/D vssd1 vssd1 vccd1 vccd1 _12163_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_57_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10904_ _10904_/A _11005_/A _17467_/D _11095_/D vssd1 vssd1 vccd1 vccd1 _11107_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_45_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17460_ fanout934/X _17460_/D vssd1 vssd1 vccd1 vccd1 _17460_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_83_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14672_ _14633_/A _14631_/A _14669_/B _14671_/X vssd1 vssd1 vccd1 vccd1 _14701_/A
+ sky130_fd_sc_hd__a31oi_2
X_11884_ _11884_/A _11884_/B vssd1 vssd1 vccd1 vccd1 _11886_/B sky130_fd_sc_hd__xnor2_1
X_16411_ _16411_/A _16505_/B vssd1 vssd1 vccd1 vccd1 _16414_/A sky130_fd_sc_hd__and2_1
X_13623_ _12705_/X _12709_/B _13627_/S vssd1 vssd1 vccd1 vccd1 _13624_/B sky130_fd_sc_hd__mux2_1
X_10835_ _10836_/A _10834_/Y _11124_/C _10933_/D vssd1 vssd1 vccd1 vccd1 _10850_/A
+ sky130_fd_sc_hd__and4bb_1
X_17391_ _17391_/A _17425_/B vssd1 vssd1 vccd1 vccd1 _17391_/X sky130_fd_sc_hd__or2_1
XFILLER_16_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16342_ _16342_/A _16342_/B vssd1 vssd1 vccd1 vccd1 _16344_/B sky130_fd_sc_hd__xnor2_1
XFILLER_13_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13554_ _13555_/A _13555_/B vssd1 vssd1 vccd1 vccd1 _13680_/B sky130_fd_sc_hd__nor2_1
X_10766_ _10764_/X _10766_/B _10766_/C vssd1 vssd1 vccd1 vccd1 _11725_/A sky130_fd_sc_hd__nand3b_2
XFILLER_160_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12505_ _17415_/A _13194_/D vssd1 vssd1 vccd1 vccd1 _12506_/B sky130_fd_sc_hd__nand2_1
X_16273_ _16273_/A _16273_/B vssd1 vssd1 vccd1 vccd1 _16276_/A sky130_fd_sc_hd__xnor2_1
X_10697_ _10694_/X _10697_/B vssd1 vssd1 vccd1 vccd1 _11036_/B sky130_fd_sc_hd__and2b_1
XFILLER_12_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13485_ _13485_/A _13485_/B vssd1 vssd1 vccd1 vccd1 _13486_/C sky130_fd_sc_hd__nand2_1
XFILLER_145_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_882 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15224_ _15222_/A _15222_/B _15225_/B vssd1 vssd1 vccd1 vccd1 _15296_/A sky130_fd_sc_hd__a21o_1
XFILLER_157_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12436_ _12437_/A _12437_/B _12437_/C vssd1 vssd1 vccd1 vccd1 _12458_/A sky130_fd_sc_hd__a21o_2
X_15155_ _15155_/A _15155_/B vssd1 vssd1 vccd1 vccd1 _15157_/B sky130_fd_sc_hd__xor2_1
X_12367_ _12198_/A _12367_/B vssd1 vssd1 vccd1 vccd1 _12368_/B sky130_fd_sc_hd__and2b_2
XFILLER_4_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14106_ _13974_/A _13974_/B _14015_/X vssd1 vssd1 vccd1 vccd1 _14108_/B sky130_fd_sc_hd__o21ai_1
X_11318_ _11423_/B _11561_/D _11317_/B _11314_/X vssd1 vssd1 vccd1 vccd1 _11320_/B
+ sky130_fd_sc_hd__a31oi_1
XFILLER_99_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12298_ _12299_/A _12299_/B vssd1 vssd1 vccd1 vccd1 _12508_/B sky130_fd_sc_hd__nor2_1
XFILLER_99_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15086_ _15726_/A _16226_/C _15085_/B vssd1 vssd1 vccd1 vccd1 _15087_/B sky130_fd_sc_hd__a21o_1
XFILLER_113_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11249_ _11249_/A _11249_/B _11249_/C vssd1 vssd1 vccd1 vccd1 _11250_/B sky130_fd_sc_hd__or3_1
XFILLER_141_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14037_ _12038_/X _14210_/B _14482_/B1 vssd1 vssd1 vccd1 vccd1 _14037_/X sky130_fd_sc_hd__o21a_1
XFILLER_79_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_900 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_302 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15988_ _15989_/A _15989_/B _15987_/X vssd1 vssd1 vccd1 vccd1 _16096_/B sky130_fd_sc_hd__o21ba_1
XFILLER_35_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14939_ _17607_/Q _17477_/D _17476_/D _17608_/Q vssd1 vssd1 vccd1 vccd1 _14939_/X
+ sky130_fd_sc_hd__and4bb_1
XFILLER_36_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_777 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16609_ _16609_/A _16609_/B _16609_/C vssd1 vssd1 vccd1 vccd1 _16610_/B sky130_fd_sc_hd__and3_1
XFILLER_23_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17589_ fanout937/X _17589_/D vssd1 vssd1 vccd1 vccd1 _17589_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_602 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09012_ _09012_/A _09012_/B _09012_/C vssd1 vssd1 vccd1 vccd1 _09013_/B sky130_fd_sc_hd__and3_1
XFILLER_128_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout602 _10792_/A vssd1 vssd1 vccd1 vccd1 _11630_/A sky130_fd_sc_hd__clkbuf_2
X_09914_ _09914_/A _09914_/B _10029_/A vssd1 vssd1 vccd1 vccd1 _09915_/B sky130_fd_sc_hd__nor3_1
Xfanout613 _11629_/B vssd1 vssd1 vccd1 vccd1 _11518_/B sky130_fd_sc_hd__buf_2
Xfanout624 _14181_/B vssd1 vssd1 vccd1 vccd1 _13844_/C sky130_fd_sc_hd__buf_2
Xfanout635 _14385_/B vssd1 vssd1 vccd1 vccd1 _14641_/C sky130_fd_sc_hd__buf_2
Xfanout646 _14765_/B vssd1 vssd1 vccd1 vccd1 _17065_/A sky130_fd_sc_hd__clkbuf_4
Xfanout657 _17505_/Q vssd1 vssd1 vccd1 vccd1 _11813_/B sky130_fd_sc_hd__buf_4
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09845_ _09845_/A _09845_/B vssd1 vssd1 vccd1 vccd1 _09847_/A sky130_fd_sc_hd__nor2_1
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout668 _14865_/B vssd1 vssd1 vccd1 vccd1 _14485_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_100_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout679 _08860_/B vssd1 vssd1 vccd1 vccd1 _14864_/A sky130_fd_sc_hd__clkbuf_4
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09776_ _09776_/A _09776_/B _09776_/C vssd1 vssd1 vccd1 vccd1 _09777_/B sky130_fd_sc_hd__and3_1
XFILLER_160_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08727_ _15008_/A vssd1 vssd1 vccd1 vccd1 _11653_/B sky130_fd_sc_hd__inv_2
XTAP_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_24 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10620_ _10963_/B _10875_/C _10962_/B _10963_/A vssd1 vssd1 vccd1 vccd1 _10621_/B
+ sky130_fd_sc_hd__a22oi_1
XFILLER_169_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10551_ _10538_/Y _10550_/X _10566_/A _10523_/Y vssd1 vssd1 vccd1 vccd1 _10566_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_128_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_115 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10482_ _10709_/A _10370_/B _10481_/X vssd1 vssd1 vccd1 vccd1 _10597_/B sky130_fd_sc_hd__o21a_1
X_13270_ _13271_/A _13271_/B vssd1 vssd1 vccd1 vccd1 _13270_/Y sky130_fd_sc_hd__nand2_1
XFILLER_108_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12221_ _11831_/Y _11835_/Y _17365_/A vssd1 vssd1 vccd1 vccd1 _12221_/X sky130_fd_sc_hd__mux2_1
XFILLER_151_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12152_ _12316_/A _12151_/B _12151_/C vssd1 vssd1 vccd1 vccd1 _12152_/X sky130_fd_sc_hd__a21o_1
XFILLER_108_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11103_ _11104_/B _11104_/C _11104_/A vssd1 vssd1 vccd1 vccd1 _11112_/B sky130_fd_sc_hd__a21o_1
XFILLER_151_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16960_ _17012_/B _16960_/B vssd1 vssd1 vccd1 vccd1 _16960_/X sky130_fd_sc_hd__xor2_1
X_12083_ _12252_/B _12083_/B vssd1 vssd1 vccd1 vccd1 _12085_/C sky130_fd_sc_hd__or2_1
XFILLER_96_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11034_ _11035_/A _11035_/B vssd1 vssd1 vccd1 vccd1 _11176_/B sky130_fd_sc_hd__and2b_1
X_15911_ _16317_/A _16054_/B vssd1 vssd1 vccd1 vccd1 _16813_/B sky130_fd_sc_hd__nand2_4
XFILLER_150_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16891_ _16807_/A _16935_/B _16808_/X _16809_/X vssd1 vssd1 vccd1 vccd1 _16893_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_103_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_806 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15842_ _15760_/A _15760_/B _15758_/X vssd1 vssd1 vccd1 vccd1 _15863_/A sky130_fd_sc_hd__o21ai_1
XFILLER_76_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15773_ _15773_/A _15773_/B vssd1 vssd1 vccd1 vccd1 _15775_/A sky130_fd_sc_hd__nor2_1
XFILLER_18_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12985_ _12985_/A _12985_/B _12985_/C vssd1 vssd1 vccd1 vccd1 _13125_/B sky130_fd_sc_hd__or3_2
XTAP_3551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17512_ fanout949/X _17512_/D vssd1 vssd1 vccd1 vccd1 _17512_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_3573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14724_ _14750_/A _14726_/C vssd1 vssd1 vccd1 vccd1 _14727_/B sky130_fd_sc_hd__and2_1
XTAP_3584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11936_ _11936_/A _11936_/B vssd1 vssd1 vccd1 vccd1 _11937_/B sky130_fd_sc_hd__nor2_1
XTAP_3595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17443_ fanout938/X _17443_/D vssd1 vssd1 vccd1 vccd1 _17443_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14655_ _14655_/A _14655_/B vssd1 vssd1 vccd1 vccd1 _14656_/B sky130_fd_sc_hd__or2_1
XTAP_2894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11867_ _12077_/A _12077_/B _12077_/D _11867_/D vssd1 vssd1 vccd1 vccd1 _12093_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_60_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13606_ _13607_/A _13607_/B _13607_/C vssd1 vssd1 vccd1 vccd1 _13718_/A sky130_fd_sc_hd__o21ai_1
X_10818_ _10823_/A _10823_/B vssd1 vssd1 vccd1 vccd1 _10829_/A sky130_fd_sc_hd__nor2_1
XFILLER_159_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17374_ input63/X _17424_/A2 _17373_/X _17388_/C1 vssd1 vssd1 vccd1 vccd1 _17515_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_158_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14586_ _14629_/C _14587_/B vssd1 vssd1 vccd1 vccd1 _14586_/X sky130_fd_sc_hd__or2_1
X_11798_ _14888_/B _11798_/B _11798_/C _11798_/D vssd1 vssd1 vccd1 vccd1 _11800_/C
+ sky130_fd_sc_hd__or4_1
XFILLER_13_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16325_ _16497_/A _16499_/B vssd1 vssd1 vccd1 vccd1 _16326_/B sky130_fd_sc_hd__nor2_1
X_13537_ _13538_/A _13538_/B vssd1 vssd1 vccd1 vccd1 _13537_/Y sky130_fd_sc_hd__nor2_1
X_10749_ _10750_/B _10750_/C _10750_/A vssd1 vssd1 vccd1 vccd1 _10760_/A sky130_fd_sc_hd__a21o_1
XFILLER_174_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16256_ _16257_/A _16257_/B vssd1 vssd1 vccd1 vccd1 _16256_/X sky130_fd_sc_hd__and2_1
X_13468_ _13977_/A _13977_/B _13866_/D _13764_/D vssd1 vssd1 vccd1 vccd1 _13469_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_127_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15207_ _15262_/C _15208_/C _15208_/D vssd1 vssd1 vccd1 vccd1 _15207_/X sky130_fd_sc_hd__or3_1
XFILLER_173_468 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12419_ _12419_/A _12419_/B vssd1 vssd1 vccd1 vccd1 _12421_/C sky130_fd_sc_hd__xnor2_1
X_16187_ _16188_/A _16188_/B _16188_/C vssd1 vssd1 vccd1 vccd1 _16187_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_142_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13399_ _13398_/C _13526_/A _13397_/Y vssd1 vssd1 vccd1 vccd1 _13401_/B sky130_fd_sc_hd__a21bo_1
XFILLER_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15138_ _16025_/A _16315_/B vssd1 vssd1 vccd1 vccd1 _15159_/A sky130_fd_sc_hd__nor2_1
XFILLER_142_844 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15069_ _16021_/A _17612_/Q vssd1 vssd1 vccd1 vccd1 _15069_/X sky130_fd_sc_hd__and2_1
XFILLER_142_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_931 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09630_ _09630_/A _09630_/B vssd1 vssd1 vccd1 vccd1 _09632_/B sky130_fd_sc_hd__xnor2_1
XFILLER_67_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09561_ _09574_/B _09574_/C _09574_/A vssd1 vssd1 vccd1 vccd1 _09576_/A sky130_fd_sc_hd__o21ai_1
XFILLER_83_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09492_ _11839_/S _11808_/B vssd1 vssd1 vccd1 vccd1 _14949_/A sky130_fd_sc_hd__and2_1
XFILLER_24_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_104 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_997 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout410 _17530_/Q vssd1 vssd1 vccd1 vccd1 _12068_/A sky130_fd_sc_hd__buf_4
Xfanout421 _13632_/B vssd1 vssd1 vccd1 vccd1 _13735_/B sky130_fd_sc_hd__buf_2
Xfanout432 _14777_/A vssd1 vssd1 vccd1 vccd1 _12722_/A sky130_fd_sc_hd__buf_2
Xfanout443 _12077_/B vssd1 vssd1 vccd1 vccd1 _17395_/A sky130_fd_sc_hd__clkbuf_4
Xfanout454 _09412_/A vssd1 vssd1 vccd1 vccd1 _17393_/A sky130_fd_sc_hd__buf_6
XFILLER_87_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout465 _17523_/Q vssd1 vssd1 vccd1 vccd1 _13414_/B sky130_fd_sc_hd__buf_2
XFILLER_24_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout476 _15393_/A vssd1 vssd1 vccd1 vccd1 _16136_/A sky130_fd_sc_hd__clkbuf_4
X_09828_ _09828_/A _09828_/B vssd1 vssd1 vccd1 vccd1 _09966_/A sky130_fd_sc_hd__xor2_2
Xfanout487 _15262_/A vssd1 vssd1 vccd1 vccd1 _10142_/A sky130_fd_sc_hd__clkbuf_4
Xfanout498 _09730_/C vssd1 vssd1 vccd1 vccd1 _17381_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_100_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_699 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09759_ _09890_/A _09898_/A _09890_/C vssd1 vssd1 vccd1 vccd1 _09891_/A sky130_fd_sc_hd__o21ai_2
XTAP_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_850 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12770_ _12770_/A _12770_/B _12923_/D _12770_/D vssd1 vssd1 vccd1 vccd1 _12771_/B
+ sky130_fd_sc_hd__and4_1
XTAP_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11721_ _10774_/A _10774_/C _10774_/B vssd1 vssd1 vccd1 vccd1 _11722_/B sky130_fd_sc_hd__o21a_1
XFILLER_15_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_566 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14440_ _14440_/A _14440_/B _14440_/C vssd1 vssd1 vccd1 vccd1 _14441_/B sky130_fd_sc_hd__nor3_1
X_11652_ _14796_/A _11675_/C vssd1 vssd1 vccd1 vccd1 _11657_/B sky130_fd_sc_hd__nor2_1
XFILLER_120_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_728 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_763 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10603_ _10603_/A _10603_/B vssd1 vssd1 vccd1 vccd1 _10610_/A sky130_fd_sc_hd__xor2_2
XFILLER_11_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14371_ _14372_/A _14372_/B _14372_/C vssd1 vssd1 vccd1 vccd1 _14445_/A sky130_fd_sc_hd__o21ai_1
X_11583_ _11583_/A _11583_/B vssd1 vssd1 vccd1 vccd1 _11583_/Y sky130_fd_sc_hd__nand2_1
XFILLER_11_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_616 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16110_ _16107_/Y _16108_/X _16001_/A _16003_/X vssd1 vssd1 vccd1 vccd1 _16111_/C
+ sky130_fd_sc_hd__o211a_1
X_13322_ _13322_/A _13322_/B vssd1 vssd1 vccd1 vccd1 _13324_/A sky130_fd_sc_hd__nor2_1
X_10534_ _10535_/A _10533_/Y _10745_/C _10534_/D vssd1 vssd1 vccd1 vccd1 _10644_/A
+ sky130_fd_sc_hd__and4bb_1
X_17090_ _17090_/A _17093_/B vssd1 vssd1 vccd1 vccd1 _17118_/B sky130_fd_sc_hd__nor2_1
XFILLER_10_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16041_ _16667_/A _16041_/B _16041_/C vssd1 vssd1 vccd1 vccd1 _16043_/A sky130_fd_sc_hd__or3_1
X_13253_ _13249_/Y _13250_/X _13121_/A _13123_/A vssd1 vssd1 vccd1 vccd1 _13253_/Y
+ sky130_fd_sc_hd__a211oi_1
X_10465_ _10465_/A _10465_/B vssd1 vssd1 vccd1 vccd1 _10469_/C sky130_fd_sc_hd__xnor2_1
XFILLER_124_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12204_ _12371_/A _12202_/Y _11967_/A _11971_/A vssd1 vssd1 vccd1 vccd1 _12206_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_163_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10396_ _10397_/B _10397_/A vssd1 vssd1 vccd1 vccd1 _10396_/X sky130_fd_sc_hd__and2b_1
X_13184_ _13184_/A _13184_/B vssd1 vssd1 vccd1 vccd1 _13186_/B sky130_fd_sc_hd__xnor2_1
XFILLER_89_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12135_ _12471_/A _14925_/A _12592_/C _12592_/D vssd1 vssd1 vccd1 vccd1 _12136_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_2_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16943_ _16943_/A _16943_/B vssd1 vssd1 vccd1 vccd1 _16944_/B sky130_fd_sc_hd__or2_1
XFILLER_49_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12066_ _15998_/A _12018_/Y _12065_/X vssd1 vssd1 vccd1 vccd1 _17577_/D sky130_fd_sc_hd__o21ai_1
XFILLER_1_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11017_ _11117_/C _10933_/D _10739_/A _10737_/Y vssd1 vssd1 vccd1 vccd1 _11018_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_78_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16874_ _16485_/A _16865_/Y _16873_/X vssd1 vssd1 vccd1 vccd1 _16874_/X sky130_fd_sc_hd__a21o_1
XFILLER_65_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15825_ _15825_/A _15825_/B vssd1 vssd1 vccd1 vccd1 _15827_/B sky130_fd_sc_hd__xnor2_1
XFILLER_37_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15756_ _15756_/A _15756_/B vssd1 vssd1 vccd1 vccd1 _15759_/A sky130_fd_sc_hd__xnor2_1
X_12968_ _12968_/A _12968_/B vssd1 vssd1 vccd1 vccd1 _12971_/A sky130_fd_sc_hd__xnor2_1
XFILLER_18_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14707_ _14708_/B _14738_/B _14708_/D _14738_/A vssd1 vssd1 vccd1 vccd1 _14713_/A
+ sky130_fd_sc_hd__a22o_1
X_11919_ _17423_/A _12127_/D _11920_/D _17425_/A vssd1 vssd1 vccd1 vccd1 _11921_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_45_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15687_ _15687_/A _16747_/A _15686_/Y vssd1 vssd1 vccd1 vccd1 _15782_/B sky130_fd_sc_hd__or3b_1
X_12899_ _13049_/A _12899_/B _12899_/C vssd1 vssd1 vccd1 vccd1 _13049_/B sky130_fd_sc_hd__nand3_1
XTAP_2691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1047 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17426_ input60/X _17426_/A2 _17425_/X _17426_/C1 vssd1 vssd1 vccd1 vccd1 _17541_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_60_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14638_ _14638_/A _14638_/B vssd1 vssd1 vccd1 vccd1 _14664_/A sky130_fd_sc_hd__nand2_1
XFILLER_20_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17357_ input59/X _17359_/B _17359_/C vssd1 vssd1 vccd1 vccd1 _17357_/X sky130_fd_sc_hd__or3_1
X_14569_ _14569_/A _14569_/B _14569_/C vssd1 vssd1 vccd1 vccd1 _14570_/C sky130_fd_sc_hd__nand3_1
XFILLER_159_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_250 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16308_ _16302_/A _17163_/A2 _16307_/X vssd1 vssd1 vccd1 vccd1 _16310_/C sky130_fd_sc_hd__o21ba_1
X_17288_ _17605_/Q _17291_/A2 _17291_/B1 vssd1 vssd1 vccd1 vccd1 _17288_/X sky130_fd_sc_hd__a21o_1
XFILLER_118_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16239_ _16239_/A _16239_/B vssd1 vssd1 vccd1 vccd1 _16239_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_173_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08992_ _08994_/A vssd1 vssd1 vccd1 vccd1 _08992_/Y sky130_fd_sc_hd__inv_2
XFILLER_87_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_836 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09613_ _09746_/A _09612_/Y _15538_/A _10180_/B vssd1 vssd1 vccd1 vccd1 _09754_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_141_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09544_ _09436_/A _09435_/C _09435_/B vssd1 vssd1 vccd1 vccd1 _09577_/B sky130_fd_sc_hd__a21o_1
XFILLER_24_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09475_ _09602_/A _09610_/A _09602_/C vssd1 vssd1 vccd1 vccd1 _09603_/A sky130_fd_sc_hd__o21ai_2
XFILLER_63_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_527 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_903 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xwire118 wire118/A vssd1 vssd1 vccd1 vccd1 wire118/X sky130_fd_sc_hd__clkbuf_1
XFILLER_149_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10250_ _10243_/B _10245_/B _10243_/A vssd1 vssd1 vccd1 vccd1 _10253_/A sky130_fd_sc_hd__o21ba_1
XFILLER_105_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10181_ _15254_/S _10431_/B _14952_/A vssd1 vssd1 vccd1 vccd1 _10181_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_133_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout240 _16401_/C1 vssd1 vssd1 vccd1 vccd1 _16494_/B1 sky130_fd_sc_hd__clkbuf_4
Xfanout251 _15108_/A vssd1 vssd1 vccd1 vccd1 _16485_/A sky130_fd_sc_hd__buf_4
XFILLER_59_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout262 _17359_/C vssd1 vssd1 vccd1 vccd1 _17355_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_47_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13940_ _14122_/A wire116/X vssd1 vssd1 vccd1 vccd1 _13940_/X sky130_fd_sc_hd__and2_1
Xfanout273 _15373_/B vssd1 vssd1 vccd1 vccd1 _16644_/B sky130_fd_sc_hd__buf_2
XFILLER_19_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout284 _15275_/C1 vssd1 vssd1 vccd1 vccd1 _17363_/A sky130_fd_sc_hd__buf_2
Xfanout295 fanout299/X vssd1 vssd1 vccd1 vccd1 _15384_/S sky130_fd_sc_hd__clkbuf_4
X_13871_ _13768_/A _13768_/B _13762_/A vssd1 vssd1 vccd1 vccd1 _13873_/B sky130_fd_sc_hd__a21o_1
XFILLER_35_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_77 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15610_ _15610_/A _15610_/B vssd1 vssd1 vccd1 vccd1 _15610_/Y sky130_fd_sc_hd__nor2_1
X_12822_ _12823_/B _12822_/B vssd1 vssd1 vccd1 vccd1 _12824_/A sky130_fd_sc_hd__nand2b_1
XFILLER_62_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16590_ _16590_/A _16686_/A vssd1 vssd1 vccd1 vccd1 _16591_/C sky130_fd_sc_hd__nor2_1
XFILLER_90_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15541_ _15541_/A _15541_/B vssd1 vssd1 vccd1 vccd1 _15541_/Y sky130_fd_sc_hd__nor2_1
X_12753_ _12907_/A _13051_/D _12754_/A vssd1 vssd1 vccd1 vccd1 _12910_/B sky130_fd_sc_hd__and3_1
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_875 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11704_ _11705_/A _11704_/B vssd1 vssd1 vccd1 vccd1 _15889_/A sky130_fd_sc_hd__xnor2_2
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15472_ _15472_/A _15472_/B vssd1 vssd1 vccd1 vccd1 _15472_/Y sky130_fd_sc_hd__nand2_1
XFILLER_43_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12684_ _12685_/A _12685_/B vssd1 vssd1 vccd1 vccd1 _12684_/X sky130_fd_sc_hd__or2_1
XFILLER_30_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17211_ _17547_/Q _17274_/B vssd1 vssd1 vccd1 vccd1 _17211_/X sky130_fd_sc_hd__and2_1
X_14423_ _14734_/A _14421_/X _14422_/X vssd1 vssd1 vccd1 vccd1 _14423_/Y sky130_fd_sc_hd__a21oi_2
X_11635_ _11635_/A _11635_/B vssd1 vssd1 vccd1 vccd1 _11659_/A sky130_fd_sc_hd__xnor2_1
XFILLER_156_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17142_ _17167_/A _17163_/A2 _17141_/X vssd1 vssd1 vccd1 vccd1 _17142_/X sky130_fd_sc_hd__o21ba_1
XFILLER_168_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14354_ _14416_/B _14354_/B vssd1 vssd1 vccd1 vccd1 _14354_/X sky130_fd_sc_hd__or2_1
XFILLER_155_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11566_ _11566_/A _11566_/B vssd1 vssd1 vccd1 vccd1 _11568_/B sky130_fd_sc_hd__xnor2_1
XFILLER_156_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13305_ _13306_/A _13306_/B vssd1 vssd1 vccd1 vccd1 _13305_/Y sky130_fd_sc_hd__nand2b_1
X_10517_ _10517_/A _10517_/B vssd1 vssd1 vccd1 vccd1 _10519_/B sky130_fd_sc_hd__nand2_1
X_17073_ _17065_/A _17029_/B _17072_/Y vssd1 vssd1 vccd1 vccd1 _17077_/B sky130_fd_sc_hd__o21a_1
XFILLER_143_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14285_ _17070_/B _14283_/X _14352_/B _14211_/X vssd1 vssd1 vccd1 vccd1 _17595_/D
+ sky130_fd_sc_hd__o31ai_1
X_11497_ _11502_/A _11497_/B vssd1 vssd1 vccd1 vccd1 _11499_/B sky130_fd_sc_hd__nand2_1
XFILLER_157_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_298 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16024_ _15913_/A _16023_/Y _16022_/X vssd1 vssd1 vccd1 vccd1 _16026_/A sky130_fd_sc_hd__o21ai_1
XFILLER_143_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13236_ _13236_/A _13236_/B vssd1 vssd1 vccd1 vccd1 _13238_/B sky130_fd_sc_hd__nor2_1
XFILLER_6_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10448_ _10685_/A _10448_/B vssd1 vssd1 vccd1 vccd1 _10563_/B sky130_fd_sc_hd__nor2_1
XFILLER_152_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13167_ _13027_/A _13029_/B _13027_/B vssd1 vssd1 vccd1 vccd1 _13174_/A sky130_fd_sc_hd__o21ba_1
X_10379_ _10379_/A _10379_/B vssd1 vssd1 vccd1 vccd1 _10487_/B sky130_fd_sc_hd__nor2_1
XFILLER_112_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12118_ _12118_/A _12118_/B _12118_/C vssd1 vssd1 vccd1 vccd1 _12118_/Y sky130_fd_sc_hd__nand3_1
XFILLER_69_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13098_ _13227_/A _14153_/B _13551_/D _13434_/D vssd1 vssd1 vccd1 vccd1 _13099_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_97_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16926_ _14080_/C _17075_/A2 _16925_/X vssd1 vssd1 vccd1 vccd1 _16926_/Y sky130_fd_sc_hd__a21oi_1
X_12049_ _14911_/B _12049_/B vssd1 vssd1 vccd1 vccd1 _12049_/Y sky130_fd_sc_hd__nand2_1
XFILLER_37_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16857_ _16931_/A _16931_/B _16856_/Y vssd1 vssd1 vccd1 vccd1 _16857_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_26_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15808_ _15808_/A _15808_/B vssd1 vssd1 vccd1 vccd1 _15808_/Y sky130_fd_sc_hd__nor2_1
X_16788_ _13689_/A _17134_/C _16789_/A vssd1 vssd1 vccd1 vccd1 _16788_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_81_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15739_ _15740_/A _15740_/B vssd1 vssd1 vccd1 vccd1 _15861_/A sky130_fd_sc_hd__and2b_1
XFILLER_34_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09260_ _09050_/A _09049_/C _09049_/B vssd1 vssd1 vccd1 vccd1 _09261_/B sky130_fd_sc_hd__a21o_1
XFILLER_61_683 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17409_ _17409_/A _17421_/B vssd1 vssd1 vccd1 vccd1 _17409_/X sky130_fd_sc_hd__or2_1
X_09191_ _09942_/A _09514_/B _12174_/D _12129_/B vssd1 vssd1 vccd1 vccd1 _09196_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_14_1003 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08975_ _17423_/A _09362_/D _09172_/B _12770_/A vssd1 vssd1 vccd1 vccd1 _08977_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_152_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_880 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09527_ _09487_/X _09488_/Y _09507_/Y _09525_/X vssd1 vssd1 vccd1 vccd1 _09530_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_71_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09458_ _09483_/B _09483_/A vssd1 vssd1 vccd1 vccd1 _09458_/X sky130_fd_sc_hd__and2b_1
XPHY_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09389_ _09387_/A _09388_/Y _09343_/X _09344_/Y vssd1 vssd1 vccd1 vccd1 _09393_/B
+ sky130_fd_sc_hd__a211oi_4
XFILLER_61_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_711 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11420_ _11408_/A _11408_/C _11408_/B vssd1 vssd1 vccd1 vccd1 _11458_/B sky130_fd_sc_hd__o21ai_1
XFILLER_138_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11351_ _11351_/A _11402_/A _11351_/C vssd1 vssd1 vccd1 vccd1 _11354_/A sky130_fd_sc_hd__and3_1
XFILLER_4_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10302_ _10411_/A _10411_/B vssd1 vssd1 vccd1 vccd1 _10305_/C sky130_fd_sc_hd__nand2_1
XFILLER_125_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14070_ _14071_/B _14071_/A vssd1 vssd1 vccd1 vccd1 _14162_/B sky130_fd_sc_hd__and2b_1
XFILLER_153_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11282_ _11283_/B _11333_/A _11283_/A vssd1 vssd1 vccd1 vccd1 _11352_/A sky130_fd_sc_hd__o21ai_1
XFILLER_4_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13021_ _13021_/A _13021_/B vssd1 vssd1 vccd1 vccd1 _13024_/A sky130_fd_sc_hd__xnor2_1
XFILLER_10_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10233_ _10111_/C _10111_/D _10112_/A _10110_/Y vssd1 vssd1 vccd1 vccd1 _10234_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_105_151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10164_ _14786_/A _14787_/A _10647_/D _10745_/D vssd1 vssd1 vccd1 vccd1 _10167_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_120_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14972_ _14875_/X _14971_/X _15147_/D vssd1 vssd1 vccd1 vccd1 _14972_/X sky130_fd_sc_hd__a21o_1
X_10095_ _10097_/A _10097_/B vssd1 vssd1 vccd1 vccd1 _10098_/A sky130_fd_sc_hd__or2_1
XFILLER_120_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16711_ _16711_/A _16711_/B _16711_/C vssd1 vssd1 vccd1 vccd1 _16712_/B sky130_fd_sc_hd__or3_1
X_13923_ _13923_/A _13923_/B vssd1 vssd1 vccd1 vccd1 _13925_/C sky130_fd_sc_hd__xor2_1
XFILLER_47_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16642_ _16644_/C _16965_/B _16651_/A vssd1 vssd1 vccd1 vccd1 _16643_/A sky130_fd_sc_hd__a21boi_2
X_13854_ _13748_/A _13748_/B _13742_/A vssd1 vssd1 vccd1 vccd1 _13856_/B sky130_fd_sc_hd__a21o_1
XFILLER_90_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12805_ _12805_/A _12805_/B vssd1 vssd1 vccd1 vccd1 _12807_/A sky130_fd_sc_hd__nor2_1
X_16573_ _16481_/A _16482_/Y _16572_/Y vssd1 vssd1 vccd1 vccd1 _16574_/B sky130_fd_sc_hd__a21o_1
XFILLER_27_190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13785_ _13891_/A _13785_/B vssd1 vssd1 vccd1 vccd1 _13787_/B sky130_fd_sc_hd__nor2_1
X_10997_ _11164_/B _10996_/B _10996_/C vssd1 vssd1 vccd1 vccd1 _10998_/B sky130_fd_sc_hd__o21ai_1
XFILLER_43_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_970 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15524_ _11624_/Y _15524_/B _15524_/C vssd1 vssd1 vccd1 vccd1 _15525_/B sky130_fd_sc_hd__nand3b_1
XFILLER_163_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12736_ _13302_/A _17505_/Q vssd1 vssd1 vccd1 vccd1 _12737_/B sky130_fd_sc_hd__nand2_1
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15455_ _14805_/A _14805_/B _14805_/C vssd1 vssd1 vccd1 vccd1 _15455_/X sky130_fd_sc_hd__a21o_1
X_12667_ _12668_/A _12668_/B vssd1 vssd1 vccd1 vccd1 _12816_/A sky130_fd_sc_hd__or2_1
X_14406_ _14405_/B _14405_/C _14405_/A vssd1 vssd1 vccd1 vccd1 _14406_/Y sky130_fd_sc_hd__a21oi_1
X_11618_ _11617_/B _11616_/Y _11583_/B _11587_/X vssd1 vssd1 vccd1 vccd1 _11624_/A
+ sky130_fd_sc_hd__o211ai_2
X_15386_ _15386_/A _15386_/B vssd1 vssd1 vccd1 vccd1 _15386_/Y sky130_fd_sc_hd__nand2_1
X_12598_ _12599_/A _12599_/B vssd1 vssd1 vccd1 vccd1 _12600_/A sky130_fd_sc_hd__nor2_1
XFILLER_128_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17125_ _17125_/A _17125_/B vssd1 vssd1 vccd1 vccd1 _17127_/B sky130_fd_sc_hd__nand2_1
X_14337_ _14337_/A _14405_/A _14337_/C vssd1 vssd1 vccd1 vccd1 _14337_/Y sky130_fd_sc_hd__nor3_1
X_11549_ _15888_/A _11549_/B vssd1 vssd1 vccd1 vccd1 _15793_/A sky130_fd_sc_hd__and2_1
XFILLER_144_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17056_ _17057_/B _17056_/B vssd1 vssd1 vccd1 vccd1 _17096_/A sky130_fd_sc_hd__and2b_1
XFILLER_171_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14268_ _14268_/A _14268_/B vssd1 vssd1 vccd1 vccd1 _14270_/C sky130_fd_sc_hd__xnor2_1
XFILLER_143_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16007_ _16007_/A _16007_/B _16007_/C vssd1 vssd1 vccd1 vccd1 _16007_/X sky130_fd_sc_hd__or3_1
X_13219_ _13220_/A _13220_/B _13220_/C vssd1 vssd1 vccd1 vccd1 _13221_/A sky130_fd_sc_hd__a21o_1
XFILLER_125_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14199_ _14200_/A _14200_/B _14198_/X vssd1 vssd1 vccd1 vccd1 _14276_/B sky130_fd_sc_hd__o21ba_1
XFILLER_140_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_912 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08760_ _12077_/B _13080_/D vssd1 vssd1 vccd1 vccd1 _08760_/Y sky130_fd_sc_hd__nand2_4
XFILLER_85_528 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16909_ _16909_/A _16909_/B vssd1 vssd1 vccd1 vccd1 _16910_/B sky130_fd_sc_hd__xnor2_1
XFILLER_93_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09312_ _09261_/A _09261_/B _09310_/B _09401_/A vssd1 vssd1 vccd1 vccd1 _09338_/B
+ sky130_fd_sc_hd__a31oi_2
XFILLER_62_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09243_ _11990_/A _09243_/B vssd1 vssd1 vccd1 vccd1 _09245_/C sky130_fd_sc_hd__nand2_1
XFILLER_90_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_366 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09174_ _09172_/A _09362_/D _09172_/B _09360_/A vssd1 vssd1 vccd1 vccd1 _09174_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_147_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08958_ _08958_/A _09084_/A vssd1 vssd1 vccd1 vccd1 _09077_/A sky130_fd_sc_hd__or2_1
XFILLER_103_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08889_ _08889_/A _08889_/B vssd1 vssd1 vccd1 vccd1 _09020_/B sky130_fd_sc_hd__xnor2_1
XFILLER_45_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10920_ _14786_/A _10920_/B vssd1 vssd1 vccd1 vccd1 _14806_/A sky130_fd_sc_hd__and2_2
XFILLER_45_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10851_ _10933_/A _10851_/B _15541_/A _14895_/B vssd1 vssd1 vccd1 vccd1 _10854_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_60_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_683 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13570_ _13569_/A _13569_/B _13569_/C vssd1 vssd1 vccd1 vccd1 _13702_/A sky130_fd_sc_hd__o21ai_1
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10782_ _10685_/B _10688_/A _10579_/B _10584_/X vssd1 vssd1 vccd1 vccd1 _11768_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_158_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12521_ _12521_/A _12521_/B vssd1 vssd1 vccd1 vccd1 _12522_/C sky130_fd_sc_hd__xor2_1
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15240_ _15241_/A _15241_/B _15241_/C vssd1 vssd1 vccd1 vccd1 _15242_/B sky130_fd_sc_hd__a21o_1
X_12452_ _12452_/A _12452_/B vssd1 vssd1 vccd1 vccd1 _12454_/C sky130_fd_sc_hd__xnor2_1
XFILLER_8_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11403_ _11403_/A _11403_/B vssd1 vssd1 vccd1 vccd1 _11406_/B sky130_fd_sc_hd__and2_1
X_15171_ _15171_/A _15171_/B vssd1 vssd1 vccd1 vccd1 _15171_/Y sky130_fd_sc_hd__xnor2_1
X_12383_ _12046_/Y _12049_/Y _12383_/S vssd1 vssd1 vccd1 vccd1 _12383_/X sky130_fd_sc_hd__mux2_1
XFILLER_165_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14122_ _14122_/A _14122_/B vssd1 vssd1 vccd1 vccd1 _14281_/A sky130_fd_sc_hd__nor2_1
X_11334_ _11561_/A _11518_/B _15617_/A _14851_/A vssd1 vssd1 vccd1 vccd1 _11337_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_126_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_972 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14053_ _14054_/A _14054_/B vssd1 vssd1 vccd1 vccd1 _14158_/B sky130_fd_sc_hd__nor2_1
X_11265_ _11506_/A _11561_/C vssd1 vssd1 vccd1 vccd1 _15244_/A sky130_fd_sc_hd__and2_2
X_13004_ _13004_/A _13004_/B vssd1 vssd1 vccd1 vccd1 _13005_/B sky130_fd_sc_hd__nor2_1
XFILLER_79_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10216_ _10216_/A _10216_/B _10216_/C vssd1 vssd1 vccd1 vccd1 _10219_/A sky130_fd_sc_hd__and3_1
X_11196_ _11088_/A _11087_/B _11087_/A vssd1 vssd1 vccd1 vccd1 _11198_/B sky130_fd_sc_hd__o21ba_1
XFILLER_122_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10147_ _10148_/B _10148_/C _10148_/A vssd1 vssd1 vccd1 vccd1 _10149_/A sky130_fd_sc_hd__o21a_1
XFILLER_94_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14955_ _14954_/A _14952_/Y _14954_/Y _14912_/Y vssd1 vssd1 vccd1 vccd1 _14955_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_36_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10078_ _10078_/A _10078_/B vssd1 vssd1 vccd1 vccd1 _10080_/B sky130_fd_sc_hd__xor2_1
XFILLER_75_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13906_ _13906_/A _13906_/B _13906_/C vssd1 vssd1 vccd1 vccd1 _13907_/B sky130_fd_sc_hd__and3_1
X_14886_ _15373_/C _15305_/C _14924_/A _14886_/D vssd1 vssd1 vccd1 vccd1 _14886_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_62_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16625_ _16625_/A _16625_/B _16623_/X vssd1 vssd1 vccd1 vccd1 _16626_/B sky130_fd_sc_hd__or3b_1
X_13837_ _17164_/A _17164_/B _13837_/C vssd1 vssd1 vccd1 vccd1 _14841_/B sky130_fd_sc_hd__or3_1
XFILLER_23_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16556_ _16638_/A vssd1 vssd1 vccd1 vccd1 _16558_/B sky130_fd_sc_hd__inv_2
X_13768_ _13768_/A _13768_/B vssd1 vssd1 vccd1 vccd1 _13770_/C sky130_fd_sc_hd__xor2_1
XFILLER_43_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12719_ _12720_/A _12720_/B vssd1 vssd1 vccd1 vccd1 _12886_/A sky130_fd_sc_hd__and2_1
X_15507_ _15507_/A _15507_/B vssd1 vssd1 vccd1 vccd1 _15510_/A sky130_fd_sc_hd__xnor2_1
X_16487_ _16480_/A _16400_/B _16579_/A vssd1 vssd1 vccd1 vccd1 _16487_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_30_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13699_ _14176_/A _16859_/A _13698_/C vssd1 vssd1 vccd1 vccd1 _13700_/B sky130_fd_sc_hd__a21o_1
XFILLER_87_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15438_ _15439_/A _15439_/B vssd1 vssd1 vccd1 vccd1 _15520_/B sky130_fd_sc_hd__and2b_1
XFILLER_30_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15369_ _15369_/A _15369_/B vssd1 vssd1 vccd1 vccd1 _15369_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_8_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17108_ _17065_/A _17029_/B _14867_/A vssd1 vssd1 vccd1 vccd1 _17109_/C sky130_fd_sc_hd__a21oi_1
XFILLER_132_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17039_ _17038_/C _17040_/B _17040_/A vssd1 vssd1 vccd1 vccd1 _17039_/X sky130_fd_sc_hd__o21a_1
X_09930_ _09930_/A _09930_/B _09930_/C vssd1 vssd1 vccd1 vccd1 _10074_/B sky130_fd_sc_hd__or3_1
XFILLER_171_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout806 _12158_/D vssd1 vssd1 vccd1 vccd1 _13067_/D sky130_fd_sc_hd__clkbuf_4
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout817 _09265_/C vssd1 vssd1 vccd1 vccd1 _12338_/C sky130_fd_sc_hd__buf_4
X_09861_ _09862_/B _09862_/A vssd1 vssd1 vccd1 vccd1 _09870_/B sky130_fd_sc_hd__nand2b_1
XFILLER_113_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout828 _17486_/Q vssd1 vssd1 vccd1 vccd1 _12770_/D sky130_fd_sc_hd__buf_4
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout839 _11387_/B vssd1 vssd1 vccd1 vccd1 _14850_/A sky130_fd_sc_hd__clkbuf_4
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08812_ _08812_/A _08812_/B vssd1 vssd1 vccd1 vccd1 _08814_/A sky130_fd_sc_hd__nor2_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09792_ _10560_/A _09937_/B _09643_/C vssd1 vssd1 vccd1 vccd1 _09793_/B sky130_fd_sc_hd__a21oi_1
XFILLER_100_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08743_ _08743_/A _14872_/A vssd1 vssd1 vccd1 vccd1 _08743_/Y sky130_fd_sc_hd__nor2_1
XFILLER_54_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_49 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_255 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_586 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09226_ _09227_/A _09227_/B _09227_/C vssd1 vssd1 vccd1 vccd1 _09228_/A sky130_fd_sc_hd__a21oi_1
XFILLER_139_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09157_ _09654_/C _11815_/B _09101_/A _09099_/Y vssd1 vssd1 vccd1 vccd1 _09165_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_147_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09088_ _09088_/A _09088_/B vssd1 vssd1 vccd1 vccd1 _09317_/C sky130_fd_sc_hd__xnor2_1
XFILLER_135_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_780 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_30 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11050_ _11051_/A _11051_/B _11051_/C vssd1 vssd1 vccd1 vccd1 _11050_/X sky130_fd_sc_hd__and3_1
XFILLER_153_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10001_ _10123_/A _10000_/B _10000_/A vssd1 vssd1 vccd1 vccd1 _10003_/B sky130_fd_sc_hd__o21ba_1
XFILLER_131_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14740_ _17151_/A _14739_/Y _14737_/X vssd1 vssd1 vccd1 vccd1 _14742_/B sky130_fd_sc_hd__o21a_1
X_11952_ _17411_/A _12158_/D _12923_/D _17413_/A vssd1 vssd1 vccd1 vccd1 _11956_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_57_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_22 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10903_ _11005_/A _17466_/D vssd1 vssd1 vccd1 vccd1 _11347_/A sky130_fd_sc_hd__nand2_1
XFILLER_72_553 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14671_ _14660_/B _14662_/A _14670_/X vssd1 vssd1 vccd1 vccd1 _14671_/X sky130_fd_sc_hd__a21o_1
X_11883_ _17387_/A _12256_/D vssd1 vssd1 vccd1 vccd1 _11884_/B sky130_fd_sc_hd__nand2_1
X_16410_ _16410_/A _16595_/B _16504_/B vssd1 vssd1 vccd1 vccd1 _16505_/B sky130_fd_sc_hd__or3_1
XFILLER_72_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13622_ _14756_/A1 _13620_/Y _13621_/X _13517_/Y _13520_/X vssd1 vssd1 vccd1 vccd1
+ _17588_/D sky130_fd_sc_hd__a32o_1
X_10834_ _11122_/B _10970_/B _10971_/B _10933_/A vssd1 vssd1 vccd1 vccd1 _10834_/Y
+ sky130_fd_sc_hd__a22oi_1
X_17390_ input40/X _17426_/A2 _17389_/X _17426_/C1 vssd1 vssd1 vccd1 vccd1 _17523_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_32_439 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16341_ _16342_/A _16342_/B vssd1 vssd1 vccd1 vccd1 _16444_/B sky130_fd_sc_hd__and2b_1
XFILLER_41_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13553_ _14215_/A _13764_/D vssd1 vssd1 vccd1 vccd1 _13555_/B sky130_fd_sc_hd__nand2_1
X_10765_ _10631_/X _10693_/Y _10712_/X _10730_/Y vssd1 vssd1 vccd1 vccd1 _10766_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_34_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12504_ _12504_/A _12504_/B vssd1 vssd1 vccd1 vccd1 _12506_/A sky130_fd_sc_hd__nor2_1
X_16272_ _16272_/A _16272_/B vssd1 vssd1 vccd1 vccd1 _16273_/B sky130_fd_sc_hd__xnor2_1
XFILLER_157_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13484_ _13485_/A _13485_/B vssd1 vssd1 vccd1 vccd1 _13603_/B sky130_fd_sc_hd__or2_1
X_10696_ _11027_/A _11027_/C _10905_/D _10694_/A vssd1 vssd1 vccd1 vccd1 _10697_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_139_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_494 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15223_ _16086_/A _15647_/A vssd1 vssd1 vccd1 vccd1 _15225_/B sky130_fd_sc_hd__nand2_1
X_12435_ _12435_/A _12588_/B vssd1 vssd1 vccd1 vccd1 _12437_/C sky130_fd_sc_hd__nand2_1
XFILLER_8_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15154_ _15155_/A _15155_/B vssd1 vssd1 vccd1 vccd1 _15222_/A sky130_fd_sc_hd__or2_1
XFILLER_5_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12366_ _12366_/A _12366_/B vssd1 vssd1 vccd1 vccd1 _12368_/A sky130_fd_sc_hd__or2_1
XFILLER_114_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14105_ _14192_/B _14105_/B vssd1 vssd1 vccd1 vccd1 _14108_/A sky130_fd_sc_hd__nand2_1
X_11317_ _11314_/X _11317_/B vssd1 vssd1 vccd1 vccd1 _11362_/B sky130_fd_sc_hd__and2b_1
XFILLER_154_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15085_ _15913_/A _15085_/B vssd1 vssd1 vccd1 vccd1 _15161_/A sky130_fd_sc_hd__nand2b_1
X_12297_ _17421_/A _12618_/D vssd1 vssd1 vccd1 vccd1 _12299_/B sky130_fd_sc_hd__nand2_1
XFILLER_4_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14036_ _12057_/X _12063_/X _16012_/S vssd1 vssd1 vccd1 vccd1 _14036_/X sky130_fd_sc_hd__mux2_1
X_11248_ _11249_/B _11249_/C _11249_/A vssd1 vssd1 vccd1 vccd1 _11255_/B sky130_fd_sc_hd__o21ai_1
XFILLER_80_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_912 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11179_ _11175_/Y _11176_/X _11015_/X _11019_/X vssd1 vssd1 vccd1 vccd1 _11182_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_94_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15987_ _15987_/A _15987_/B vssd1 vssd1 vccd1 vccd1 _15987_/X sky130_fd_sc_hd__xor2_1
XFILLER_36_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14938_ _17607_/Q _14938_/B vssd1 vssd1 vccd1 vccd1 _14938_/X sky130_fd_sc_hd__or2_1
XFILLER_36_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14869_ _08967_/B _15248_/C _17140_/B _14838_/X _14842_/X vssd1 vssd1 vccd1 vccd1
+ _14869_/X sky130_fd_sc_hd__a311o_1
XFILLER_23_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16608_ _16609_/A _16609_/B _16609_/C vssd1 vssd1 vccd1 vccd1 _16697_/A sky130_fd_sc_hd__a21oi_1
XFILLER_35_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17588_ fanout935/X _17588_/D vssd1 vssd1 vccd1 vccd1 _17588_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16539_ _16541_/A _16541_/B vssd1 vssd1 vccd1 vccd1 _16627_/A sky130_fd_sc_hd__nand2_1
XFILLER_31_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_472 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09011_ _09012_/A _09012_/B _09012_/C vssd1 vssd1 vccd1 vccd1 _09013_/A sky130_fd_sc_hd__a21oi_1
XFILLER_12_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_227 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09913_ _09913_/A _09913_/B vssd1 vssd1 vccd1 vccd1 _09973_/A sky130_fd_sc_hd__nand2_1
XFILLER_99_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout603 _14982_/A vssd1 vssd1 vccd1 vccd1 _10792_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_113_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout614 _11132_/B vssd1 vssd1 vccd1 vccd1 _11629_/B sky130_fd_sc_hd__clkbuf_2
Xfanout625 _13051_/D vssd1 vssd1 vccd1 vccd1 _14181_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_98_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout636 _14867_/A vssd1 vssd1 vccd1 vccd1 _14385_/B sky130_fd_sc_hd__buf_2
XFILLER_59_826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout647 _09350_/B vssd1 vssd1 vccd1 vccd1 _12447_/B sky130_fd_sc_hd__clkbuf_4
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09844_ _10241_/B _09843_/C _09843_/D _10694_/A vssd1 vssd1 vccd1 vccd1 _09845_/B
+ sky130_fd_sc_hd__a22oi_1
Xfanout658 _13802_/B vssd1 vssd1 vccd1 vccd1 _13632_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_59_848 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout669 _14865_/B vssd1 vssd1 vccd1 vccd1 _13993_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_86_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09775_ _09776_/A _09776_/B _09776_/C vssd1 vssd1 vccd1 vccd1 _09777_/A sky130_fd_sc_hd__a21oi_1
XFILLER_86_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08726_ _15402_/A vssd1 vssd1 vccd1 vccd1 _15274_/A sky130_fd_sc_hd__inv_2
XFILLER_73_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_36 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_973 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10550_ _10550_/A _10550_/B _10550_/C vssd1 vssd1 vccd1 vccd1 _10550_/X sky130_fd_sc_hd__and3_1
XFILLER_10_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09209_ _17407_/A _09555_/D _09209_/C vssd1 vssd1 vccd1 vccd1 _09373_/A sky130_fd_sc_hd__and3_1
XFILLER_154_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10481_ _10236_/B _11027_/C _11027_/D _10366_/A vssd1 vssd1 vccd1 vccd1 _10481_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_154_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12220_ _11826_/Y _11829_/Y _17365_/A vssd1 vssd1 vccd1 vccd1 _12220_/X sky130_fd_sc_hd__mux2_1
XFILLER_108_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12151_ _12316_/A _12151_/B _12151_/C vssd1 vssd1 vccd1 vccd1 _12316_/B sky130_fd_sc_hd__nand3_2
XFILLER_162_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11102_ _11238_/A _11238_/B vssd1 vssd1 vccd1 vccd1 _11104_/C sky130_fd_sc_hd__nand2_1
XFILLER_2_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12082_ _12082_/A _12082_/B vssd1 vssd1 vccd1 vccd1 _12083_/B sky130_fd_sc_hd__nor2_1
XFILLER_104_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_303 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11033_ _11005_/A _11005_/B _11007_/X _11006_/X _10805_/D vssd1 vssd1 vccd1 vccd1
+ _11035_/B sky130_fd_sc_hd__a32o_1
X_15910_ _16317_/A _16054_/B vssd1 vssd1 vccd1 vccd1 _16129_/B sky130_fd_sc_hd__and2_1
XFILLER_78_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16890_ _16890_/A _16952_/A vssd1 vssd1 vccd1 vccd1 _16895_/A sky130_fd_sc_hd__nand2_1
X_15841_ _15841_/A _15841_/B vssd1 vssd1 vccd1 vccd1 _15864_/A sky130_fd_sc_hd__xnor2_1
XFILLER_77_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_818 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12984_ _12984_/A _12984_/B vssd1 vssd1 vccd1 vccd1 _12985_/C sky130_fd_sc_hd__nand2_1
XFILLER_91_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15772_ _15772_/A _15772_/B _15772_/C vssd1 vssd1 vccd1 vccd1 _15773_/B sky130_fd_sc_hd__and3_1
XTAP_3541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17511_ fanout949/X _17511_/D vssd1 vssd1 vccd1 vccd1 _17511_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_851 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11935_ _11935_/A _11935_/B vssd1 vssd1 vccd1 vccd1 _11936_/B sky130_fd_sc_hd__nor2_1
X_14723_ _14723_/A _14723_/B _14723_/C vssd1 vssd1 vccd1 vccd1 _14726_/C sky130_fd_sc_hd__or3_1
XFILLER_91_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17442_ fanout938/X _17442_/D vssd1 vssd1 vccd1 vccd1 _17442_/Q sky130_fd_sc_hd__dfxtp_1
X_14654_ _14655_/A _14655_/B vssd1 vssd1 vccd1 vccd1 _14691_/A sky130_fd_sc_hd__nand2_1
XTAP_2884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11866_ _12077_/B _12077_/D _11867_/D _12077_/A vssd1 vssd1 vccd1 vccd1 _11868_/A
+ sky130_fd_sc_hd__a22oi_1
XTAP_2895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13605_ _13605_/A _13605_/B vssd1 vssd1 vccd1 vccd1 _13607_/C sky130_fd_sc_hd__xor2_1
X_10817_ _11097_/C _11115_/C _10812_/A _10810_/Y vssd1 vssd1 vccd1 vccd1 _10823_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_17373_ _17373_/A _17389_/B vssd1 vssd1 vccd1 vccd1 _17373_/X sky130_fd_sc_hd__or2_1
X_14585_ _14585_/A _14585_/B vssd1 vssd1 vccd1 vccd1 _14587_/B sky130_fd_sc_hd__nand2_1
XFILLER_159_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11797_ _14832_/A _17134_/A _17100_/C _14765_/A vssd1 vssd1 vccd1 vccd1 _11798_/D
+ sky130_fd_sc_hd__or4_1
XFILLER_13_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16324_ _16324_/A _16324_/B vssd1 vssd1 vccd1 vccd1 _16326_/A sky130_fd_sc_hd__nand2_1
XFILLER_13_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13536_ _13403_/B _13409_/B _13403_/A vssd1 vssd1 vccd1 vccd1 _13538_/B sky130_fd_sc_hd__a21boi_1
X_10748_ _11160_/A _11160_/B vssd1 vssd1 vccd1 vccd1 _10750_/C sky130_fd_sc_hd__nand2_1
XFILLER_159_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16255_ _16158_/A _16158_/B _16145_/Y vssd1 vssd1 vccd1 vccd1 _16257_/B sky130_fd_sc_hd__a21bo_1
XFILLER_145_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13467_ _13352_/B _13866_/D _13764_/D _14153_/A vssd1 vssd1 vccd1 vccd1 _13469_/A
+ sky130_fd_sc_hd__a22oi_1
X_10679_ _10681_/A _10681_/B vssd1 vssd1 vccd1 vccd1 _10679_/X sky130_fd_sc_hd__and2_1
XFILLER_173_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15206_ _15206_/A _15206_/B vssd1 vssd1 vccd1 vccd1 _15206_/X sky130_fd_sc_hd__and2_1
X_12418_ _12419_/A _12419_/B vssd1 vssd1 vccd1 vccd1 _12572_/B sky130_fd_sc_hd__and2_1
X_16186_ _16188_/A _16188_/B _16188_/C vssd1 vssd1 vccd1 vccd1 _16189_/A sky130_fd_sc_hd__o21a_1
XFILLER_154_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13398_ _13397_/Y _13526_/A _13398_/C vssd1 vssd1 vccd1 vccd1 _13526_/B sky130_fd_sc_hd__nand3b_1
XFILLER_154_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15137_ _15116_/B _14944_/A _15133_/X _15136_/X vssd1 vssd1 vccd1 vccd1 _17546_/D
+ sky130_fd_sc_hd__a22oi_1
X_12349_ _12349_/A _12349_/B vssd1 vssd1 vccd1 vccd1 _12350_/B sky130_fd_sc_hd__nand2_1
XFILLER_142_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15068_ _15274_/A _16977_/A _15065_/Y _15067_/X vssd1 vssd1 vccd1 vccd1 _17545_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_141_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14019_ _14113_/A _14019_/B vssd1 vssd1 vccd1 vccd1 _14021_/B sky130_fd_sc_hd__and2_1
XFILLER_4_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09560_ _09689_/A _09689_/B vssd1 vssd1 vccd1 vccd1 _09574_/C sky130_fd_sc_hd__and2_1
XFILLER_67_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09491_ _09491_/A _09491_/B vssd1 vssd1 vccd1 vccd1 _09619_/A sky130_fd_sc_hd__nor2_1
XFILLER_82_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_792 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout400 _12171_/A vssd1 vssd1 vccd1 vccd1 _17405_/A sky130_fd_sc_hd__buf_4
XFILLER_63_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout411 _09979_/A vssd1 vssd1 vccd1 vccd1 _10236_/A sky130_fd_sc_hd__buf_2
Xfanout422 _13948_/B vssd1 vssd1 vccd1 vccd1 _13632_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_87_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout433 _17527_/Q vssd1 vssd1 vccd1 vccd1 _14777_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_101_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout444 _10242_/A1 vssd1 vssd1 vccd1 vccd1 _12077_/B sky130_fd_sc_hd__buf_4
XFILLER_58_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout455 _17525_/Q vssd1 vssd1 vccd1 vccd1 _09412_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_86_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout466 _17523_/Q vssd1 vssd1 vccd1 vccd1 _12734_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_150_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout477 _10255_/A vssd1 vssd1 vccd1 vccd1 _11005_/A sky130_fd_sc_hd__clkbuf_4
X_09827_ _09827_/A _09827_/B vssd1 vssd1 vccd1 vccd1 _09968_/A sky130_fd_sc_hd__xnor2_1
XFILLER_24_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout488 _17521_/Q vssd1 vssd1 vccd1 vccd1 _15262_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_150_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout499 _12907_/A vssd1 vssd1 vccd1 vccd1 _09730_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_58_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09758_ _09758_/A _09758_/B vssd1 vssd1 vccd1 vccd1 _09890_/C sky130_fd_sc_hd__xnor2_1
XTAP_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09689_ _09689_/A _09689_/B vssd1 vssd1 vccd1 vccd1 _09718_/A sky130_fd_sc_hd__xnor2_1
XFILLER_73_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11720_ _11726_/A _11726_/B vssd1 vssd1 vccd1 vccd1 _11732_/A sky130_fd_sc_hd__or2_1
XTAP_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11651_ _11651_/A _15008_/B vssd1 vssd1 vccd1 vccd1 _11675_/C sky130_fd_sc_hd__nand2_2
XFILLER_168_720 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_34 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10602_ _10603_/A _10603_/B vssd1 vssd1 vccd1 vccd1 _10615_/A sky130_fd_sc_hd__nand2_1
X_14370_ _14370_/A _14370_/B vssd1 vssd1 vccd1 vccd1 _14372_/C sky130_fd_sc_hd__nor2_1
X_11582_ _11582_/A _11583_/A _11582_/C vssd1 vssd1 vccd1 vccd1 _11583_/B sky130_fd_sc_hd__nand3_1
XFILLER_168_775 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13321_ _14213_/A _13434_/B _13434_/D _13321_/D vssd1 vssd1 vccd1 vccd1 _13322_/B
+ sky130_fd_sc_hd__and4_1
X_10533_ _10851_/B _10647_/D _10745_/D _11122_/A vssd1 vssd1 vccd1 vccd1 _10533_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_127_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16040_ _16040_/A _16040_/B vssd1 vssd1 vccd1 vccd1 _16041_/C sky130_fd_sc_hd__xnor2_1
XFILLER_10_497 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13252_ _13252_/A vssd1 vssd1 vccd1 vccd1 _13252_/Y sky130_fd_sc_hd__inv_2
XFILLER_109_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10464_ _10465_/B _10465_/A vssd1 vssd1 vccd1 vccd1 _10467_/A sky130_fd_sc_hd__and2b_1
XFILLER_164_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12203_ _11967_/A _11971_/A _12371_/A _12202_/Y vssd1 vssd1 vccd1 vccd1 _12371_/B
+ sky130_fd_sc_hd__a211oi_2
XFILLER_89_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13183_ _13184_/A _13184_/B vssd1 vssd1 vccd1 vccd1 _13326_/A sky130_fd_sc_hd__and2_1
XFILLER_89_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10395_ _10395_/A _10505_/A vssd1 vssd1 vccd1 vccd1 _10397_/B sky130_fd_sc_hd__nor2_1
XFILLER_151_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12134_ _14356_/S _08967_/B _17134_/B _11849_/A vssd1 vssd1 vccd1 vccd1 _12136_/A
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_150_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16942_ _16943_/A _16943_/B vssd1 vssd1 vccd1 vccd1 _16994_/B sky130_fd_sc_hd__nand2_1
XFILLER_1_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12065_ _11849_/A _12058_/X _12064_/X _13625_/B vssd1 vssd1 vccd1 vccd1 _12065_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_150_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11016_ _11016_/A _11016_/B vssd1 vssd1 vccd1 vccd1 _11020_/A sky130_fd_sc_hd__xnor2_1
X_16873_ _11766_/X _16922_/A _16866_/Y _16872_/X vssd1 vssd1 vccd1 vccd1 _16873_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_93_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15824_ _15825_/A _15825_/B vssd1 vssd1 vccd1 vccd1 _15926_/A sky130_fd_sc_hd__nand2_1
XFILLER_64_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15755_ _16262_/A _15755_/B vssd1 vssd1 vccd1 vccd1 _15756_/B sky130_fd_sc_hd__nor2_1
X_12967_ _12968_/A _12968_/B vssd1 vssd1 vccd1 vccd1 _13107_/A sky130_fd_sc_hd__and2b_1
XFILLER_52_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11918_ _11914_/X _11916_/A _08874_/A _08873_/X vssd1 vssd1 vccd1 vccd1 _11918_/Y
+ sky130_fd_sc_hd__a211oi_1
X_14706_ _14735_/A1 _12548_/B _13625_/Y _12853_/X vssd1 vssd1 vccd1 vccd1 _14706_/X
+ sky130_fd_sc_hd__a31o_1
XTAP_2670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12898_ _13049_/A _12899_/B _12899_/C vssd1 vssd1 vccd1 vccd1 _12900_/A sky130_fd_sc_hd__a21o_1
XFILLER_60_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15686_ _15686_/A _15686_/B vssd1 vssd1 vccd1 vccd1 _15686_/Y sky130_fd_sc_hd__xnor2_1
XTAP_2681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17425_ _17425_/A _17425_/B vssd1 vssd1 vccd1 vccd1 _17425_/X sky130_fd_sc_hd__or2_1
XFILLER_21_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14637_ _14735_/A1 _12218_/A _13625_/Y _12853_/X vssd1 vssd1 vccd1 vccd1 _14637_/X
+ sky130_fd_sc_hd__a31o_1
X_11849_ _11849_/A _13626_/B vssd1 vssd1 vccd1 vccd1 _11849_/Y sky130_fd_sc_hd__nand2_1
XFILLER_21_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17356_ _11815_/B _17356_/A2 _17355_/X _17422_/C1 vssd1 vssd1 vccd1 vccd1 _17507_/D
+ sky130_fd_sc_hd__o211a_1
X_14568_ _14569_/A _14569_/B _14569_/C vssd1 vssd1 vccd1 vccd1 _14621_/A sky130_fd_sc_hd__a21o_1
XFILLER_158_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16307_ _16302_/B _16799_/A2 _16580_/B1 _16298_/A _16869_/C1 vssd1 vssd1 vccd1 vccd1
+ _16307_/X sky130_fd_sc_hd__a221o_1
XFILLER_9_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13519_ _14757_/S _13519_/B vssd1 vssd1 vccd1 vccd1 _13519_/Y sky130_fd_sc_hd__nor2_1
X_14499_ _17023_/A _14492_/A _14438_/B vssd1 vssd1 vccd1 vccd1 _14500_/B sky130_fd_sc_hd__o21ba_1
X_17287_ _17463_/Q _17290_/A2 _17285_/X _17286_/X _17293_/C1 vssd1 vssd1 vccd1 vccd1
+ _17463_/D sky130_fd_sc_hd__o221a_1
XFILLER_146_447 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16238_ _16238_/A _16238_/B vssd1 vssd1 vccd1 vccd1 _16239_/B sky130_fd_sc_hd__xor2_1
XFILLER_146_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16169_ _16695_/A _16589_/B _16065_/B _16352_/A vssd1 vssd1 vccd1 vccd1 _16170_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_142_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08991_ _08991_/A _08991_/B vssd1 vssd1 vccd1 vccd1 _08994_/A sky130_fd_sc_hd__xnor2_1
XFILLER_173_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09612_ _09755_/B _10309_/B _10311_/D _09755_/A vssd1 vssd1 vccd1 vccd1 _09612_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_83_412 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09543_ _09543_/A _09543_/B vssd1 vssd1 vccd1 vccd1 _09624_/A sky130_fd_sc_hd__xnor2_1
XFILLER_55_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09474_ _09478_/B _09474_/B vssd1 vssd1 vccd1 vccd1 _09602_/C sky130_fd_sc_hd__and2_1
XFILLER_93_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_740 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10180_ _10180_/A _10180_/B _10180_/C vssd1 vssd1 vccd1 vccd1 _10183_/A sky130_fd_sc_hd__and3_1
XFILLER_106_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout230 fanout230/A vssd1 vssd1 vccd1 vccd1 _17075_/A2 sky130_fd_sc_hd__clkbuf_4
Xfanout241 _14871_/Y vssd1 vssd1 vccd1 vccd1 _16401_/C1 sky130_fd_sc_hd__clkbuf_2
XFILLER_87_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout252 _15998_/A vssd1 vssd1 vccd1 vccd1 _17070_/B sky130_fd_sc_hd__clkbuf_8
Xfanout263 _17429_/C vssd1 vssd1 vccd1 vccd1 _17359_/C sky130_fd_sc_hd__clkbuf_2
Xfanout274 _15373_/B vssd1 vssd1 vccd1 vccd1 _16209_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_47_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_475 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout285 _08723_/Y vssd1 vssd1 vccd1 vccd1 _15275_/C1 sky130_fd_sc_hd__clkbuf_4
Xfanout296 _15130_/S vssd1 vssd1 vccd1 vccd1 _15312_/S sky130_fd_sc_hd__buf_4
X_13870_ _13870_/A _13870_/B vssd1 vssd1 vccd1 vccd1 _13873_/A sky130_fd_sc_hd__xnor2_1
XFILLER_28_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12821_ _12821_/A _12821_/B vssd1 vssd1 vccd1 vccd1 _12823_/B sky130_fd_sc_hd__or2_1
XFILLER_75_89 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12752_ _12907_/A _13051_/D vssd1 vssd1 vccd1 vccd1 _12754_/B sky130_fd_sc_hd__nand2_1
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15540_ _16012_/S _15537_/X _15539_/X _15808_/A vssd1 vssd1 vccd1 vccd1 _15540_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11703_ _11703_/A _11703_/B vssd1 vssd1 vccd1 vccd1 _11704_/B sky130_fd_sc_hd__xor2_2
X_15471_ _15472_/A _15472_/B vssd1 vssd1 vccd1 vccd1 _16604_/B sky130_fd_sc_hd__and2_4
XFILLER_42_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12683_ _12519_/A _12519_/B _12520_/Y vssd1 vssd1 vccd1 vccd1 _12685_/B sky130_fd_sc_hd__o21a_1
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17210_ _17579_/Q _17225_/A2 _17225_/B1 vssd1 vssd1 vccd1 vccd1 _17210_/X sky130_fd_sc_hd__a21o_1
X_14422_ _12849_/X _14210_/B _14482_/B1 vssd1 vssd1 vccd1 vccd1 _14422_/X sky130_fd_sc_hd__o21a_1
X_11634_ _11635_/B _11635_/A vssd1 vssd1 vccd1 vccd1 _11662_/A sky130_fd_sc_hd__nand2b_1
XFILLER_156_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14353_ _14416_/B _14354_/B vssd1 vssd1 vccd1 vccd1 _14353_/Y sky130_fd_sc_hd__nand2_1
X_17141_ _14829_/X _17162_/A2 _16974_/B _14829_/B _17162_/C1 vssd1 vssd1 vccd1 vccd1
+ _17141_/X sky130_fd_sc_hd__a221o_1
X_11565_ _11565_/A _11565_/B _11566_/B vssd1 vssd1 vccd1 vccd1 _11610_/A sky130_fd_sc_hd__or3_1
XFILLER_156_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13304_ _13304_/A _13304_/B vssd1 vssd1 vccd1 vccd1 _13306_/B sky130_fd_sc_hd__xor2_1
XFILLER_155_244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10516_ _10502_/X _10503_/Y _10510_/X _10514_/X vssd1 vssd1 vccd1 vccd1 _10517_/B
+ sky130_fd_sc_hd__a211o_1
X_17072_ _17065_/A _17029_/B _17140_/A vssd1 vssd1 vccd1 vccd1 _17072_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_156_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14284_ _14283_/B _14284_/B vssd1 vssd1 vccd1 vccd1 _14352_/B sky130_fd_sc_hd__and2b_1
XFILLER_109_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11496_ _11496_/A _11496_/B vssd1 vssd1 vccd1 vccd1 _11497_/B sky130_fd_sc_hd__nand2_1
XFILLER_143_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16023_ _16938_/A _17119_/C vssd1 vssd1 vccd1 vccd1 _16023_/Y sky130_fd_sc_hd__nand2_1
XFILLER_6_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13235_ _13235_/A _13235_/B vssd1 vssd1 vccd1 vccd1 _13238_/A sky130_fd_sc_hd__xor2_1
XFILLER_40_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10447_ _10560_/B _10446_/B _10446_/C vssd1 vssd1 vccd1 vccd1 _10448_/B sky130_fd_sc_hd__a21oi_1
XFILLER_124_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13166_ _13036_/A _13038_/B _13036_/B vssd1 vssd1 vccd1 vccd1 _13176_/A sky130_fd_sc_hd__o21ba_1
X_10378_ _11006_/B _10799_/B _14788_/B _10954_/A vssd1 vssd1 vccd1 vccd1 _10379_/B
+ sky130_fd_sc_hd__a22oi_1
XFILLER_151_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12117_ _12118_/A _12118_/B _12118_/C vssd1 vssd1 vccd1 vccd1 _12309_/A sky130_fd_sc_hd__a21o_1
XFILLER_112_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13097_ _14153_/B _13551_/D _13434_/D _14153_/A vssd1 vssd1 vccd1 vccd1 _13099_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_111_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16925_ _16918_/B _17162_/A2 _16974_/B _13993_/B _17162_/C1 vssd1 vssd1 vccd1 vccd1
+ _16925_/X sky130_fd_sc_hd__a221o_1
X_12048_ _12487_/D _12320_/D _12050_/S vssd1 vssd1 vccd1 vccd1 _12049_/B sky130_fd_sc_hd__mux2_1
XFILLER_77_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_20 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16856_ _16931_/A _16931_/B _17131_/A vssd1 vssd1 vccd1 vccd1 _16856_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_92_220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15807_ _16011_/A _15180_/X _15628_/A vssd1 vssd1 vccd1 vccd1 _15808_/B sky130_fd_sc_hd__o21a_1
XFILLER_37_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16787_ _16787_/A _16853_/C vssd1 vssd1 vccd1 vccd1 _16787_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_65_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13999_ _13897_/A _14485_/D _13898_/A _13896_/B vssd1 vssd1 vccd1 vccd1 _14001_/B
+ sky130_fd_sc_hd__a31o_1
XTAP_3190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15738_ _15647_/A _16152_/A _15644_/X _15645_/Y vssd1 vssd1 vccd1 vccd1 _15740_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_52_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15669_ _15568_/A _15570_/B _15568_/B vssd1 vssd1 vccd1 vccd1 _15671_/B sky130_fd_sc_hd__a21bo_1
XFILLER_21_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_695 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17408_ input50/X _17422_/A2 _17407_/X _17408_/C1 vssd1 vssd1 vccd1 vccd1 _17532_/D
+ sky130_fd_sc_hd__o211a_1
X_09190_ _09190_/A _09221_/B vssd1 vssd1 vccd1 vccd1 _09196_/A sky130_fd_sc_hd__nor2_1
XFILLER_60_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1015 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17339_ input49/X _17353_/B _17353_/C vssd1 vssd1 vccd1 vccd1 _17339_/X sky130_fd_sc_hd__or3_1
XFILLER_119_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08974_ _09242_/A _08974_/B vssd1 vssd1 vccd1 vccd1 _08983_/A sky130_fd_sc_hd__and2_1
XFILLER_130_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1046 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_795 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09526_ _09507_/Y _09525_/X _09487_/X _09488_/Y vssd1 vssd1 vccd1 vccd1 _09530_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_71_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09457_ _09455_/A _09455_/B _09543_/B _09437_/X vssd1 vssd1 vccd1 vccd1 _09483_/B
+ sky130_fd_sc_hd__a31oi_1
XPHY_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_504 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09388_ _09388_/A vssd1 vssd1 vccd1 vccd1 _09388_/Y sky130_fd_sc_hd__inv_2
XFILLER_138_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_570 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11350_ _11291_/B _11288_/C _11288_/A vssd1 vssd1 vccd1 vccd1 _11351_/C sky130_fd_sc_hd__a21o_1
XFILLER_153_704 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10301_ _10301_/A _10301_/B vssd1 vssd1 vccd1 vccd1 _10411_/B sky130_fd_sc_hd__xnor2_1
X_11281_ _11281_/A _11281_/B _11281_/C vssd1 vssd1 vccd1 vccd1 _11333_/A sky130_fd_sc_hd__and3_1
X_13020_ _13950_/A _14213_/C vssd1 vssd1 vccd1 vccd1 _13021_/B sky130_fd_sc_hd__nand2_1
XFILLER_3_246 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10232_ _10232_/A _10232_/B vssd1 vssd1 vccd1 vccd1 _10261_/A sky130_fd_sc_hd__xnor2_1
XFILLER_152_269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10163_ _10163_/A _10163_/B vssd1 vssd1 vccd1 vccd1 _10177_/A sky130_fd_sc_hd__nand2_1
XFILLER_121_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14971_ _15147_/C _11789_/X _14877_/Y vssd1 vssd1 vccd1 vccd1 _14971_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_250 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10094_ _10094_/A _10348_/A vssd1 vssd1 vccd1 vccd1 _10097_/B sky130_fd_sc_hd__nor2_1
XFILLER_47_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16710_ _16711_/A _16711_/B _16711_/C vssd1 vssd1 vccd1 vccd1 _16786_/A sky130_fd_sc_hd__o21ai_1
XFILLER_102_892 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13922_ _13922_/A _13922_/B vssd1 vssd1 vccd1 vccd1 _13923_/B sky130_fd_sc_hd__nand2_1
XFILLER_19_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16641_ _16641_/A _16641_/B vssd1 vssd1 vccd1 vccd1 _16641_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_74_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13853_ _13853_/A _13853_/B vssd1 vssd1 vccd1 vccd1 _13856_/A sky130_fd_sc_hd__xor2_1
XFILLER_90_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12804_ _12804_/A _12804_/B _13321_/D _13194_/D vssd1 vssd1 vccd1 vccd1 _12805_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_90_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16572_ _16572_/A _16572_/B vssd1 vssd1 vccd1 vccd1 _16572_/Y sky130_fd_sc_hd__nand2_1
X_10996_ _11164_/B _10996_/B _10996_/C vssd1 vssd1 vccd1 vccd1 _11159_/A sky130_fd_sc_hd__or3_1
X_13784_ _13784_/A _13784_/B vssd1 vssd1 vccd1 vccd1 _13785_/B sky130_fd_sc_hd__and2_1
XFILLER_163_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15523_ _15523_/A _15523_/B vssd1 vssd1 vccd1 vccd1 _15523_/X sky130_fd_sc_hd__or2_1
X_12735_ _12735_/A _12735_/B vssd1 vssd1 vccd1 vccd1 _12737_/A sky130_fd_sc_hd__nor2_1
XFILLER_35_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_982 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_8 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12666_ _12509_/B _12511_/B _12509_/A vssd1 vssd1 vccd1 vccd1 _12668_/B sky130_fd_sc_hd__o21ba_1
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15454_ _15454_/A _15454_/B _15532_/B vssd1 vssd1 vccd1 vccd1 _15454_/X sky130_fd_sc_hd__and3_1
XFILLER_30_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11617_ _11617_/A _11617_/B _11617_/C vssd1 vssd1 vccd1 vccd1 _11672_/A sky130_fd_sc_hd__or3_1
X_14405_ _14405_/A _14405_/B _14405_/C vssd1 vssd1 vccd1 vccd1 _14424_/B sky130_fd_sc_hd__and3_1
X_12597_ _12907_/A _13037_/B vssd1 vssd1 vccd1 vccd1 _12599_/B sky130_fd_sc_hd__and2_1
XFILLER_30_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15385_ _12858_/Y _17164_/D _15384_/X _16011_/A vssd1 vssd1 vccd1 vccd1 _15386_/B
+ sky130_fd_sc_hd__o22ai_2
X_17124_ _17124_/A _17124_/B vssd1 vssd1 vccd1 vccd1 _17125_/B sky130_fd_sc_hd__or2_1
X_11548_ _11705_/A _11547_/C _11586_/A vssd1 vssd1 vccd1 vccd1 _11549_/B sky130_fd_sc_hd__a21bo_1
X_14336_ _14405_/A _14337_/C _14337_/A vssd1 vssd1 vccd1 vccd1 _14336_/X sky130_fd_sc_hd__o21a_1
XFILLER_156_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17055_ _17093_/B _17055_/B vssd1 vssd1 vccd1 vccd1 _17057_/B sky130_fd_sc_hd__xor2_1
X_14267_ _14268_/A _14268_/B vssd1 vssd1 vccd1 vccd1 _14344_/B sky130_fd_sc_hd__and2_1
X_11479_ _11479_/A _11479_/B vssd1 vssd1 vccd1 vccd1 _11484_/A sky130_fd_sc_hd__nor2_1
XFILLER_171_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13218_ _13346_/B _13218_/B vssd1 vssd1 vccd1 vccd1 _13220_/C sky130_fd_sc_hd__nand2_1
X_16006_ _17119_/B _16005_/B _16005_/C vssd1 vssd1 vccd1 vccd1 _16007_/C sky130_fd_sc_hd__a21oi_1
X_14198_ _14276_/A _14198_/B vssd1 vssd1 vccd1 vccd1 _14198_/X sky130_fd_sc_hd__or2_1
XFILLER_98_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13149_ _13149_/A _13149_/B vssd1 vssd1 vccd1 vccd1 _13151_/A sky130_fd_sc_hd__nor2_1
XFILLER_83_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_924 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16908_ _16908_/A _16908_/B vssd1 vssd1 vccd1 vccd1 _16909_/B sky130_fd_sc_hd__xnor2_1
XFILLER_111_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16839_ _16775_/A _16775_/B _16771_/A vssd1 vssd1 vccd1 vccd1 _16841_/B sky130_fd_sc_hd__a21bo_1
XFILLER_93_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_595 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09311_ _09311_/A _09316_/B _09311_/C vssd1 vssd1 vccd1 vccd1 _09401_/A sky130_fd_sc_hd__and3_1
XFILLER_22_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09242_ _09242_/A _09242_/B _09242_/C vssd1 vssd1 vccd1 vccd1 _09243_/B sky130_fd_sc_hd__nand3_1
XFILLER_21_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09173_ _09360_/A _10446_/B _09502_/C vssd1 vssd1 vccd1 vccd1 _09357_/A sky130_fd_sc_hd__and3_1
XFILLER_31_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_704 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08957_ _11932_/A _11895_/C _08957_/C _08957_/D vssd1 vssd1 vccd1 vccd1 _09084_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_29_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08888_ _16315_/A _08888_/B vssd1 vssd1 vccd1 vccd1 _09020_/A sky130_fd_sc_hd__xnor2_1
XFILLER_5_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10850_ _10850_/A _10855_/A _10850_/C vssd1 vssd1 vccd1 vccd1 _10859_/B sky130_fd_sc_hd__or3_1
XFILLER_72_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09509_ _10559_/A _09555_/D vssd1 vssd1 vccd1 vccd1 _09524_/A sky130_fd_sc_hd__nand2_1
XFILLER_169_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10781_ _10682_/Y _10689_/X _10779_/B _10780_/Y vssd1 vssd1 vccd1 vccd1 _10784_/B
+ sky130_fd_sc_hd__o31a_2
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_695 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12520_ _12521_/B _12521_/A vssd1 vssd1 vccd1 vccd1 _12520_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_158_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12451_ _12451_/A _12451_/B vssd1 vssd1 vccd1 vccd1 _12452_/B sky130_fd_sc_hd__xnor2_1
XFILLER_12_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11402_ _11402_/A _11402_/B _11451_/A vssd1 vssd1 vccd1 vccd1 _11408_/A sky130_fd_sc_hd__nor3b_1
XFILLER_172_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15170_ _15170_/A _15170_/B _15170_/C vssd1 vssd1 vccd1 vccd1 _15171_/B sky130_fd_sc_hd__and3_1
X_12382_ _12042_/Y _12044_/Y _12383_/S vssd1 vssd1 vccd1 vccd1 _12382_/X sky130_fd_sc_hd__mux2_1
XANTENNA_90 _10016_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14121_ _14032_/A _14029_/Y _14031_/B vssd1 vssd1 vccd1 vccd1 _14121_/X sky130_fd_sc_hd__o21a_1
X_11333_ _11333_/A _11333_/B vssd1 vssd1 vccd1 vccd1 _11340_/A sky130_fd_sc_hd__nor2_1
XFILLER_21_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14052_ _14215_/A _14213_/D vssd1 vssd1 vccd1 vccd1 _14054_/B sky130_fd_sc_hd__nand2_1
X_11264_ _11264_/A _11270_/A _11264_/C vssd1 vssd1 vccd1 vccd1 _11274_/B sky130_fd_sc_hd__or3_1
XFILLER_153_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13003_ _13003_/A _13003_/B vssd1 vssd1 vccd1 vccd1 _13004_/B sky130_fd_sc_hd__or2_1
XFILLER_134_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10215_ _10214_/A _10215_/B vssd1 vssd1 vccd1 vccd1 _10216_/C sky130_fd_sc_hd__nand2b_1
XFILLER_106_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11195_ _11195_/A _11195_/B vssd1 vssd1 vccd1 vccd1 _11198_/A sky130_fd_sc_hd__xnor2_1
XFILLER_133_291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10146_ _10271_/A _10146_/B _10268_/B vssd1 vssd1 vccd1 vccd1 _10148_/C sky130_fd_sc_hd__and3_1
XFILLER_130_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10077_ _10033_/B _10055_/B _10033_/A vssd1 vssd1 vccd1 vccd1 _10080_/A sky130_fd_sc_hd__o21bai_1
X_14954_ _14954_/A _15038_/B vssd1 vssd1 vccd1 vccd1 _14954_/Y sky130_fd_sc_hd__nor2_1
XFILLER_94_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_787 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13905_ _13906_/A _13906_/B _13906_/C vssd1 vssd1 vccd1 vccd1 _14027_/A sky130_fd_sc_hd__a21oi_1
XFILLER_63_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14885_ _15396_/A _14888_/B _14888_/C _14888_/D vssd1 vssd1 vccd1 vccd1 _14886_/D
+ sky130_fd_sc_hd__or4_1
X_16624_ _16625_/A _16625_/B _16623_/X vssd1 vssd1 vccd1 vccd1 _16624_/X sky130_fd_sc_hd__o21ba_1
X_13836_ _14756_/A1 _13829_/Y _13830_/X _13835_/X vssd1 vssd1 vccd1 vccd1 _17590_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_51_919 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16555_ _16557_/A _16557_/B _16557_/C vssd1 vssd1 vccd1 vccd1 _16638_/A sky130_fd_sc_hd__o21a_1
XFILLER_50_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10979_ _11049_/A _11049_/B _11049_/C vssd1 vssd1 vccd1 vccd1 _11051_/A sky130_fd_sc_hd__o21ai_2
X_13767_ _13767_/A _13767_/B vssd1 vssd1 vccd1 vccd1 _13768_/B sky130_fd_sc_hd__xnor2_1
XFILLER_31_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_807 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15506_ _16056_/A _16812_/A _15414_/A _15416_/Y vssd1 vssd1 vccd1 vccd1 _15507_/B
+ sky130_fd_sc_hd__a31o_1
X_12718_ _12871_/A _13334_/C _12557_/X _12869_/C _12235_/C vssd1 vssd1 vccd1 vccd1
+ _12720_/B sky130_fd_sc_hd__a32o_1
XFILLER_148_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16486_ _12560_/A _14775_/X _14816_/X _16485_/Y vssd1 vssd1 vccd1 vccd1 _16493_/B
+ sky130_fd_sc_hd__a31o_1
X_13698_ _14176_/A _16859_/A _13698_/C vssd1 vssd1 vccd1 vccd1 _13800_/B sky130_fd_sc_hd__nand3_1
XFILLER_30_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15437_ _15358_/A _15358_/B _15356_/A vssd1 vssd1 vccd1 vccd1 _15439_/B sky130_fd_sc_hd__o21ai_1
XFILLER_129_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12649_ _12650_/B _12649_/B vssd1 vssd1 vccd1 vccd1 _12651_/A sky130_fd_sc_hd__nand2b_1
XFILLER_30_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15368_ _15233_/X _15299_/Y _15298_/Y vssd1 vssd1 vccd1 vccd1 _15369_/B sky130_fd_sc_hd__o21bai_1
XFILLER_11_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17107_ _11775_/Y _17105_/Y _17106_/Y vssd1 vssd1 vccd1 vccd1 _17107_/X sky130_fd_sc_hd__a21o_1
X_14319_ _14319_/A _14389_/A vssd1 vssd1 vccd1 vccd1 _14321_/C sky130_fd_sc_hd__nor2_1
XFILLER_7_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15299_ _15299_/A _15299_/B vssd1 vssd1 vccd1 vccd1 _15299_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_116_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_718 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17038_ _17081_/A _17038_/B _17038_/C vssd1 vssd1 vccd1 vccd1 _17040_/B sky130_fd_sc_hd__nor3_1
XFILLER_144_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout807 _12158_/D vssd1 vssd1 vccd1 vccd1 _12340_/B sky130_fd_sc_hd__buf_4
X_09860_ _09994_/A _15801_/A _09855_/X vssd1 vssd1 vccd1 vccd1 _09862_/B sky130_fd_sc_hd__o21ba_2
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout818 _09265_/C vssd1 vssd1 vccd1 vccd1 _12923_/D sky130_fd_sc_hd__clkbuf_4
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout829 _14851_/A vssd1 vssd1 vccd1 vccd1 _15463_/A sky130_fd_sc_hd__buf_4
XFILLER_140_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08811_ _17397_/A _17395_/A _11861_/B _11859_/D vssd1 vssd1 vccd1 vccd1 _08812_/B
+ sky130_fd_sc_hd__and4_1
X_09791_ _10559_/A _09843_/D vssd1 vssd1 vccd1 vccd1 _09808_/A sky130_fd_sc_hd__nand2_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_838 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08742_ _17607_/Q _17608_/Q vssd1 vssd1 vccd1 vccd1 _14872_/A sky130_fd_sc_hd__or2_1
XFILLER_38_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09225_ _09225_/A _09225_/B vssd1 vssd1 vccd1 vccd1 _09227_/C sky130_fd_sc_hd__xor2_1
XFILLER_158_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_840 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09156_ _09152_/A _09153_/X _09131_/X _09138_/X vssd1 vssd1 vccd1 vccd1 _09156_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_147_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09087_ _09317_/A _09086_/Y _09327_/C _11895_/D vssd1 vssd1 vccd1 vccd1 _09323_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_174_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_910 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10000_ _10000_/A _10000_/B vssd1 vssd1 vccd1 vccd1 _10123_/B sky130_fd_sc_hd__nor2_1
XFILLER_88_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09989_ _09989_/A _09989_/B vssd1 vssd1 vccd1 vccd1 _10106_/B sky130_fd_sc_hd__xnor2_1
XFILLER_88_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_242 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11951_ _09014_/A _09013_/B _09013_/A vssd1 vssd1 vccd1 vccd1 _11993_/A sky130_fd_sc_hd__o21ba_1
XFILLER_83_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10902_ _10995_/B _10902_/B _10902_/C vssd1 vssd1 vccd1 vccd1 _10953_/A sky130_fd_sc_hd__or3_1
XFILLER_17_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11882_ _11882_/A _11882_/B vssd1 vssd1 vccd1 vccd1 _11884_/A sky130_fd_sc_hd__nor2_1
XFILLER_45_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14670_ _14633_/A _14631_/B _14669_/B _14669_/X vssd1 vssd1 vccd1 vccd1 _14670_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_72_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10833_ _10933_/A _11122_/B _10970_/B _10971_/B vssd1 vssd1 vccd1 vccd1 _10836_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_44_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13621_ _13729_/B _13621_/B vssd1 vssd1 vccd1 vccd1 _13621_/X sky130_fd_sc_hd__or2_1
XFILLER_72_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_1023 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16340_ _16444_/A _16340_/B vssd1 vssd1 vccd1 vccd1 _16342_/B sky130_fd_sc_hd__nor2_1
XFILLER_25_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10764_ _10771_/B _10764_/B vssd1 vssd1 vccd1 vccd1 _10764_/X sky130_fd_sc_hd__or2_1
X_13552_ _13552_/A _13680_/A vssd1 vssd1 vccd1 vccd1 _13555_/A sky130_fd_sc_hd__or2_1
XFILLER_160_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12503_ _12804_/A _12804_/B _13067_/D _12923_/D vssd1 vssd1 vccd1 vccd1 _12504_/B
+ sky130_fd_sc_hd__and4_1
X_16271_ _16271_/A _16271_/B vssd1 vssd1 vccd1 vccd1 _16272_/B sky130_fd_sc_hd__nor2_1
X_13483_ _13603_/A _13483_/B vssd1 vssd1 vccd1 vccd1 _13485_/B sky130_fd_sc_hd__nand2_1
XFILLER_40_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10695_ _11027_/B _11006_/C vssd1 vssd1 vccd1 vccd1 _11036_/A sky130_fd_sc_hd__nand2_1
XFILLER_12_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_647 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12434_ _12588_/A _12434_/B _12434_/C vssd1 vssd1 vccd1 vccd1 _12588_/B sky130_fd_sc_hd__nand3_2
X_15222_ _15222_/A _15222_/B vssd1 vssd1 vccd1 vccd1 _15225_/A sky130_fd_sc_hd__nand2_1
XFILLER_173_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15153_ _14881_/X _14889_/X _15932_/A _15275_/C1 vssd1 vssd1 vccd1 vccd1 _15155_/B
+ sky130_fd_sc_hd__a211o_1
X_12365_ _12364_/A _12364_/B _12364_/C vssd1 vssd1 vccd1 vccd1 _12366_/B sky130_fd_sc_hd__a21oi_1
XFILLER_126_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11316_ _15373_/C _11592_/B _17467_/D _11370_/A vssd1 vssd1 vccd1 vccd1 _11317_/B
+ sky130_fd_sc_hd__a22o_1
X_14104_ _14104_/A _14104_/B vssd1 vssd1 vccd1 vccd1 _14105_/B sky130_fd_sc_hd__or2_1
X_15084_ _15081_/A _15734_/A _15157_/A _15083_/X vssd1 vssd1 vccd1 vccd1 _15085_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_126_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12296_ _12296_/A _12508_/A vssd1 vssd1 vccd1 vccd1 _12299_/A sky130_fd_sc_hd__or2_1
XFILLER_5_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_770 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14035_ _14763_/S _14033_/X _14034_/Y _13945_/Y vssd1 vssd1 vccd1 vccd1 _17592_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_107_792 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11247_ _11308_/A _11308_/B vssd1 vssd1 vccd1 vccd1 _11249_/C sky130_fd_sc_hd__and2b_1
XFILLER_79_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11178_ _11015_/X _11019_/X _11175_/Y _11176_/X vssd1 vssd1 vccd1 vccd1 _11178_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_79_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10129_ _10255_/A _10270_/B vssd1 vssd1 vccd1 vccd1 _10251_/B sky130_fd_sc_hd__nand2_1
XFILLER_110_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_808 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15986_ _15987_/A _15987_/B vssd1 vssd1 vccd1 vccd1 _16096_/A sky130_fd_sc_hd__and2b_1
XFILLER_94_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14937_ _17607_/Q _14938_/B vssd1 vssd1 vccd1 vccd1 _15454_/A sky130_fd_sc_hd__nor2_1
XFILLER_82_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14868_ _17139_/A _17139_/B vssd1 vssd1 vccd1 vccd1 _17140_/B sky130_fd_sc_hd__and2_1
XFILLER_35_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16607_ _16607_/A _16607_/B vssd1 vssd1 vccd1 vccd1 _16609_/C sky130_fd_sc_hd__xor2_1
XFILLER_23_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_982 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13819_ _13820_/A _13820_/B vssd1 vssd1 vccd1 vccd1 _13930_/A sky130_fd_sc_hd__and2b_1
XFILLER_51_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17587_ fanout940/X _17587_/D vssd1 vssd1 vccd1 vccd1 _17587_/Q sky130_fd_sc_hd__dfxtp_1
X_14799_ _14790_/Y _14798_/Y _11321_/X vssd1 vssd1 vccd1 vccd1 _15244_/C sky130_fd_sc_hd__o21ba_1
XFILLER_51_749 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16538_ _16447_/Y _16450_/B _16446_/X vssd1 vssd1 vccd1 vccd1 _16541_/B sky130_fd_sc_hd__o21ai_1
XFILLER_32_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16469_ _16469_/A _16469_/B vssd1 vssd1 vccd1 vccd1 _16470_/C sky130_fd_sc_hd__xor2_2
XFILLER_31_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_607 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09010_ _09010_/A _09010_/B vssd1 vssd1 vccd1 vccd1 _09012_/C sky130_fd_sc_hd__nand2_1
XFILLER_136_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09912_ _09912_/A _09912_/B _09912_/C vssd1 vssd1 vccd1 vccd1 _09913_/B sky130_fd_sc_hd__or3_1
XFILLER_144_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout604 _17511_/Q vssd1 vssd1 vccd1 vccd1 _14982_/A sky130_fd_sc_hd__buf_2
Xfanout615 _17510_/Q vssd1 vssd1 vccd1 vccd1 _11132_/B sky130_fd_sc_hd__clkbuf_2
Xfanout626 _14829_/B vssd1 vssd1 vccd1 vccd1 _13051_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_113_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09843_ _10694_/A _10241_/B _09843_/C _09843_/D vssd1 vssd1 vccd1 vccd1 _09845_/A
+ sky130_fd_sc_hd__and4_1
Xfanout637 _15033_/A3 vssd1 vssd1 vccd1 vccd1 _14867_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_112_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout648 _14765_/B vssd1 vssd1 vccd1 vccd1 _09350_/B sky130_fd_sc_hd__clkbuf_4
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout659 _17504_/Q vssd1 vssd1 vccd1 vccd1 _13802_/B sky130_fd_sc_hd__clkbuf_4
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09774_ _09774_/A _09774_/B vssd1 vssd1 vccd1 vccd1 _09776_/C sky130_fd_sc_hd__xnor2_1
XTAP_3008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_702 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08725_ _14893_/B vssd1 vssd1 vccd1 vccd1 _15206_/A sky130_fd_sc_hd__inv_2
XTAP_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_985 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09208_ _09208_/A _09208_/B vssd1 vssd1 vccd1 vccd1 _09209_/C sky130_fd_sc_hd__xnor2_1
X_10480_ _10480_/A _10480_/B vssd1 vssd1 vccd1 vccd1 _10597_/A sky130_fd_sc_hd__xnor2_1
XFILLER_136_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09139_ _09139_/A _09139_/B vssd1 vssd1 vccd1 vccd1 _09150_/A sky130_fd_sc_hd__nor2_1
X_12150_ _12150_/A _12150_/B vssd1 vssd1 vccd1 vccd1 _12151_/C sky130_fd_sc_hd__xnor2_1
XFILLER_118_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11101_ _11101_/A _11101_/B vssd1 vssd1 vccd1 vccd1 _11238_/B sky130_fd_sc_hd__xnor2_1
XFILLER_1_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12081_ _12082_/A _12082_/B vssd1 vssd1 vccd1 vccd1 _12252_/B sky130_fd_sc_hd__and2_1
XFILLER_89_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11032_ _11032_/A _11032_/B vssd1 vssd1 vccd1 vccd1 _11035_/A sky130_fd_sc_hd__xnor2_1
XFILLER_1_366 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15840_ _15841_/A _15841_/B vssd1 vssd1 vccd1 vccd1 _15840_/Y sky130_fd_sc_hd__nand2_1
XFILLER_94_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15771_ _15772_/A _15772_/B _15772_/C vssd1 vssd1 vccd1 vccd1 _15773_/A sky130_fd_sc_hd__a21oi_1
XTAP_3531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12983_ _12982_/B _12983_/B vssd1 vssd1 vccd1 vccd1 _12984_/B sky130_fd_sc_hd__nand2b_1
XTAP_3542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17510_ fanout949/X _17510_/D vssd1 vssd1 vccd1 vccd1 _17510_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_73_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_543 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14722_ _14723_/A _14723_/B _14723_/C vssd1 vssd1 vccd1 vccd1 _14750_/A sky130_fd_sc_hd__o21ai_1
XTAP_3564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11934_ _11935_/A _11935_/B vssd1 vssd1 vccd1 vccd1 _11936_/A sky130_fd_sc_hd__and2_1
XTAP_3575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17441_ fanout937/X _17441_/D vssd1 vssd1 vccd1 vccd1 _17441_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_150_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14653_ _14693_/B _14653_/B vssd1 vssd1 vccd1 vccd1 _14655_/B sky130_fd_sc_hd__xnor2_1
XTAP_2874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11865_ _11865_/A _11865_/B vssd1 vssd1 vccd1 vccd1 _11874_/A sky130_fd_sc_hd__xor2_1
XTAP_2885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13604_ _13604_/A _13604_/B vssd1 vssd1 vccd1 vccd1 _13605_/B sky130_fd_sc_hd__nor2_1
X_10816_ _10816_/A _10816_/B vssd1 vssd1 vccd1 vccd1 _11072_/A sky130_fd_sc_hd__xnor2_1
X_17372_ input62/X _17377_/B _17371_/Y _17378_/C1 vssd1 vssd1 vccd1 vccd1 _17514_/D
+ sky130_fd_sc_hd__o211a_1
X_14584_ _14584_/A _14584_/B vssd1 vssd1 vccd1 vccd1 _14629_/C sky130_fd_sc_hd__nor2_1
X_11796_ _14766_/A _14554_/A _16913_/C _14383_/A vssd1 vssd1 vccd1 vccd1 _11798_/C
+ sky130_fd_sc_hd__or4_1
XFILLER_14_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16323_ _16410_/A _16595_/A _16662_/C _16662_/D vssd1 vssd1 vccd1 vccd1 _16324_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_14_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13535_ _13535_/A _13535_/B vssd1 vssd1 vccd1 vccd1 _13538_/A sky130_fd_sc_hd__xnor2_1
X_10747_ _10747_/A _10747_/B vssd1 vssd1 vccd1 vccd1 _11160_/B sky130_fd_sc_hd__xnor2_1
XFILLER_41_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16254_ _16254_/A _16254_/B vssd1 vssd1 vccd1 vccd1 _16257_/A sky130_fd_sc_hd__xor2_1
X_10678_ _10678_/A _10678_/B vssd1 vssd1 vccd1 vccd1 _10681_/B sky130_fd_sc_hd__nand2_1
X_13466_ _13322_/A _13324_/B _13322_/B vssd1 vssd1 vccd1 vccd1 _13473_/A sky130_fd_sc_hd__o21ba_1
XFILLER_174_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15205_ _15205_/A _15205_/B vssd1 vssd1 vccd1 vccd1 _15206_/B sky130_fd_sc_hd__nor2_1
XFILLER_126_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12417_ _12417_/A _12417_/B vssd1 vssd1 vccd1 vccd1 _12419_/B sky130_fd_sc_hd__xnor2_1
XFILLER_154_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16185_ _16165_/A _16533_/B _16060_/A _16058_/A vssd1 vssd1 vccd1 vccd1 _16188_/C
+ sky130_fd_sc_hd__a31o_1
X_13397_ _13846_/A _13522_/D vssd1 vssd1 vccd1 vccd1 _13397_/Y sky130_fd_sc_hd__nand2_1
XFILLER_142_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15136_ _15628_/A _15104_/X _15135_/Y _15808_/A vssd1 vssd1 vccd1 vccd1 _15136_/X
+ sky130_fd_sc_hd__a211o_1
X_12348_ _12349_/A _12349_/B vssd1 vssd1 vccd1 vccd1 _12517_/A sky130_fd_sc_hd__or2_1
XFILLER_154_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12279_ _12108_/A _12110_/B _12108_/B vssd1 vssd1 vccd1 vccd1 _12281_/B sky130_fd_sc_hd__o21ba_1
XFILLER_4_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15067_ _17131_/A _15093_/B _15031_/X _15066_/Y vssd1 vssd1 vccd1 vccd1 _15067_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_114_559 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14018_ _14018_/A _14018_/B _14018_/C vssd1 vssd1 vccd1 vccd1 _14019_/B sky130_fd_sc_hd__nand3_1
XFILLER_68_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15969_ _15969_/A _15969_/B vssd1 vssd1 vccd1 vccd1 _15970_/B sky130_fd_sc_hd__nor2_1
X_09490_ _09654_/C _11813_/B _09353_/A _09351_/Y vssd1 vssd1 vccd1 vccd1 _09491_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_63_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout401 _10559_/A vssd1 vssd1 vccd1 vccd1 _10560_/B sky130_fd_sc_hd__buf_2
Xfanout412 _17530_/Q vssd1 vssd1 vccd1 vccd1 _09979_/A sky130_fd_sc_hd__clkbuf_2
Xfanout423 _12869_/A vssd1 vssd1 vccd1 vccd1 _13948_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_99_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout434 _12077_/A vssd1 vssd1 vccd1 vccd1 _17397_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_101_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1006 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout445 _10241_/B vssd1 vssd1 vccd1 vccd1 _11027_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_86_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout456 _13035_/A vssd1 vssd1 vccd1 vccd1 _13658_/A sky130_fd_sc_hd__buf_2
Xfanout467 _08791_/B vssd1 vssd1 vccd1 vccd1 _17389_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_58_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09826_ _09826_/A _09826_/B vssd1 vssd1 vccd1 vccd1 _12016_/B sky130_fd_sc_hd__nor2_1
XFILLER_47_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout478 _15393_/A vssd1 vssd1 vccd1 vccd1 _10255_/A sky130_fd_sc_hd__buf_6
Xfanout489 _12275_/B vssd1 vssd1 vccd1 vccd1 _13051_/B sky130_fd_sc_hd__buf_2
XFILLER_100_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09757_ _09890_/A _09756_/Y _15538_/A _14863_/B vssd1 vssd1 vccd1 vccd1 _09898_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_100_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_47 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09688_ _09721_/A _09721_/B vssd1 vssd1 vccd1 vccd1 _09739_/A sky130_fd_sc_hd__nand2_1
XFILLER_55_874 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11650_ _11651_/A _15042_/B _15008_/B _11518_/A vssd1 vssd1 vccd1 vccd1 _11650_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_42_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_732 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10601_ _10601_/A _10601_/B vssd1 vssd1 vccd1 vccd1 _10603_/B sky130_fd_sc_hd__xnor2_1
X_11581_ _11538_/B _11551_/X _11579_/A _11614_/A vssd1 vssd1 vccd1 vccd1 _11582_/C
+ sky130_fd_sc_hd__o211ai_1
XFILLER_120_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_787 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10532_ _11122_/A _10851_/B _10647_/D _10532_/D vssd1 vssd1 vccd1 vccd1 _10535_/A
+ sky130_fd_sc_hd__and4_1
X_13320_ _13434_/B _13434_/D _13321_/D _14213_/A vssd1 vssd1 vccd1 vccd1 _13322_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_11_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13251_ _13121_/A _13123_/A _13249_/Y _13250_/X vssd1 vssd1 vccd1 vccd1 _13252_/A
+ sky130_fd_sc_hd__o211a_1
X_10463_ _10463_/A _10463_/B vssd1 vssd1 vccd1 vccd1 _10465_/B sky130_fd_sc_hd__nor2_1
XFILLER_6_447 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12202_ _12367_/B _12201_/B _12201_/C vssd1 vssd1 vccd1 vccd1 _12202_/Y sky130_fd_sc_hd__a21oi_2
X_13182_ _13182_/A _13948_/C _13182_/C vssd1 vssd1 vccd1 vccd1 _13184_/B sky130_fd_sc_hd__and3_1
XFILLER_164_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10394_ _10395_/A _10393_/Y _10719_/C _10525_/D vssd1 vssd1 vccd1 vccd1 _10505_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_163_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12133_ _11932_/A _12592_/C _11933_/A _11931_/B vssd1 vssd1 vccd1 vccd1 _12141_/A
+ sky130_fd_sc_hd__a31o_1
X_16941_ _16813_/Y _16986_/A _16940_/X _16994_/A vssd1 vssd1 vccd1 vccd1 _16943_/B
+ sky130_fd_sc_hd__o211a_1
X_12064_ _14356_/S _12063_/X _15457_/A vssd1 vssd1 vccd1 vccd1 _12064_/X sky130_fd_sc_hd__o21a_1
XFILLER_151_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_890 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11015_ _11016_/B _11016_/A vssd1 vssd1 vccd1 vccd1 _11015_/X sky130_fd_sc_hd__and2b_1
XFILLER_78_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16872_ _16872_/A _16872_/B _16871_/X vssd1 vssd1 vccd1 vccd1 _16872_/X sky130_fd_sc_hd__or3b_2
XFILLER_78_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15823_ _15821_/X _15823_/B vssd1 vssd1 vccd1 vccd1 _15825_/B sky130_fd_sc_hd__and2b_1
XFILLER_38_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15754_ _15666_/B _15853_/A _15753_/X vssd1 vssd1 vccd1 vccd1 _15756_/A sky130_fd_sc_hd__a21oi_1
X_12966_ _12966_/A _12966_/B vssd1 vssd1 vccd1 vccd1 _12968_/B sky130_fd_sc_hd__xnor2_1
XFILLER_46_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14705_ _14734_/A _14705_/B vssd1 vssd1 vccd1 vccd1 _14705_/Y sky130_fd_sc_hd__nand2_1
XTAP_3394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11917_ _08874_/A _08873_/X _11914_/X _11916_/A vssd1 vssd1 vccd1 vccd1 _11917_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15685_ _15686_/B _15685_/B _15587_/B vssd1 vssd1 vccd1 vccd1 _15782_/A sky130_fd_sc_hd__or3b_1
XTAP_2671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12897_ _12897_/A _12897_/B vssd1 vssd1 vccd1 vccd1 _12899_/C sky130_fd_sc_hd__xnor2_1
XTAP_2682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17424_ input59/X _17424_/A2 _17423_/X _17426_/C1 vssd1 vssd1 vccd1 vccd1 _17540_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_2693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14636_ _14636_/A _14636_/B vssd1 vssd1 vccd1 vccd1 _14636_/Y sky130_fd_sc_hd__nand2_1
X_11848_ _14636_/A _13625_/B vssd1 vssd1 vccd1 vccd1 _11848_/Y sky130_fd_sc_hd__nor2_2
XFILLER_60_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17355_ input57/X _17355_/B _17355_/C vssd1 vssd1 vccd1 vccd1 _17355_/X sky130_fd_sc_hd__or3_1
XFILLER_159_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14567_ _14567_/A _14567_/B vssd1 vssd1 vccd1 vccd1 _14569_/C sky130_fd_sc_hd__xnor2_1
X_11779_ _11778_/A _17138_/A _17138_/B _11777_/Y vssd1 vssd1 vccd1 vccd1 _11781_/B
+ sky130_fd_sc_hd__a31o_2
XFILLER_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16306_ _16579_/A _16399_/B _16306_/C vssd1 vssd1 vccd1 vccd1 _16310_/B sky130_fd_sc_hd__or3_1
XFILLER_146_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13518_ _12544_/X _12547_/X _13833_/S vssd1 vssd1 vccd1 vccd1 _13519_/B sky130_fd_sc_hd__mux2_1
XFILLER_119_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17286_ _17572_/Q _17289_/B vssd1 vssd1 vccd1 vccd1 _17286_/X sky130_fd_sc_hd__and2_1
X_14498_ _14562_/A _14498_/B vssd1 vssd1 vccd1 vccd1 _14501_/B sky130_fd_sc_hd__and2_1
XFILLER_174_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16237_ _16238_/A _16238_/B vssd1 vssd1 vccd1 vccd1 _16339_/B sky130_fd_sc_hd__nand2_1
XFILLER_146_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13449_ _13450_/B _13450_/C _14050_/D _14167_/A vssd1 vssd1 vccd1 vccd1 _13451_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16168_ _16168_/A _16938_/B _16168_/C vssd1 vssd1 vccd1 vccd1 _16170_/A sky130_fd_sc_hd__or3_1
XFILLER_126_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15119_ _15119_/A _15119_/B vssd1 vssd1 vccd1 vccd1 _15119_/Y sky130_fd_sc_hd__nor2_1
XFILLER_5_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08990_ _11922_/A _12127_/D vssd1 vssd1 vccd1 vccd1 _08991_/B sky130_fd_sc_hd__nand2_1
XFILLER_88_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16099_ _15994_/A _15994_/B _16100_/B _15991_/X vssd1 vssd1 vccd1 vccd1 _16099_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_134_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_903 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09611_ _09755_/A _09755_/B _10309_/B _10311_/D vssd1 vssd1 vccd1 vccd1 _09746_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_110_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09542_ _09484_/A _09484_/B _09484_/C vssd1 vssd1 vccd1 vccd1 _09628_/B sky130_fd_sc_hd__a21oi_1
XFILLER_83_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_991 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09473_ _09473_/A _09591_/A _09473_/C vssd1 vssd1 vccd1 vccd1 _09474_/B sky130_fd_sc_hd__or3_1
XFILLER_70_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_960 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_708 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout220 _15148_/Y vssd1 vssd1 vccd1 vccd1 _17083_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_114_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout231 _14930_/Y vssd1 vssd1 vccd1 vccd1 _15804_/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_87_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout242 _16869_/C1 vssd1 vssd1 vccd1 vccd1 _14944_/A sky130_fd_sc_hd__clkbuf_4
Xfanout253 _15998_/A vssd1 vssd1 vccd1 vccd1 _16207_/B sky130_fd_sc_hd__clkbuf_4
Xfanout264 _17295_/X vssd1 vssd1 vccd1 vccd1 _17429_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_115_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout275 _14939_/X vssd1 vssd1 vccd1 vccd1 _15373_/B sky130_fd_sc_hd__buf_2
Xfanout286 _12212_/S vssd1 vssd1 vccd1 vccd1 _17365_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_87_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09809_ _09919_/A _09919_/B vssd1 vssd1 vccd1 vccd1 _09920_/A sky130_fd_sc_hd__nand2_1
Xfanout297 _15130_/S vssd1 vssd1 vccd1 vccd1 _15103_/S sky130_fd_sc_hd__buf_2
XFILLER_101_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12820_ _12820_/A _12820_/B _12820_/C vssd1 vssd1 vccd1 vccd1 _12821_/B sky130_fd_sc_hd__and3_1
XFILLER_90_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12751_ _12751_/A _12910_/A vssd1 vssd1 vccd1 vccd1 _12754_/A sky130_fd_sc_hd__nor2_1
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11702_ _15793_/A _15793_/B vssd1 vssd1 vccd1 vccd1 _15888_/B sky130_fd_sc_hd__nand2_1
XFILLER_15_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15470_ _15442_/Y _15443_/X _15441_/X vssd1 vssd1 vccd1 vccd1 _15522_/A sky130_fd_sc_hd__a21o_1
X_12682_ _12682_/A _12682_/B vssd1 vssd1 vccd1 vccd1 _12685_/A sky130_fd_sc_hd__xnor2_1
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14421_ _12847_/B _12852_/X _14421_/S vssd1 vssd1 vccd1 vccd1 _14421_/X sky130_fd_sc_hd__mux2_1
X_11633_ _11649_/A _11632_/B _11632_/A vssd1 vssd1 vccd1 vccd1 _11635_/B sky130_fd_sc_hd__o21ba_1
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17140_ _17140_/A _17140_/B _17140_/C vssd1 vssd1 vccd1 vccd1 _17140_/X sky130_fd_sc_hd__or3_1
X_14352_ _14352_/A _14352_/B vssd1 vssd1 vccd1 vccd1 _14354_/B sky130_fd_sc_hd__or2_1
X_11564_ _11564_/A _11590_/A vssd1 vssd1 vccd1 vccd1 _11566_/B sky130_fd_sc_hd__nor2_1
XFILLER_11_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13303_ _13303_/A _13303_/B vssd1 vssd1 vccd1 vccd1 _13304_/B sky130_fd_sc_hd__xnor2_1
X_10515_ _10510_/X _10514_/X _10502_/X _10503_/Y vssd1 vssd1 vccd1 vccd1 _10517_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_128_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17071_ _11773_/A _11773_/B _17070_/Y vssd1 vssd1 vccd1 vccd1 _17077_/A sky130_fd_sc_hd__o21a_1
X_11495_ _11495_/A _11495_/B _11532_/A vssd1 vssd1 vccd1 vccd1 _11499_/A sky130_fd_sc_hd__nor3b_2
XFILLER_144_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14283_ _14284_/B _14283_/B vssd1 vssd1 vccd1 vccd1 _14283_/X sky130_fd_sc_hd__and2b_1
XFILLER_155_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16022_ _16226_/C _16165_/B _17119_/C _15726_/A vssd1 vssd1 vccd1 vccd1 _16022_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_109_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13234_ _13235_/B _13235_/A vssd1 vssd1 vccd1 vccd1 _13361_/B sky130_fd_sc_hd__and2b_1
X_10446_ _10560_/B _10446_/B _10446_/C vssd1 vssd1 vccd1 vccd1 _10685_/A sky130_fd_sc_hd__and3_1
XFILLER_136_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10377_ _15393_/A _10920_/B vssd1 vssd1 vccd1 vccd1 _10487_/A sky130_fd_sc_hd__nand2_1
X_13165_ _13165_/A _13165_/B _13165_/C vssd1 vssd1 vccd1 vccd1 _13178_/B sky130_fd_sc_hd__nand3_1
XFILLER_97_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12116_ _12116_/A _12116_/B vssd1 vssd1 vccd1 vccd1 _12118_/C sky130_fd_sc_hd__or2_1
XFILLER_124_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13096_ _12924_/A _12926_/B _12924_/B vssd1 vssd1 vccd1 vccd1 _13103_/A sky130_fd_sc_hd__o21ba_1
XFILLER_111_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12047_ _12040_/Y _12042_/Y _12044_/Y _12046_/Y _12383_/S _12865_/S vssd1 vssd1 vccd1
+ vccd1 _12047_/X sky130_fd_sc_hd__mux4_1
X_16924_ _13993_/B _16868_/A _16923_/Y vssd1 vssd1 vccd1 vccd1 _16924_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_66_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16855_ _16716_/Y _16854_/D _16854_/X _16852_/Y vssd1 vssd1 vccd1 vccd1 _16931_/B
+ sky130_fd_sc_hd__a211oi_4
XFILLER_120_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_32 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15806_ _15901_/S _15179_/X _15175_/A vssd1 vssd1 vccd1 vccd1 _15806_/Y sky130_fd_sc_hd__o21ai_1
X_16786_ _16786_/A _16786_/B vssd1 vssd1 vccd1 vccd1 _16853_/C sky130_fd_sc_hd__xor2_1
XFILLER_18_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13998_ _13998_/A _13998_/B vssd1 vssd1 vccd1 vccd1 _14001_/A sky130_fd_sc_hd__nor2_1
XFILLER_92_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15737_ _15737_/A _15737_/B vssd1 vssd1 vccd1 vccd1 _15740_/A sky130_fd_sc_hd__xnor2_1
XFILLER_18_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_90 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12949_ _12949_/A _13092_/A vssd1 vssd1 vccd1 vccd1 _12950_/C sky130_fd_sc_hd__and2_1
XFILLER_92_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15668_ _15668_/A _15668_/B vssd1 vssd1 vccd1 vccd1 _15671_/A sky130_fd_sc_hd__xor2_1
XFILLER_33_354 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17407_ _17407_/A _17425_/B vssd1 vssd1 vccd1 vccd1 _17407_/X sky130_fd_sc_hd__or2_1
X_14619_ _14658_/B _14619_/B vssd1 vssd1 vccd1 vccd1 _14621_/C sky130_fd_sc_hd__or2_1
XFILLER_21_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15599_ _15599_/A _15599_/B vssd1 vssd1 vccd1 vccd1 _15601_/B sky130_fd_sc_hd__nand2_1
XFILLER_159_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_1013 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17338_ _09319_/D _17360_/A2 _17337_/X _17406_/C1 vssd1 vssd1 vccd1 vccd1 _17498_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_146_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17269_ _17457_/Q _17290_/A2 _17267_/X _17268_/X _17293_/C1 vssd1 vssd1 vccd1 vccd1
+ _17457_/D sky130_fd_sc_hd__o221a_1
XFILLER_134_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_278 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_470 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08973_ _08973_/A _08973_/B _09095_/A vssd1 vssd1 vccd1 vccd1 _08974_/B sky130_fd_sc_hd__or3_1
XFILLER_114_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_608 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09525_ _09630_/A _09630_/B vssd1 vssd1 vccd1 vccd1 _09525_/X sky130_fd_sc_hd__and2_1
XFILLER_71_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09456_ _09456_/A _09456_/B vssd1 vssd1 vccd1 vccd1 _09543_/B sky130_fd_sc_hd__xnor2_1
XPHY_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09387_ _09387_/A _09387_/B _09387_/C vssd1 vssd1 vccd1 vccd1 _09388_/A sky130_fd_sc_hd__and3_1
XFILLER_40_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10300_ _10300_/A _10418_/A vssd1 vssd1 vccd1 vccd1 _10411_/A sky130_fd_sc_hd__or2_1
X_11280_ _11283_/B _11280_/B vssd1 vssd1 vccd1 vccd1 _11281_/C sky130_fd_sc_hd__nor2_1
XFILLER_152_215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10231_ _10134_/A _10134_/C _10134_/B vssd1 vssd1 vccd1 vccd1 _10231_/X sky130_fd_sc_hd__a21o_1
XFILLER_10_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10162_ _10162_/A _10170_/A _10162_/C vssd1 vssd1 vccd1 vccd1 _10163_/B sky130_fd_sc_hd__or3_1
XFILLER_160_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_34 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14970_ _14899_/X _14968_/X _11675_/B vssd1 vssd1 vccd1 vccd1 _16025_/A sky130_fd_sc_hd__a21o_2
X_10093_ _09806_/A _09807_/Y _10094_/A _10092_/X vssd1 vssd1 vccd1 vccd1 _10348_/A
+ sky130_fd_sc_hd__a211oi_1
XFILLER_48_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13921_ _13921_/A _13921_/B _13921_/C vssd1 vssd1 vccd1 vccd1 _13922_/B sky130_fd_sc_hd__nand3_1
XFILLER_74_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16640_ _11756_/A _11756_/B _16568_/B _16568_/A vssd1 vssd1 vccd1 vccd1 _16641_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_19_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13852_ _13852_/A _13852_/B _13853_/B vssd1 vssd1 vccd1 vccd1 _13958_/B sky130_fd_sc_hd__and3_1
XFILLER_16_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12803_ _12804_/B _13321_/D _13194_/D _12804_/A vssd1 vssd1 vccd1 vccd1 _12805_/A
+ sky130_fd_sc_hd__a22oi_1
X_16571_ _16571_/A _16571_/B _14774_/A vssd1 vssd1 vccd1 vccd1 _16572_/B sky130_fd_sc_hd__or3b_1
X_13783_ _13784_/A _13784_/B vssd1 vssd1 vccd1 vccd1 _13891_/A sky130_fd_sc_hd__nor2_1
X_10995_ _10995_/A _10995_/B vssd1 vssd1 vccd1 vccd1 _10996_/C sky130_fd_sc_hd__nor2_1
XFILLER_43_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1043 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15522_ _15522_/A _15522_/B vssd1 vssd1 vccd1 vccd1 _15523_/B sky130_fd_sc_hd__xor2_1
X_12734_ _13035_/A _12734_/B _13802_/B _13704_/B vssd1 vssd1 vccd1 vccd1 _12735_/B
+ sky130_fd_sc_hd__and4_1
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_994 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15453_ _15532_/A _15453_/B _15453_/C vssd1 vssd1 vccd1 vccd1 _15532_/B sky130_fd_sc_hd__nand3_1
X_12665_ _12665_/A _12665_/B vssd1 vssd1 vccd1 vccd1 _12668_/A sky130_fd_sc_hd__xor2_1
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14404_ _14399_/X _14466_/B _14296_/X _14404_/C1 vssd1 vssd1 vccd1 vccd1 _14405_/C
+ sky130_fd_sc_hd__a211o_1
X_11616_ _11617_/A _11617_/B _11617_/C vssd1 vssd1 vccd1 vccd1 _11616_/Y sky130_fd_sc_hd__nor3_1
XFILLER_168_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15384_ _15097_/X _15100_/Y _15384_/S vssd1 vssd1 vccd1 vccd1 _15384_/X sky130_fd_sc_hd__mux2_1
X_12596_ _12596_/A _12755_/A vssd1 vssd1 vccd1 vccd1 _12599_/A sky130_fd_sc_hd__nor2_1
XFILLER_168_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17123_ _17124_/A _17124_/B vssd1 vssd1 vccd1 vccd1 _17125_/A sky130_fd_sc_hd__nand2_1
XFILLER_7_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14335_ _14332_/X _14333_/Y _14239_/A _14256_/X vssd1 vssd1 vccd1 vccd1 _14337_/C
+ sky130_fd_sc_hd__a211oi_1
X_11547_ _11586_/A _11705_/A _11547_/C vssd1 vssd1 vccd1 vccd1 _15888_/A sky130_fd_sc_hd__nand3b_1
XFILLER_11_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17054_ _17090_/A _17093_/A vssd1 vssd1 vccd1 vccd1 _17055_/B sky130_fd_sc_hd__nand2_1
XFILLER_116_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14266_ _14266_/A _14266_/B vssd1 vssd1 vccd1 vccd1 _14268_/B sky130_fd_sc_hd__xnor2_1
X_11478_ _11520_/C _14850_/A _11440_/A _11438_/Y vssd1 vssd1 vccd1 vccd1 _11479_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_143_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16005_ _17119_/B _16005_/B _16005_/C vssd1 vssd1 vccd1 vccd1 _16007_/B sky130_fd_sc_hd__and3_1
X_13217_ _13903_/A _13968_/B _13216_/C vssd1 vssd1 vccd1 vccd1 _13218_/B sky130_fd_sc_hd__a21o_1
X_10429_ _10429_/A _10429_/B vssd1 vssd1 vccd1 vccd1 _10436_/A sky130_fd_sc_hd__nor2_1
X_14197_ _14197_/A _14197_/B _14197_/C vssd1 vssd1 vccd1 vccd1 _14198_/B sky130_fd_sc_hd__and3_1
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13148_ _13632_/A _13735_/B _14065_/B _14213_/C vssd1 vssd1 vccd1 vccd1 _13149_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_44_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13079_ _13450_/B _13080_/C _13080_/D _13080_/A vssd1 vssd1 vccd1 vccd1 _13083_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_111_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16907_ _16906_/A _16906_/B _16908_/A vssd1 vssd1 vccd1 vccd1 _17012_/A sky130_fd_sc_hd__a21o_1
XFILLER_111_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16838_ _16838_/A _16838_/B vssd1 vssd1 vccd1 vccd1 _16841_/A sky130_fd_sc_hd__xnor2_1
XFILLER_20_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16769_ _16770_/A _16770_/B _16770_/C vssd1 vssd1 vccd1 vccd1 _16771_/A sky130_fd_sc_hd__o21ai_1
XFILLER_19_693 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09310_ _09310_/A _09310_/B vssd1 vssd1 vccd1 vccd1 _09311_/C sky130_fd_sc_hd__xnor2_1
XFILLER_34_663 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09241_ _09242_/A _09242_/B _09242_/C vssd1 vssd1 vccd1 vccd1 _11990_/A sky130_fd_sc_hd__a21o_1
XFILLER_33_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09172_ _09172_/A _09172_/B vssd1 vssd1 vccd1 vccd1 _09502_/C sky130_fd_sc_hd__and2_1
XFILLER_135_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_749 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_911 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08956_ _09325_/B _12445_/D _11902_/B _09755_/A vssd1 vssd1 vccd1 vccd1 _08957_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_56_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08887_ _08887_/A _08887_/B vssd1 vssd1 vccd1 vccd1 _08888_/B sky130_fd_sc_hd__nor2_1
XFILLER_84_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09508_ _09508_/A _09508_/B vssd1 vssd1 vccd1 vccd1 _09630_/A sky130_fd_sc_hd__xor2_1
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10780_ _11749_/A _11749_/B vssd1 vssd1 vccd1 vccd1 _10780_/Y sky130_fd_sc_hd__nand2_1
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09439_ _09439_/A _09439_/B vssd1 vssd1 vccd1 vccd1 _09441_/C sky130_fd_sc_hd__or2_1
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12450_ _12451_/B _12451_/A vssd1 vssd1 vccd1 vccd1 _12450_/X sky130_fd_sc_hd__and2b_1
XFILLER_40_677 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11401_ _11349_/A _11349_/B _11349_/C vssd1 vssd1 vccd1 vccd1 _11402_/B sky130_fd_sc_hd__a21oi_1
X_12381_ _12696_/A _12379_/B _12380_/Y vssd1 vssd1 vccd1 vccd1 _12403_/A sky130_fd_sc_hd__a21o_1
XANTENNA_80 _16880_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_91 _10743_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14120_ _14279_/A _14120_/B vssd1 vssd1 vccd1 vccd1 _14278_/A sky130_fd_sc_hd__nand2b_1
X_11332_ _11281_/A _15617_/A _11281_/C vssd1 vssd1 vccd1 vccd1 _11333_/B sky130_fd_sc_hd__a21oi_1
XFILLER_126_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14051_ _14051_/A _14158_/A vssd1 vssd1 vccd1 vccd1 _14054_/A sky130_fd_sc_hd__or2_1
X_11263_ _11264_/A _11264_/C vssd1 vssd1 vccd1 vccd1 _11270_/B sky130_fd_sc_hd__nor2_1
XFILLER_141_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13002_ _13002_/A _13002_/B vssd1 vssd1 vccd1 vccd1 _13268_/A sky130_fd_sc_hd__or2_1
XFILLER_122_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10214_ _10214_/A _10214_/B _10214_/C vssd1 vssd1 vccd1 vccd1 _10215_/B sky130_fd_sc_hd__or3_1
X_11194_ _11194_/A _11194_/B vssd1 vssd1 vccd1 vccd1 _11195_/B sky130_fd_sc_hd__nor2_1
XFILLER_133_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10145_ _10145_/A _10145_/B vssd1 vssd1 vccd1 vccd1 _10268_/B sky130_fd_sc_hd__xnor2_1
XFILLER_43_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14953_ _17363_/A _10308_/B _10180_/C vssd1 vssd1 vccd1 vccd1 _15038_/B sky130_fd_sc_hd__a21o_1
X_10076_ _10208_/A _10208_/B vssd1 vssd1 vccd1 vccd1 _10209_/A sky130_fd_sc_hd__nor2_1
XFILLER_130_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13904_ _13904_/A _13904_/B vssd1 vssd1 vccd1 vccd1 _13906_/C sky130_fd_sc_hd__xnor2_1
XFILLER_48_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14884_ _14888_/B _14888_/C _14888_/D vssd1 vssd1 vccd1 vccd1 _14887_/B sky130_fd_sc_hd__or3_2
XFILLER_35_416 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16623_ _16699_/A _16623_/B vssd1 vssd1 vccd1 vccd1 _16623_/X sky130_fd_sc_hd__or2_1
XFILLER_75_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13835_ _14421_/S _11848_/Y _13834_/Y _13832_/Y _12853_/X vssd1 vssd1 vccd1 vccd1
+ _13835_/X sky130_fd_sc_hd__a32o_1
XFILLER_90_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16554_ _16554_/A _16554_/B vssd1 vssd1 vccd1 vccd1 _16557_/C sky130_fd_sc_hd__xnor2_1
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13766_ _14215_/A _13966_/D vssd1 vssd1 vccd1 vccd1 _13767_/B sky130_fd_sc_hd__nand2_1
XFILLER_15_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10978_ _10978_/A _10978_/B vssd1 vssd1 vccd1 vccd1 _11049_/C sky130_fd_sc_hd__xor2_1
XFILLER_16_674 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15505_ _15505_/A _15505_/B vssd1 vssd1 vccd1 vccd1 _15512_/A sky130_fd_sc_hd__xnor2_1
X_12717_ _12717_/A _12717_/B vssd1 vssd1 vccd1 vccd1 _12720_/A sky130_fd_sc_hd__xnor2_1
X_16485_ _16485_/A _16485_/B vssd1 vssd1 vccd1 vccd1 _16485_/Y sky130_fd_sc_hd__nand2_1
X_13697_ _13697_/A _13800_/A vssd1 vssd1 vccd1 vccd1 _13698_/C sky130_fd_sc_hd__and2_1
X_15436_ _15436_/A _15436_/B vssd1 vssd1 vccd1 vccd1 _15439_/A sky130_fd_sc_hd__xnor2_1
XFILLER_129_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12648_ _12795_/A _12942_/D _12496_/A _12494_/B vssd1 vssd1 vccd1 vccd1 _12649_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_169_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15367_ _15365_/X _15367_/B vssd1 vssd1 vccd1 vccd1 _15369_/A sky130_fd_sc_hd__nand2b_1
XFILLER_156_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12579_ _12579_/A _12579_/B vssd1 vssd1 vccd1 vccd1 _12581_/B sky130_fd_sc_hd__xnor2_1
XFILLER_50_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_502 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17106_ _11775_/Y _17105_/Y _16922_/A vssd1 vssd1 vccd1 vccd1 _17106_/Y sky130_fd_sc_hd__o21ai_1
X_14318_ _14318_/A _14318_/B _14385_/B _14433_/B vssd1 vssd1 vccd1 vccd1 _14389_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_171_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15298_ _15299_/A _15299_/B vssd1 vssd1 vccd1 vccd1 _15298_/Y sky130_fd_sc_hd__nor2_1
X_17037_ _17037_/A _17037_/B vssd1 vssd1 vccd1 vccd1 _17056_/B sky130_fd_sc_hd__nor2_1
X_14249_ _16723_/A _14383_/B _14248_/C vssd1 vssd1 vccd1 vccd1 _14250_/B sky130_fd_sc_hd__a21o_1
XFILLER_98_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout808 _12158_/D vssd1 vssd1 vccd1 vccd1 _09555_/C sky130_fd_sc_hd__buf_2
XFILLER_112_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout819 _09265_/C vssd1 vssd1 vccd1 vccd1 _15541_/A sky130_fd_sc_hd__buf_4
XFILLER_124_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08810_ _17395_/A _11861_/B _11859_/D _17397_/A vssd1 vssd1 vccd1 vccd1 _08812_/A
+ sky130_fd_sc_hd__a22oi_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09790_ _09933_/A _09790_/B vssd1 vssd1 vccd1 vccd1 _09919_/A sky130_fd_sc_hd__xnor2_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08741_ _17612_/Q _08743_/A _08740_/Y vssd1 vssd1 vccd1 vccd1 _17612_/D sky130_fd_sc_hd__a21o_1
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_906 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_522 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09224_ _17407_/A _09557_/B vssd1 vssd1 vccd1 vccd1 _09225_/B sky130_fd_sc_hd__nand2_1
XFILLER_148_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09155_ _09155_/A vssd1 vssd1 vccd1 vccd1 _09155_/Y sky130_fd_sc_hd__inv_2
XFILLER_147_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09086_ _09325_/B _11902_/B _09926_/B _17373_/A vssd1 vssd1 vccd1 vccd1 _09086_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_174_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_515 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_590 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_36 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09988_ _09988_/A _09988_/B vssd1 vssd1 vccd1 vccd1 _10106_/A sky130_fd_sc_hd__xnor2_1
XFILLER_107_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08939_ _09325_/B _09350_/B _11895_/C _17373_/A vssd1 vssd1 vccd1 vccd1 _08941_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_29_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11950_ _11947_/X _11948_/Y _09016_/A _09016_/Y vssd1 vssd1 vccd1 vccd1 _11998_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_85_872 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10901_ _10901_/A _10901_/B vssd1 vssd1 vccd1 vccd1 _10902_/C sky130_fd_sc_hd__nor2_1
XFILLER_123_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11881_ _17391_/A _17389_/A _12088_/D _12079_/B vssd1 vssd1 vccd1 vccd1 _11882_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_44_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13620_ _13729_/B _13621_/B vssd1 vssd1 vccd1 vccd1 _13620_/Y sky130_fd_sc_hd__nand2_1
X_10832_ _10863_/A vssd1 vssd1 vccd1 vccd1 _11075_/A sky130_fd_sc_hd__inv_2
XFILLER_26_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13551_ _13966_/A _14213_/B _13664_/D _13551_/D vssd1 vssd1 vccd1 vccd1 _13680_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_73_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10763_ _10771_/A _10734_/X _10760_/A _10761_/Y vssd1 vssd1 vccd1 vccd1 _10764_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_41_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12502_ _12804_/B _13067_/D _12923_/D _12804_/A vssd1 vssd1 vccd1 vccd1 _12504_/A
+ sky130_fd_sc_hd__a22oi_1
X_16270_ _16270_/A _16270_/B _16270_/C vssd1 vssd1 vccd1 vccd1 _16271_/B sky130_fd_sc_hd__nor3_1
XFILLER_41_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13482_ _13482_/A _13482_/B vssd1 vssd1 vccd1 vccd1 _13483_/B sky130_fd_sc_hd__or2_1
XFILLER_160_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10694_ _10694_/A _11027_/A _10954_/D _10905_/D vssd1 vssd1 vccd1 vccd1 _10694_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_139_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15221_ _15221_/A _15221_/B vssd1 vssd1 vccd1 vccd1 _15226_/A sky130_fd_sc_hd__xnor2_1
X_12433_ _12588_/A _12434_/B _12434_/C vssd1 vssd1 vccd1 vccd1 _12435_/A sky130_fd_sc_hd__a21o_1
XFILLER_32_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_384 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15152_ _16315_/D _15152_/B _15151_/B vssd1 vssd1 vccd1 vccd1 _15932_/A sky130_fd_sc_hd__or3b_4
XFILLER_153_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12364_ _12364_/A _12364_/B _12364_/C vssd1 vssd1 vccd1 vccd1 _12366_/A sky130_fd_sc_hd__and3_1
XFILLER_148_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14103_ _14104_/A _14104_/B vssd1 vssd1 vccd1 vccd1 _14192_/B sky130_fd_sc_hd__nand2_1
X_11315_ _11423_/B _11561_/D vssd1 vssd1 vccd1 vccd1 _11362_/A sky130_fd_sc_hd__nand2_1
XFILLER_99_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15083_ _15278_/A _16226_/B _15647_/A _15846_/A vssd1 vssd1 vccd1 vccd1 _15083_/X
+ sky130_fd_sc_hd__a22o_1
X_12295_ _12770_/A _12770_/B _12463_/D _12295_/D vssd1 vssd1 vccd1 vccd1 _12508_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_107_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14034_ _14122_/B _14034_/B vssd1 vssd1 vccd1 vccd1 _14034_/Y sky130_fd_sc_hd__nand2_1
X_11246_ _11246_/A _11246_/B vssd1 vssd1 vccd1 vccd1 _11308_/B sky130_fd_sc_hd__nor2_1
XFILLER_164_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11177_ _11015_/X _11019_/X _11175_/Y _11176_/X vssd1 vssd1 vccd1 vccd1 _11182_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_95_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10128_ _10128_/A _10128_/B vssd1 vssd1 vccd1 vccd1 _10251_/A sky130_fd_sc_hd__nor2_1
X_15985_ _15867_/B _15875_/B _15867_/A vssd1 vssd1 vccd1 vccd1 _15987_/B sky130_fd_sc_hd__a21bo_1
XFILLER_67_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10059_ _10059_/A _10059_/B _10059_/C vssd1 vssd1 vccd1 vccd1 _10086_/A sky130_fd_sc_hd__nor3_1
XFILLER_94_168 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14936_ _14942_/A _10062_/B _15248_/C _16799_/A2 _14935_/X vssd1 vssd1 vccd1 vccd1
+ _14944_/B sky130_fd_sc_hd__o32a_1
XFILLER_36_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14867_ _14867_/A _17065_/A _17029_/B vssd1 vssd1 vccd1 vccd1 _17139_/B sky130_fd_sc_hd__and3_1
XFILLER_24_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16606_ _16807_/A _16606_/B vssd1 vssd1 vccd1 vccd1 _16607_/B sky130_fd_sc_hd__nand2_1
XFILLER_17_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13818_ _13818_/A _13818_/B vssd1 vssd1 vccd1 vccd1 _13820_/B sky130_fd_sc_hd__nand2_1
X_17586_ fanout938/X _17586_/D vssd1 vssd1 vccd1 vccd1 _17586_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14798_ _14791_/X _14797_/X _11469_/X vssd1 vssd1 vccd1 vccd1 _14798_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_17_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_791 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16537_ _16537_/A _16537_/B vssd1 vssd1 vccd1 vccd1 _16541_/A sky130_fd_sc_hd__xnor2_1
XFILLER_50_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13749_ _13749_/A _13749_/B vssd1 vssd1 vccd1 vccd1 _13751_/B sky130_fd_sc_hd__nand2_1
XFILLER_92_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16468_ _16469_/A _16469_/B vssd1 vssd1 vccd1 vccd1 _16558_/A sky130_fd_sc_hd__and2b_1
XFILLER_148_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15419_ _15419_/A _15419_/B vssd1 vssd1 vccd1 vccd1 _15422_/A sky130_fd_sc_hd__xor2_1
XFILLER_164_619 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16399_ _16399_/A _16399_/B vssd1 vssd1 vccd1 vccd1 _16400_/C sky130_fd_sc_hd__nor2_1
XFILLER_157_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09911_ _09912_/A _09912_/B _09912_/C vssd1 vssd1 vccd1 vccd1 _09913_/A sky130_fd_sc_hd__o21ai_1
XFILLER_171_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout605 _12050_/S vssd1 vssd1 vccd1 vccd1 _11839_/S sky130_fd_sc_hd__buf_2
Xfanout616 _13948_/C vssd1 vssd1 vccd1 vccd1 _13852_/B sky130_fd_sc_hd__buf_2
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09842_ _09842_/A _09842_/B _09848_/B vssd1 vssd1 vccd1 vccd1 _09863_/B sky130_fd_sc_hd__or3_1
Xfanout627 _14383_/B vssd1 vssd1 vccd1 vccd1 _14708_/D sky130_fd_sc_hd__buf_2
XFILLER_140_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout638 _11815_/B vssd1 vssd1 vccd1 vccd1 _12439_/D sky130_fd_sc_hd__buf_2
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout649 _17506_/Q vssd1 vssd1 vccd1 vccd1 _14765_/B sky130_fd_sc_hd__buf_6
XFILLER_113_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09773_ _09773_/A _09773_/B _09773_/C vssd1 vssd1 vccd1 vccd1 _09813_/A sky130_fd_sc_hd__or3_1
XFILLER_100_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08724_ _17508_/Q vssd1 vssd1 vccd1 vccd1 _17134_/B sky130_fd_sc_hd__clkinv_2
XFILLER_160_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_1046 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09207_ _09208_/B _09208_/A vssd1 vssd1 vccd1 vccd1 _09211_/B sky130_fd_sc_hd__and2b_1
XFILLER_10_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09138_ _09170_/B _09170_/A vssd1 vssd1 vccd1 vccd1 _09138_/X sky130_fd_sc_hd__and2b_1
XFILLER_135_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09069_ _09069_/A _09076_/B vssd1 vssd1 vccd1 vccd1 _09071_/B sky130_fd_sc_hd__nand2_1
XFILLER_2_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11100_ _11100_/A _11100_/B vssd1 vssd1 vccd1 vccd1 _11238_/A sky130_fd_sc_hd__xnor2_1
XFILLER_123_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12080_ _12080_/A _12080_/B vssd1 vssd1 vccd1 vccd1 _12082_/B sky130_fd_sc_hd__xnor2_1
XFILLER_1_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11031_ _11032_/A _11032_/B vssd1 vssd1 vccd1 vccd1 _11176_/A sky130_fd_sc_hd__and2_1
XFILLER_89_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15770_ _15750_/A _16065_/B _15663_/A _15660_/X vssd1 vssd1 vccd1 vccd1 _15772_/C
+ sky130_fd_sc_hd__a31oi_1
XTAP_3510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12982_ _12983_/B _12982_/B vssd1 vssd1 vccd1 vccd1 _12984_/A sky130_fd_sc_hd__nand2b_1
XFILLER_91_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14721_ _14747_/B _14721_/B vssd1 vssd1 vccd1 vccd1 _14723_/C sky130_fd_sc_hd__and2_1
XTAP_3554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11933_ _11933_/A _11933_/B vssd1 vssd1 vccd1 vccd1 _11935_/B sky130_fd_sc_hd__xnor2_1
XFILLER_57_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_51 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17440_ fanout939/X _17440_/D vssd1 vssd1 vccd1 vccd1 _17440_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_72_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_577 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14652_ _14683_/A _14693_/A vssd1 vssd1 vccd1 vccd1 _14653_/B sky130_fd_sc_hd__nor2_1
XTAP_2864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11864_ _11865_/A _11865_/B vssd1 vssd1 vccd1 vccd1 _12085_/A sky130_fd_sc_hd__nand2_1
XFILLER_73_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13603_ _13603_/A _13603_/B _13603_/C vssd1 vssd1 vccd1 vccd1 _13604_/B sky130_fd_sc_hd__and3_1
X_10815_ _10816_/A _10816_/B vssd1 vssd1 vccd1 vccd1 _11057_/B sky130_fd_sc_hd__nand2_1
XTAP_2897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17371_ _17371_/A _17371_/B vssd1 vssd1 vccd1 vccd1 _17371_/Y sky130_fd_sc_hd__nand2_1
XFILLER_32_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14583_ _14583_/A _14583_/B _14583_/C vssd1 vssd1 vccd1 vccd1 _14584_/B sky130_fd_sc_hd__and3_1
X_11795_ _14775_/A _14776_/A _14777_/A _16209_/C vssd1 vssd1 vccd1 vccd1 _11799_/B
+ sky130_fd_sc_hd__or4_1
X_16322_ _16505_/A _16743_/C _17043_/B _15397_/A vssd1 vssd1 vccd1 vccd1 _16324_/A
+ sky130_fd_sc_hd__a22o_1
X_13534_ _13534_/A _13534_/B vssd1 vssd1 vccd1 vccd1 _13535_/B sky130_fd_sc_hd__xnor2_1
X_10746_ _10746_/A _10984_/A vssd1 vssd1 vccd1 vccd1 _11160_/A sky130_fd_sc_hd__or2_1
XFILLER_41_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16253_ _16254_/A _16254_/B vssd1 vssd1 vccd1 vccd1 _16347_/B sky130_fd_sc_hd__nor2_1
XFILLER_173_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13465_ _13465_/A _13465_/B vssd1 vssd1 vccd1 vccd1 _13485_/A sky130_fd_sc_hd__xor2_1
X_10677_ _10678_/A _10677_/B _10677_/C vssd1 vssd1 vccd1 vccd1 _10678_/B sky130_fd_sc_hd__nand3_1
X_15204_ _16935_/A _15204_/B _15270_/A vssd1 vssd1 vccd1 vccd1 _15205_/B sky130_fd_sc_hd__or3b_1
XFILLER_9_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12416_ _13028_/A _13348_/B vssd1 vssd1 vccd1 vccd1 _12417_/B sky130_fd_sc_hd__nand2_1
XFILLER_173_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16184_ _16184_/A _16184_/B vssd1 vssd1 vccd1 vccd1 _16192_/A sky130_fd_sc_hd__nor2_1
XFILLER_127_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13396_ _13632_/A _13735_/B _13632_/D _14065_/B vssd1 vssd1 vccd1 vccd1 _13526_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_154_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15135_ _15805_/A _15711_/B _15134_/X vssd1 vssd1 vccd1 vccd1 _15135_/Y sky130_fd_sc_hd__a21oi_1
X_12347_ _12180_/B _12182_/B _12180_/A vssd1 vssd1 vccd1 vccd1 _12349_/B sky130_fd_sc_hd__o21ba_1
XFILLER_126_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15066_ _16582_/A _15064_/X _15055_/X vssd1 vssd1 vccd1 vccd1 _15066_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_114_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12278_ _12278_/A _12278_/B vssd1 vssd1 vccd1 vccd1 _12281_/A sky130_fd_sc_hd__xnor2_1
XFILLER_4_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14017_ _14018_/A _14018_/B _14018_/C vssd1 vssd1 vccd1 vccd1 _14113_/A sky130_fd_sc_hd__a21o_1
XFILLER_141_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11229_ _11229_/A _11229_/B vssd1 vssd1 vccd1 vccd1 _11229_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_122_560 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_883 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15968_ _15969_/A _15969_/B vssd1 vssd1 vccd1 vccd1 _16084_/B sky130_fd_sc_hd__and2_1
XFILLER_64_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14919_ _14916_/X _14918_/Y _15103_/S vssd1 vssd1 vccd1 vccd1 _14919_/X sky130_fd_sc_hd__mux2_1
X_15899_ _15895_/B _16008_/A2 _16008_/B1 _15898_/A _14944_/A vssd1 vssd1 vccd1 vccd1
+ _15899_/X sky130_fd_sc_hd__a221o_1
XFILLER_64_875 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17569_ fanout934/X _17569_/D vssd1 vssd1 vccd1 vccd1 _17569_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_424 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout402 _12171_/A vssd1 vssd1 vccd1 vccd1 _10559_/A sky130_fd_sc_hd__clkbuf_4
Xfanout413 _13950_/A vssd1 vssd1 vccd1 vccd1 _13846_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_99_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout424 _14776_/A vssd1 vssd1 vccd1 vccd1 _12869_/A sky130_fd_sc_hd__buf_2
Xfanout435 _12077_/A vssd1 vssd1 vccd1 vccd1 _09414_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_59_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout446 _10242_/A1 vssd1 vssd1 vccd1 vccd1 _10241_/B sky130_fd_sc_hd__buf_2
XFILLER_24_1018 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout457 _17524_/Q vssd1 vssd1 vccd1 vccd1 _13035_/A sky130_fd_sc_hd__buf_2
X_09825_ _09825_/A _09825_/B vssd1 vssd1 vccd1 vccd1 _09826_/B sky130_fd_sc_hd__and2_1
Xfanout468 _17523_/Q vssd1 vssd1 vccd1 vccd1 _08791_/B sky130_fd_sc_hd__buf_2
XFILLER_171_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout479 _17522_/Q vssd1 vssd1 vccd1 vccd1 _15393_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_86_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09756_ _09755_/B _10311_/D _10308_/B _09755_/A vssd1 vssd1 vccd1 vccd1 _09756_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_55_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_55 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09687_ _09576_/A _09575_/C _09575_/B vssd1 vssd1 vccd1 vccd1 _09721_/B sky130_fd_sc_hd__a21o_1
XTAP_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_59 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10600_ _11027_/B _10805_/D _10593_/A _10592_/A vssd1 vssd1 vccd1 vccd1 _10603_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_168_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11580_ _11579_/A _11614_/A _11538_/B _11551_/X vssd1 vssd1 vccd1 vccd1 _11583_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_23_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10531_ _10531_/A _10536_/A _10531_/C vssd1 vssd1 vccd1 vccd1 _10540_/B sky130_fd_sc_hd__or3_1
XFILLER_168_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13250_ _13249_/A _13249_/B _13249_/C _13249_/D vssd1 vssd1 vccd1 vccd1 _13250_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_155_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10462_ _10454_/A _10455_/X _10463_/A _10461_/X vssd1 vssd1 vccd1 vccd1 _10463_/B
+ sky130_fd_sc_hd__a211oi_2
XFILLER_171_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12201_ _12367_/B _12201_/B _12201_/C vssd1 vssd1 vccd1 vccd1 _12371_/A sky130_fd_sc_hd__and3_1
XFILLER_170_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13181_ _13181_/A _13181_/B vssd1 vssd1 vccd1 vccd1 _13184_/A sky130_fd_sc_hd__nand2_1
XFILLER_108_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10393_ _10963_/B _10508_/D _10736_/D _10963_/A vssd1 vssd1 vccd1 vccd1 _10393_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_123_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12132_ _12343_/B _12132_/B vssd1 vssd1 vccd1 vccd1 _12145_/A sky130_fd_sc_hd__nor2_1
XFILLER_124_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16940_ _16317_/A _16165_/B _17119_/C _16809_/C vssd1 vssd1 vccd1 vccd1 _16940_/X
+ sky130_fd_sc_hd__a22o_1
X_12063_ _16011_/A _16011_/B _12063_/C vssd1 vssd1 vccd1 vccd1 _12063_/X sky130_fd_sc_hd__or3_2
XFILLER_77_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11014_ _10966_/A _10965_/B _10965_/A vssd1 vssd1 vccd1 vccd1 _11016_/B sky130_fd_sc_hd__o21ba_1
XFILLER_77_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16871_ _16735_/A _14481_/X _17164_/C _15460_/X vssd1 vssd1 vccd1 vccd1 _16871_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_65_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15822_ _16129_/A _16591_/B _15821_/C _15821_/D vssd1 vssd1 vccd1 vccd1 _15823_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_38_60 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15753_ _16446_/A _16416_/A _16619_/A _16410_/A vssd1 vssd1 vccd1 vccd1 _15753_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_18_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12965_ _16965_/C _13551_/D vssd1 vssd1 vccd1 vccd1 _12966_/B sky130_fd_sc_hd__nand2_1
XTAP_3351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11916_ _11916_/A vssd1 vssd1 vccd1 vccd1 _11916_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_363 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14704_ _13516_/X _13519_/B _14757_/S vssd1 vssd1 vccd1 vccd1 _14705_/B sky130_fd_sc_hd__mux2_1
XTAP_3384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15684_ _15580_/B _15582_/B _15580_/A vssd1 vssd1 vccd1 vccd1 _15686_/B sky130_fd_sc_hd__o21ba_1
XTAP_3395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12896_ _12897_/A _12897_/B vssd1 vssd1 vccd1 vccd1 _13057_/B sky130_fd_sc_hd__and2b_1
XFILLER_45_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17423_ _17423_/A _17425_/B vssd1 vssd1 vccd1 vccd1 _17423_/X sky130_fd_sc_hd__or2_1
X_14635_ _13273_/X _13276_/B _14757_/S vssd1 vssd1 vccd1 vccd1 _14636_/B sky130_fd_sc_hd__mux2_1
XTAP_2694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11847_ _12442_/A _14933_/A _14924_/C vssd1 vssd1 vccd1 vccd1 _13625_/B sky130_fd_sc_hd__or3_2
XTAP_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17354_ _12447_/B _17356_/A2 _17353_/X _17420_/C1 vssd1 vssd1 vccd1 vccd1 _17506_/D
+ sky130_fd_sc_hd__o211a_1
X_14566_ _14566_/A _14566_/B vssd1 vssd1 vccd1 vccd1 _14567_/B sky130_fd_sc_hd__nor2_1
XTAP_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11778_ _11778_/A _11778_/B vssd1 vssd1 vccd1 vccd1 _11778_/Y sky130_fd_sc_hd__nand2_1
XFILLER_159_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13517_ _12710_/A _13516_/X _16653_/A vssd1 vssd1 vccd1 vccd1 _13517_/Y sky130_fd_sc_hd__o21ai_1
X_16305_ _14778_/B _16115_/B _16298_/A vssd1 vssd1 vccd1 vccd1 _16306_/C sky130_fd_sc_hd__a21oi_1
X_10729_ _10729_/A _10729_/B vssd1 vssd1 vccd1 vccd1 _11212_/B sky130_fd_sc_hd__xor2_2
X_17285_ _17604_/Q _17291_/A2 _17291_/B1 vssd1 vssd1 vccd1 vccd1 _17285_/X sky130_fd_sc_hd__a21o_1
X_14497_ _14497_/A _14497_/B _14497_/C vssd1 vssd1 vccd1 vccd1 _14498_/B sky130_fd_sc_hd__or3_1
XFILLER_173_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16236_ _16416_/A _16499_/B vssd1 vssd1 vccd1 vccd1 _16238_/B sky130_fd_sc_hd__nor2_1
XFILLER_118_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13448_ _16723_/A _13691_/C vssd1 vssd1 vccd1 vccd1 _13459_/A sky130_fd_sc_hd__and2_2
XFILLER_174_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16167_ _16168_/A _16938_/B vssd1 vssd1 vccd1 vccd1 _16259_/C sky130_fd_sc_hd__nor2_1
XFILLER_86_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13379_ _13252_/Y _13256_/A _13500_/B _13378_/X vssd1 vssd1 vccd1 vccd1 _13504_/A
+ sky130_fd_sc_hd__a211oi_2
XFILLER_86_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15118_ _15042_/X _15043_/X _15041_/X vssd1 vssd1 vccd1 vccd1 _15119_/B sky130_fd_sc_hd__a21boi_1
XFILLER_47_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16098_ _16098_/A vssd1 vssd1 vccd1 vccd1 _16100_/B sky130_fd_sc_hd__inv_2
XFILLER_88_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15049_ _16731_/B1 _15110_/B _15046_/Y _15048_/Y vssd1 vssd1 vccd1 vccd1 _15049_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_123_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09610_ _09610_/A _09614_/A _09610_/C vssd1 vssd1 vccd1 vccd1 _09618_/B sky130_fd_sc_hd__or3_1
XFILLER_68_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09541_ _09530_/B _09530_/C _09528_/Y _09485_/X vssd1 vssd1 vccd1 vccd1 _09541_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_83_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09472_ _09602_/A _09471_/Y _15538_/A _09926_/B vssd1 vssd1 vccd1 vccd1 _09610_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_51_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_279 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_8 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout210 _17362_/C vssd1 vssd1 vccd1 vccd1 _17321_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_59_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout221 _17156_/B vssd1 vssd1 vccd1 vccd1 _16111_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_59_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout243 _14871_/Y vssd1 vssd1 vccd1 vccd1 _16869_/C1 sky130_fd_sc_hd__clkbuf_4
Xfanout254 _11784_/X vssd1 vssd1 vccd1 vccd1 _15998_/A sky130_fd_sc_hd__buf_4
Xfanout265 _15147_/Y vssd1 vssd1 vccd1 vccd1 _16315_/D sky130_fd_sc_hd__buf_2
XFILLER_115_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout276 _17063_/A vssd1 vssd1 vccd1 vccd1 _08743_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_47_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout287 _15096_/S vssd1 vssd1 vccd1 vccd1 _14948_/A sky130_fd_sc_hd__clkbuf_4
X_09808_ _09808_/A _09808_/B vssd1 vssd1 vccd1 vccd1 _09919_/B sky130_fd_sc_hd__xnor2_1
Xfanout298 fanout299/X vssd1 vssd1 vccd1 vccd1 _15130_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_46_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09739_ _09739_/A _09739_/B vssd1 vssd1 vccd1 vccd1 _09740_/C sky130_fd_sc_hd__xnor2_1
XFILLER_15_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12750_ _13182_/A _13051_/B _13037_/B _13035_/C vssd1 vssd1 vccd1 vccd1 _12910_/A
+ sky130_fd_sc_hd__and4_1
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11701_ _11700_/B _11700_/C _11700_/A vssd1 vssd1 vccd1 vccd1 _15793_/B sky130_fd_sc_hd__a21bo_1
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12681_ _12682_/A _12682_/B vssd1 vssd1 vccd1 vccd1 _12681_/Y sky130_fd_sc_hd__nor2_1
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14420_ _14763_/S _14418_/X _14419_/Y _14358_/Y vssd1 vssd1 vccd1 vccd1 _17597_/D
+ sky130_fd_sc_hd__a31o_1
X_11632_ _11632_/A _11632_/B vssd1 vssd1 vccd1 vccd1 _11649_/B sky130_fd_sc_hd__or2_1
XFILLER_42_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14351_ _14349_/X _14351_/B vssd1 vssd1 vccd1 vccd1 _14416_/B sky130_fd_sc_hd__and2b_1
X_11563_ _11564_/A _11562_/Y _11630_/A _11563_/D vssd1 vssd1 vccd1 vccd1 _11590_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_155_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13302_ _13302_/A _13852_/B vssd1 vssd1 vccd1 vccd1 _13303_/B sky130_fd_sc_hd__nand2_1
X_10514_ _10613_/A _10613_/B vssd1 vssd1 vccd1 vccd1 _10514_/X sky130_fd_sc_hd__and2_1
X_17070_ _17105_/B _17070_/B vssd1 vssd1 vccd1 vccd1 _17070_/Y sky130_fd_sc_hd__nor2_1
XFILLER_128_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_223 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14282_ wire116/X _14281_/Y _14280_/X vssd1 vssd1 vccd1 vccd1 _14284_/B sky130_fd_sc_hd__o21ai_1
X_11494_ _11453_/B _11449_/B _11449_/C vssd1 vssd1 vccd1 vccd1 _11495_/B sky130_fd_sc_hd__a21oi_1
XFILLER_171_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16021_ _16021_/A _16021_/B vssd1 vssd1 vccd1 vccd1 _16595_/B sky130_fd_sc_hd__nand2_1
XFILLER_10_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13233_ _13099_/A _13101_/B _13099_/B vssd1 vssd1 vccd1 vccd1 _13235_/B sky130_fd_sc_hd__o21ba_1
X_10445_ _10445_/A _10445_/B vssd1 vssd1 vccd1 vccd1 _10446_/C sky130_fd_sc_hd__nor2_1
XFILLER_170_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_94 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13164_ _13178_/A vssd1 vssd1 vccd1 vccd1 _13312_/A sky130_fd_sc_hd__inv_2
XFILLER_108_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10376_ _10954_/A _11006_/B _10799_/B _14788_/B vssd1 vssd1 vccd1 vccd1 _10379_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_123_143 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12115_ _12115_/A _12115_/B vssd1 vssd1 vccd1 vccd1 _12116_/B sky130_fd_sc_hd__nor2_1
XFILLER_97_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_528 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13095_ _13095_/A _13095_/B vssd1 vssd1 vccd1 vccd1 _13114_/A sky130_fd_sc_hd__xnor2_1
XFILLER_123_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16923_ _13993_/B _16868_/A _17140_/A vssd1 vssd1 vccd1 vccd1 _16923_/Y sky130_fd_sc_hd__a21oi_1
X_12046_ _12046_/A _12046_/B vssd1 vssd1 vccd1 vccd1 _12046_/Y sky130_fd_sc_hd__nand2_1
X_16854_ _16566_/A _16566_/B _16854_/C _16854_/D vssd1 vssd1 vccd1 vccd1 _16854_/X
+ sky130_fd_sc_hd__and4bb_1
XFILLER_37_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15805_ _15805_/A _15805_/B vssd1 vssd1 vccd1 vccd1 _15805_/Y sky130_fd_sc_hd__nor2_1
XFILLER_19_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16785_ _16850_/A _16785_/B vssd1 vssd1 vccd1 vccd1 _16786_/B sky130_fd_sc_hd__or2_1
X_13997_ _13997_/A _13997_/B vssd1 vssd1 vccd1 vccd1 _13998_/B sky130_fd_sc_hd__and2_1
XFILLER_80_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15736_ _16136_/B _16152_/A vssd1 vssd1 vccd1 vccd1 _15737_/B sky130_fd_sc_hd__nand2_1
XFILLER_19_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12948_ _12947_/A _12947_/B _12947_/C vssd1 vssd1 vccd1 vccd1 _13092_/A sky130_fd_sc_hd__o21ai_1
XFILLER_80_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15667_ _16536_/A _16505_/A vssd1 vssd1 vccd1 vccd1 _15668_/B sky130_fd_sc_hd__nand2_1
X_12879_ _13643_/A _13704_/B vssd1 vssd1 vccd1 vccd1 _12881_/B sky130_fd_sc_hd__nand2_1
XTAP_2480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17406_ input49/X _17422_/A2 _17405_/X _17406_/C1 vssd1 vssd1 vccd1 vccd1 _17531_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_60_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14618_ _14618_/A _14618_/B vssd1 vssd1 vccd1 vccd1 _14619_/B sky130_fd_sc_hd__nor2_1
X_15598_ _15598_/A _15598_/B vssd1 vssd1 vccd1 vccd1 _15599_/B sky130_fd_sc_hd__nand2_1
XTAP_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17337_ input48/X _17353_/B _17353_/C vssd1 vssd1 vccd1 vccd1 _17337_/X sky130_fd_sc_hd__or3_1
XFILLER_53_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14549_ _14549_/A _14601_/B vssd1 vssd1 vccd1 vccd1 _14570_/A sky130_fd_sc_hd__nor2_1
XFILLER_140_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_596 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17268_ _17566_/Q _17289_/B vssd1 vssd1 vccd1 vccd1 _17268_/X sky130_fd_sc_hd__and2_1
XFILLER_101_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16219_ _16219_/A1 _13839_/X _17164_/C _14961_/X vssd1 vssd1 vccd1 vccd1 _16219_/Y
+ sky130_fd_sc_hd__o22ai_1
X_17199_ _17543_/Q _17199_/B vssd1 vssd1 vccd1 vccd1 _17199_/X sky130_fd_sc_hd__and2_1
XFILLER_127_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08972_ _08973_/B _09095_/A _08973_/A vssd1 vssd1 vccd1 vccd1 _09242_/A sky130_fd_sc_hd__o21ai_1
XFILLER_114_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09524_ _09524_/A _09524_/B vssd1 vssd1 vccd1 vccd1 _09630_/B sky130_fd_sc_hd__xnor2_1
XFILLER_52_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09455_ _09455_/A _09455_/B vssd1 vssd1 vccd1 vccd1 _09543_/A sky130_fd_sc_hd__nand2_1
XFILLER_101_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09386_ _09386_/A _09386_/B vssd1 vssd1 vccd1 vccd1 _09387_/C sky130_fd_sc_hd__xnor2_1
XFILLER_61_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_227 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10230_ _10157_/C _10157_/B _10155_/Y vssd1 vssd1 vccd1 vccd1 _10230_/X sky130_fd_sc_hd__a21bo_1
XFILLER_105_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10161_ _10054_/B _10159_/Y _10155_/A _10137_/X vssd1 vssd1 vccd1 vccd1 _10161_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10092_ _10091_/A _10091_/B _10091_/C vssd1 vssd1 vccd1 vccd1 _10092_/X sky130_fd_sc_hd__o21a_1
XFILLER_86_46 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13920_ _13921_/A _13921_/B _13921_/C vssd1 vssd1 vccd1 vccd1 _13922_/A sky130_fd_sc_hd__a21o_1
XFILLER_48_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13851_ _13851_/A _13958_/A vssd1 vssd1 vccd1 vccd1 _13853_/B sky130_fd_sc_hd__nor2_1
XFILLER_19_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12802_ _12619_/A _12621_/B _12619_/B vssd1 vssd1 vccd1 vccd1 _12809_/A sky130_fd_sc_hd__o21ba_1
XFILLER_62_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13782_ _13681_/B _13683_/B _13681_/A vssd1 vssd1 vccd1 vccd1 _13784_/B sky130_fd_sc_hd__o21ba_1
X_16570_ _14774_/A _16644_/B _16571_/A vssd1 vssd1 vccd1 vccd1 _16572_/A sky130_fd_sc_hd__a21bo_1
X_10994_ _10545_/C _10993_/D _11164_/A _10992_/Y vssd1 vssd1 vccd1 vccd1 _10996_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_27_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12733_ _12734_/B _13802_/B _13704_/B _13035_/A vssd1 vssd1 vccd1 vccd1 _12735_/A
+ sky130_fd_sc_hd__a22oi_1
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15521_ _15519_/X _15521_/B vssd1 vssd1 vccd1 vccd1 _15522_/B sky130_fd_sc_hd__nand2b_1
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15452_ _15532_/A _15453_/B _15453_/C vssd1 vssd1 vccd1 vccd1 _15454_/B sky130_fd_sc_hd__a21o_1
X_12664_ _12504_/A _12506_/B _12504_/B vssd1 vssd1 vccd1 vccd1 _12665_/B sky130_fd_sc_hd__o21ba_1
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14403_ _14424_/A vssd1 vssd1 vccd1 vccd1 _14405_/B sky130_fd_sc_hd__inv_2
X_11615_ _11614_/A _11614_/B _11614_/C vssd1 vssd1 vccd1 vccd1 _11617_/C sky130_fd_sc_hd__a21oi_1
XFILLER_168_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15383_ _10799_/Y _17163_/A2 _15382_/X _16977_/A vssd1 vssd1 vccd1 vccd1 _15383_/X
+ sky130_fd_sc_hd__o211a_1
X_12595_ _13182_/A _13051_/B _13035_/C _13908_/B vssd1 vssd1 vccd1 vccd1 _12755_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_168_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17122_ _17091_/A _17118_/A _17089_/A vssd1 vssd1 vccd1 vccd1 _17124_/B sky130_fd_sc_hd__a21o_1
X_14334_ _14239_/A _14256_/X _14332_/X _14333_/Y vssd1 vssd1 vccd1 vccd1 _14405_/A
+ sky130_fd_sc_hd__o211a_1
X_11546_ _11461_/B _11544_/Y _11543_/A _11502_/B vssd1 vssd1 vccd1 vccd1 _11547_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_7_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17053_ _17091_/A _17053_/B vssd1 vssd1 vccd1 vccd1 _17093_/B sky130_fd_sc_hd__nand2b_1
X_14265_ _14265_/A _14265_/B _14266_/B vssd1 vssd1 vccd1 vccd1 _14344_/A sky130_fd_sc_hd__and3_1
XFILLER_116_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11477_ _11477_/A _11514_/A _11477_/C vssd1 vssd1 vccd1 vccd1 _11487_/A sky130_fd_sc_hd__and3_1
X_16004_ _16004_/A _16004_/B vssd1 vssd1 vccd1 vccd1 _16004_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_125_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13216_ _13903_/A _13968_/B _13216_/C vssd1 vssd1 vccd1 vccd1 _13346_/B sky130_fd_sc_hd__nand3_1
XFILLER_125_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10428_ _14958_/A _10311_/D _10312_/A _10310_/Y vssd1 vssd1 vccd1 vccd1 _10429_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_14196_ _14197_/A _14197_/B _14197_/C vssd1 vssd1 vccd1 vccd1 _14276_/A sky130_fd_sc_hd__a21oi_1
XFILLER_98_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13147_ _13735_/B _14065_/B _14213_/C _13632_/A vssd1 vssd1 vccd1 vccd1 _13149_/A
+ sky130_fd_sc_hd__a22oi_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10359_ _11027_/B _10359_/B vssd1 vssd1 vccd1 vccd1 _10364_/A sky130_fd_sc_hd__nand2_1
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13078_ _12979_/A _12978_/B _12978_/A vssd1 vssd1 vccd1 vccd1 _13120_/A sky130_fd_sc_hd__a21bo_1
XFILLER_140_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16906_ _16906_/A _16906_/B vssd1 vssd1 vccd1 vccd1 _16908_/B sky130_fd_sc_hd__nand2_1
X_12029_ _12700_/C _14911_/B vssd1 vssd1 vccd1 vccd1 _12035_/C sky130_fd_sc_hd__nand2_1
XFILLER_38_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16837_ _16762_/A _16762_/B _16765_/A vssd1 vssd1 vccd1 vccd1 _16838_/B sky130_fd_sc_hd__a21o_1
XFILLER_66_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16768_ _16768_/A _16835_/B vssd1 vssd1 vccd1 vccd1 _16770_/C sky130_fd_sc_hd__nor2_1
X_15719_ _16917_/A _15705_/Y _15706_/X _15718_/X vssd1 vssd1 vccd1 vccd1 _15719_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_80_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16699_ _16699_/A _16699_/B vssd1 vssd1 vccd1 vccd1 _16701_/B sky130_fd_sc_hd__xnor2_1
XFILLER_61_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09240_ _09240_/A _09240_/B vssd1 vssd1 vccd1 vccd1 _09242_/C sky130_fd_sc_hd__xnor2_1
XFILLER_34_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09171_ _09178_/A _09178_/B _09178_/C vssd1 vssd1 vccd1 vccd1 _09179_/A sky130_fd_sc_hd__a21oi_2
XFILLER_159_360 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_780 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_923 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08955_ _08958_/A vssd1 vssd1 vccd1 vccd1 _08957_/C sky130_fd_sc_hd__inv_2
XFILLER_130_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_499 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08886_ _17397_/A _17395_/A _11859_/D _09030_/C vssd1 vssd1 vccd1 vccd1 _08887_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_56_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_726 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09507_ _09508_/A _09508_/B vssd1 vssd1 vccd1 vccd1 _09507_/Y sky130_fd_sc_hd__nor2_1
XFILLER_24_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09438_ _09438_/A _09438_/B vssd1 vssd1 vccd1 vccd1 _09439_/B sky130_fd_sc_hd__nor2_1
XFILLER_12_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09369_ _09370_/B _09370_/C _09370_/A vssd1 vssd1 vccd1 vccd1 _09387_/A sky130_fd_sc_hd__a21o_1
XFILLER_8_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11400_ _11403_/B _11400_/B _11400_/C vssd1 vssd1 vccd1 vccd1 _11451_/A sky130_fd_sc_hd__and3_1
XFILLER_138_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12380_ _16922_/A _12380_/B vssd1 vssd1 vccd1 vccd1 _12380_/Y sky130_fd_sc_hd__nand2_1
XANTENNA_70 _15151_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_81 _17496_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11331_ _11331_/A _11331_/B _11331_/C vssd1 vssd1 vccd1 vccd1 _11341_/B sky130_fd_sc_hd__nand3_1
XFILLER_126_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_30 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_92 _10743_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14050_ _14213_/A _14050_/B _14141_/D _14050_/D vssd1 vssd1 vccd1 vccd1 _14158_/A
+ sky130_fd_sc_hd__and4_1
X_11262_ _11124_/C _14851_/A _11125_/A _11123_/Y vssd1 vssd1 vccd1 vccd1 _11264_/C
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_107_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13001_ _13001_/A _13001_/B _13001_/C vssd1 vssd1 vccd1 vccd1 _13002_/B sky130_fd_sc_hd__and3_1
X_10213_ _10194_/A _10194_/B _10194_/C vssd1 vssd1 vccd1 vccd1 _10214_/C sky130_fd_sc_hd__o21a_1
XFILLER_106_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11193_ _11222_/B _11191_/X _11067_/Y _11069_/X vssd1 vssd1 vccd1 vccd1 _11194_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_133_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_807 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10144_ _10271_/A _10146_/B vssd1 vssd1 vccd1 vccd1 _10268_/A sky130_fd_sc_hd__nand2_1
XFILLER_48_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10075_ _10075_/A _10075_/B vssd1 vssd1 vccd1 vccd1 _10208_/B sky130_fd_sc_hd__nand2_1
X_14952_ _14952_/A _14952_/B vssd1 vssd1 vccd1 vccd1 _14952_/Y sky130_fd_sc_hd__nor2_1
XFILLER_153_84 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13903_ _13903_/A _14301_/C vssd1 vssd1 vccd1 vccd1 _13904_/B sky130_fd_sc_hd__nand2_1
XFILLER_36_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14883_ _15262_/B _15472_/A _15071_/A vssd1 vssd1 vccd1 vccd1 _14888_/D sky130_fd_sc_hd__or3b_1
X_16622_ _16622_/A _16622_/B _16622_/C vssd1 vssd1 vccd1 vccd1 _16623_/B sky130_fd_sc_hd__nor3_1
XFILLER_35_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13834_ _13834_/A vssd1 vssd1 vccd1 vccd1 _13834_/Y sky130_fd_sc_hd__inv_2
XFILLER_90_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16553_ _16554_/A _16554_/B vssd1 vssd1 vccd1 vccd1 _16636_/B sky130_fd_sc_hd__nand2b_1
X_13765_ _13765_/A _13765_/B vssd1 vssd1 vccd1 vccd1 _13767_/A sky130_fd_sc_hd__nor2_1
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10977_ _10978_/A _10978_/B vssd1 vssd1 vccd1 vccd1 _10977_/X sky130_fd_sc_hd__or2_1
XFILLER_16_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15504_ _15504_/A _15504_/B vssd1 vssd1 vccd1 vccd1 _15505_/B sky130_fd_sc_hd__xor2_1
XFILLER_16_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12716_ _12871_/A _13450_/C vssd1 vssd1 vccd1 vccd1 _12717_/B sky130_fd_sc_hd__nand2_1
XFILLER_71_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13696_ _13695_/A _13695_/B _13695_/C vssd1 vssd1 vccd1 vccd1 _13800_/A sky130_fd_sc_hd__o21ai_1
X_16484_ _12560_/A _14775_/X _14816_/X vssd1 vssd1 vccd1 vccd1 _16485_/B sky130_fd_sc_hd__a21o_1
X_12647_ _12798_/B _12647_/B vssd1 vssd1 vccd1 vccd1 _12650_/B sky130_fd_sc_hd__nand2_1
X_15435_ _15436_/A _15436_/B vssd1 vssd1 vccd1 vccd1 _15520_/A sky130_fd_sc_hd__and2_1
XFILLER_62_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1003 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15366_ _15365_/B _15366_/B vssd1 vssd1 vccd1 vccd1 _15367_/B sky130_fd_sc_hd__nand2b_1
X_12578_ _13302_/A _13802_/B vssd1 vssd1 vccd1 vccd1 _12579_/B sky130_fd_sc_hd__nand2_1
XFILLER_11_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17105_ _17105_/A _17105_/B vssd1 vssd1 vccd1 vccd1 _17105_/Y sky130_fd_sc_hd__nor2_1
X_11529_ _11529_/A _11529_/B vssd1 vssd1 vccd1 vccd1 _11530_/C sky130_fd_sc_hd__xnor2_1
XFILLER_171_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14317_ _14318_/B _14385_/B _14433_/B _14318_/A vssd1 vssd1 vccd1 vccd1 _14319_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_129_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15297_ _15228_/A _15228_/B _15231_/A vssd1 vssd1 vccd1 vccd1 _15299_/B sky130_fd_sc_hd__o21a_1
XFILLER_7_87 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14248_ _14772_/A _14383_/B _14248_/C vssd1 vssd1 vccd1 vccd1 _14330_/B sky130_fd_sc_hd__nand3_1
X_17036_ _17028_/A _17170_/B1 _17035_/X vssd1 vssd1 vccd1 vccd1 _17570_/D sky130_fd_sc_hd__a21oi_1
XFILLER_125_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14179_ _14180_/A _14180_/B vssd1 vssd1 vccd1 vccd1 _14273_/A sky130_fd_sc_hd__nand2b_1
XFILLER_98_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout809 _11281_/B vssd1 vssd1 vccd1 vccd1 _12158_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_98_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_967 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08740_ _08743_/A _14933_/A vssd1 vssd1 vccd1 vccd1 _08740_/Y sky130_fd_sc_hd__nor2_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_940 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09223_ _09223_/A _09223_/B vssd1 vssd1 vccd1 vccd1 _09225_/A sky130_fd_sc_hd__nor2_1
XFILLER_22_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09154_ _09131_/X _09138_/X _09152_/A _09153_/X vssd1 vssd1 vccd1 vccd1 _09155_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_148_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09085_ _17373_/A _09325_/B _11902_/B _09926_/B vssd1 vssd1 vccd1 vccd1 _09317_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_162_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_8 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_818 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09987_ _10244_/A _10920_/B vssd1 vssd1 vccd1 vccd1 _09988_/B sky130_fd_sc_hd__nand2_1
XFILLER_153_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08938_ _08923_/A _08922_/A _08922_/B vssd1 vssd1 vccd1 vccd1 _08945_/A sky130_fd_sc_hd__o21ba_1
XFILLER_76_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08869_ _08869_/A _08869_/B _08869_/C vssd1 vssd1 vccd1 vccd1 _08869_/Y sky130_fd_sc_hd__nand3_1
XFILLER_123_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10900_ _10993_/C _10899_/D _10995_/A _10898_/Y vssd1 vssd1 vccd1 vccd1 _10902_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_17_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11880_ _17389_/A _12088_/D _12079_/B _17391_/A vssd1 vssd1 vccd1 vccd1 _11882_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_83_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10831_ _11072_/B _11072_/C _11072_/A vssd1 vssd1 vccd1 vccd1 _10863_/A sky130_fd_sc_hd__a21o_1
XFILLER_26_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13550_ _14213_/B _13664_/D _13551_/D _13966_/A vssd1 vssd1 vccd1 vccd1 _13552_/A
+ sky130_fd_sc_hd__a22oi_1
X_10762_ _10760_/A _10761_/Y _10771_/A _10734_/X vssd1 vssd1 vccd1 vccd1 _10771_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_16_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_606 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12501_ _12501_/A _12501_/B vssd1 vssd1 vccd1 vccd1 _12518_/A sky130_fd_sc_hd__xnor2_1
XFILLER_73_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13481_ _13482_/A _13482_/B vssd1 vssd1 vccd1 vccd1 _13603_/A sky130_fd_sc_hd__nand2_1
XFILLER_40_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10693_ _10632_/B _10632_/C _10632_/D _10632_/A vssd1 vssd1 vccd1 vccd1 _10693_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_13_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15220_ _15220_/A _15220_/B vssd1 vssd1 vccd1 vccd1 _15221_/B sky130_fd_sc_hd__xnor2_1
X_12432_ _12432_/A _12432_/B vssd1 vssd1 vccd1 vccd1 _12434_/C sky130_fd_sc_hd__xnor2_1
XFILLER_138_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15151_ _15152_/B _15151_/B _16054_/B vssd1 vssd1 vccd1 vccd1 _15151_/X sky130_fd_sc_hd__and3b_1
X_12363_ _12190_/A _12189_/A _12189_/B _12191_/X vssd1 vssd1 vccd1 vccd1 _12364_/C
+ sky130_fd_sc_hd__a31o_1
XFILLER_138_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14102_ _14194_/A _14102_/B vssd1 vssd1 vccd1 vccd1 _14104_/B sky130_fd_sc_hd__xnor2_1
X_11314_ _11370_/A _15373_/C _11592_/B _17467_/D vssd1 vssd1 vccd1 vccd1 _11314_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_4_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15082_ _15278_/A _16226_/B _15342_/A vssd1 vssd1 vccd1 vccd1 _15164_/B sky130_fd_sc_hd__and3_1
XFILLER_153_355 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12294_ _12770_/B _12463_/D _12295_/D _17425_/A vssd1 vssd1 vccd1 vccd1 _12296_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_5_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14033_ _14122_/B _14034_/B vssd1 vssd1 vccd1 vccd1 _14033_/X sky130_fd_sc_hd__or2_1
X_11245_ _11117_/C _11117_/D _11118_/A _11116_/Y vssd1 vssd1 vccd1 vccd1 _11246_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_4_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11176_ _11176_/A _11176_/B _11176_/C vssd1 vssd1 vccd1 vccd1 _11176_/X sky130_fd_sc_hd__or3_1
XFILLER_79_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10127_ _10126_/B _10255_/B _10920_/B _10254_/A vssd1 vssd1 vccd1 vccd1 _10128_/B
+ sky130_fd_sc_hd__a22oi_1
XFILLER_110_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15984_ _15984_/A _15984_/B vssd1 vssd1 vccd1 vccd1 _15987_/A sky130_fd_sc_hd__xnor2_1
XFILLER_48_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10058_ _10057_/B _10057_/C _10057_/A vssd1 vssd1 vccd1 vccd1 _10059_/C sky130_fd_sc_hd__a21boi_1
X_14935_ _10062_/B _15108_/A _15248_/C _14934_/X vssd1 vssd1 vccd1 vccd1 _14935_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_91_810 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14866_ _17028_/A _17028_/B vssd1 vssd1 vccd1 vccd1 _17029_/B sky130_fd_sc_hd__and2_1
XFILLER_17_940 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16605_ _16827_/B _16681_/C _16514_/C _16603_/X vssd1 vssd1 vccd1 vccd1 _16607_/A
+ sky130_fd_sc_hd__o31a_1
X_13817_ _13817_/A _13817_/B vssd1 vssd1 vccd1 vccd1 _13820_/A sky130_fd_sc_hd__xnor2_1
XFILLER_90_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17585_ fanout939/X _17585_/D vssd1 vssd1 vccd1 vccd1 _17585_/Q sky130_fd_sc_hd__dfxtp_1
X_14797_ _14796_/B _14796_/C _14796_/D _11595_/B vssd1 vssd1 vccd1 vccd1 _14797_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_51_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16536_ _16536_/A _16695_/B _16537_/A vssd1 vssd1 vccd1 vccd1 _16622_/B sky130_fd_sc_hd__and3_1
X_13748_ _13748_/A _13748_/B vssd1 vssd1 vccd1 vccd1 _13751_/A sky130_fd_sc_hd__xnor2_1
XFILLER_149_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16467_ _16369_/A _16369_/B _16371_/Y vssd1 vssd1 vccd1 vccd1 _16469_/B sky130_fd_sc_hd__a21bo_1
X_13679_ _13680_/A _13680_/B _13680_/C vssd1 vssd1 vccd1 vccd1 _13681_/A sky130_fd_sc_hd__o21a_1
XFILLER_85_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15418_ _15501_/A _15418_/B _15419_/B vssd1 vssd1 vccd1 vccd1 _15501_/B sky130_fd_sc_hd__and3b_1
XFILLER_129_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16398_ _16398_/A _16398_/B vssd1 vssd1 vccd1 vccd1 _16398_/X sky130_fd_sc_hd__xor2_1
XFILLER_117_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15349_ _15350_/A _15350_/B vssd1 vssd1 vccd1 vccd1 _15426_/A sky130_fd_sc_hd__nor2_1
XFILLER_156_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17019_ _17028_/A _17153_/B _14766_/A vssd1 vssd1 vccd1 vccd1 _17066_/A sky130_fd_sc_hd__or3b_1
X_09910_ _09910_/A _09910_/B vssd1 vssd1 vccd1 vccd1 _09912_/C sky130_fd_sc_hd__nor2_1
XFILLER_99_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout606 _15058_/S0 vssd1 vssd1 vccd1 vccd1 _12050_/S sky130_fd_sc_hd__buf_2
XFILLER_99_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout617 _08967_/B vssd1 vssd1 vccd1 vccd1 _13948_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_59_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09841_ _09841_/A _09983_/A vssd1 vssd1 vccd1 vccd1 _09848_/B sky130_fd_sc_hd__nor2_1
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout628 _14829_/B vssd1 vssd1 vccd1 vccd1 _14383_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_86_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout639 _15033_/A3 vssd1 vssd1 vccd1 vccd1 _11815_/B sky130_fd_sc_hd__clkbuf_4
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_328 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09772_ _09773_/C _09812_/A vssd1 vssd1 vccd1 vccd1 _09772_/X sky130_fd_sc_hd__and2b_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08723_ _11651_/A vssd1 vssd1 vccd1 vccd1 _08723_/Y sky130_fd_sc_hd__inv_2
XFILLER_85_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09206_ _09206_/A _09375_/A vssd1 vssd1 vccd1 vccd1 _09208_/B sky130_fd_sc_hd__nor2_1
XFILLER_167_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09137_ _09167_/A _09137_/B vssd1 vssd1 vccd1 vccd1 _09170_/B sky130_fd_sc_hd__xnor2_1
XFILLER_135_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09068_ _09062_/X _09294_/A _09076_/A _09055_/Y vssd1 vssd1 vccd1 vccd1 _09076_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_162_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11030_ _11030_/A _11030_/B vssd1 vssd1 vccd1 vccd1 _11032_/B sky130_fd_sc_hd__xnor2_1
XFILLER_2_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12981_ _12981_/A _12981_/B vssd1 vssd1 vccd1 vccd1 _12983_/B sky130_fd_sc_hd__xnor2_1
XFILLER_64_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14720_ _14719_/A _14719_/B _14719_/C vssd1 vssd1 vccd1 vccd1 _14721_/B sky130_fd_sc_hd__o21ai_1
XTAP_3544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11932_ _11932_/A _11932_/B vssd1 vssd1 vccd1 vccd1 _11933_/B sky130_fd_sc_hd__nand2_1
XFILLER_17_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_876 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11863_ _12070_/A _11859_/D _08748_/A _08747_/A vssd1 vssd1 vccd1 vccd1 _11865_/B
+ sky130_fd_sc_hd__a31o_1
X_14651_ _14710_/C _14651_/B vssd1 vssd1 vccd1 vccd1 _14693_/B sky130_fd_sc_hd__xnor2_2
XTAP_3599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10814_ _10814_/A _10814_/B vssd1 vssd1 vccd1 vccd1 _10816_/B sky130_fd_sc_hd__xnor2_1
XTAP_2887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13602_ _13603_/A _13603_/B _13603_/C vssd1 vssd1 vccd1 vccd1 _13604_/A sky130_fd_sc_hd__a21oi_1
XTAP_2898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17370_ input61/X _17371_/B _17369_/Y _17378_/C1 vssd1 vssd1 vccd1 vccd1 _17513_/D
+ sky130_fd_sc_hd__o211a_1
X_14582_ _14582_/A vssd1 vssd1 vccd1 vccd1 _14584_/A sky130_fd_sc_hd__inv_2
X_11794_ _13689_/A _16723_/A _16644_/C _14774_/A vssd1 vssd1 vccd1 vccd1 _11798_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_158_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16321_ _16321_/A _16321_/B vssd1 vssd1 vccd1 vccd1 _16328_/A sky130_fd_sc_hd__xor2_1
XFILLER_43_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10745_ _10746_/A _10744_/Y _10745_/C _10745_/D vssd1 vssd1 vccd1 vccd1 _10984_/A
+ sky130_fd_sc_hd__and4bb_1
X_13533_ _13643_/A _13844_/C vssd1 vssd1 vccd1 vccd1 _13534_/B sky130_fd_sc_hd__nand2_1
XFILLER_40_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16252_ _16252_/A _16252_/B vssd1 vssd1 vccd1 vccd1 _16254_/B sky130_fd_sc_hd__xnor2_1
XFILLER_9_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13464_ _13578_/A _13464_/B vssd1 vssd1 vccd1 vccd1 _13465_/B sky130_fd_sc_hd__nand2_1
X_10676_ _10556_/B _10587_/Y _10667_/A _10667_/Y vssd1 vssd1 vccd1 vccd1 _10677_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_173_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15203_ _14877_/Y _14967_/D _08731_/A vssd1 vssd1 vccd1 vccd1 _15203_/X sky130_fd_sc_hd__a21o_1
X_12415_ _12415_/A _12415_/B vssd1 vssd1 vccd1 vccd1 _12417_/A sky130_fd_sc_hd__nor2_1
X_16183_ _16183_/A _16183_/B _16183_/C vssd1 vssd1 vccd1 vccd1 _16184_/B sky130_fd_sc_hd__nor3_1
X_13395_ _13735_/B _13632_/D _14065_/B _13632_/A vssd1 vssd1 vccd1 vccd1 _13398_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_166_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_867 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12346_ _12346_/A _12346_/B vssd1 vssd1 vccd1 vccd1 _12349_/A sky130_fd_sc_hd__xor2_1
X_15134_ _15116_/A _15131_/A _15130_/X _10419_/B vssd1 vssd1 vccd1 vccd1 _15134_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_126_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_388 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15065_ _14963_/X _15040_/X _15044_/Y _15045_/X vssd1 vssd1 vccd1 vccd1 _15065_/Y
+ sky130_fd_sc_hd__o22ai_1
X_12277_ _12907_/A _12445_/C vssd1 vssd1 vccd1 vccd1 _12278_/B sky130_fd_sc_hd__nand2_1
XFILLER_107_580 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14016_ _14016_/A _14016_/B vssd1 vssd1 vccd1 vccd1 _14018_/C sky130_fd_sc_hd__xor2_1
X_11228_ _11228_/A _11228_/B vssd1 vssd1 vccd1 vccd1 _11229_/B sky130_fd_sc_hd__xor2_1
XFILLER_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11159_ _11159_/A _11159_/B vssd1 vssd1 vccd1 vccd1 _11190_/A sky130_fd_sc_hd__xnor2_1
XFILLER_49_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15967_ _16084_/A _15967_/B vssd1 vssd1 vccd1 vccd1 _15969_/B sky130_fd_sc_hd__nor2_1
XFILLER_67_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14918_ _15102_/A _14918_/B vssd1 vssd1 vccd1 vccd1 _14918_/Y sky130_fd_sc_hd__nand2_1
XFILLER_64_843 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15898_ _15898_/A _15898_/B vssd1 vssd1 vccd1 vccd1 _15898_/Y sky130_fd_sc_hd__nor2_1
XFILLER_91_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14849_ _14849_/A _15314_/B vssd1 vssd1 vccd1 vccd1 _15381_/B sky130_fd_sc_hd__and2_1
XFILLER_23_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17568_ fanout940/X _17568_/D vssd1 vssd1 vccd1 vccd1 _17568_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16519_ _16519_/A _16519_/B _16519_/C vssd1 vssd1 vccd1 vccd1 _16520_/B sky130_fd_sc_hd__and3_1
XFILLER_20_902 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17499_ fanout946/X _17499_/D vssd1 vssd1 vccd1 vccd1 _17499_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_143_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_804 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout403 _17531_/Q vssd1 vssd1 vccd1 vccd1 _12171_/A sky130_fd_sc_hd__buf_2
XFILLER_87_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout414 _12871_/A vssd1 vssd1 vccd1 vccd1 _13950_/A sky130_fd_sc_hd__buf_2
Xfanout425 _17528_/Q vssd1 vssd1 vccd1 vccd1 _14776_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_113_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout436 _17527_/Q vssd1 vssd1 vccd1 vccd1 _12077_/A sky130_fd_sc_hd__buf_4
XFILLER_150_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_637 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout447 _17526_/Q vssd1 vssd1 vccd1 vccd1 _10242_/A1 sky130_fd_sc_hd__buf_4
X_09824_ _09825_/A _09825_/B vssd1 vssd1 vccd1 vccd1 _09826_/A sky130_fd_sc_hd__nor2_1
Xfanout458 _08791_/A vssd1 vssd1 vccd1 vccd1 _17391_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_101_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout469 _11790_/A vssd1 vssd1 vccd1 vccd1 _16809_/A sky130_fd_sc_hd__buf_4
XFILLER_150_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09755_ _09755_/A _09755_/B _10311_/D _10308_/B vssd1 vssd1 vccd1 vccd1 _09890_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_86_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_523 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09686_ _09686_/A _09686_/B vssd1 vssd1 vccd1 vccd1 _09768_/A sky130_fd_sc_hd__xnor2_1
XTAP_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_386 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10530_ _10531_/A _10531_/C vssd1 vssd1 vccd1 vccd1 _10536_/B sky130_fd_sc_hd__nor2_1
XFILLER_149_970 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10461_ _10336_/Y _10353_/X _10459_/A _10459_/Y vssd1 vssd1 vccd1 vccd1 _10461_/X
+ sky130_fd_sc_hd__o211a_1
X_12200_ _12200_/A _12200_/B vssd1 vssd1 vccd1 vccd1 _12201_/C sky130_fd_sc_hd__or2_1
XFILLER_89_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13180_ _13177_/Y _13312_/B _13046_/A _13047_/B vssd1 vssd1 vccd1 vccd1 _13189_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_164_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10392_ _10963_/A _10963_/B _10508_/D _10736_/D vssd1 vssd1 vccd1 vccd1 _10395_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_151_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12131_ _12131_/A _12131_/B vssd1 vssd1 vccd1 vccd1 _12132_/B sky130_fd_sc_hd__and2_1
XFILLER_108_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12062_ _12397_/B _12061_/Y _12383_/S vssd1 vssd1 vccd1 vccd1 _12063_/C sky130_fd_sc_hd__mux2_1
XFILLER_96_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_166 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11013_ _11013_/A _11013_/B vssd1 vssd1 vccd1 vccd1 _11016_/A sky130_fd_sc_hd__nor2_1
X_16870_ _14770_/A _14864_/A _17075_/A2 _16869_/X vssd1 vssd1 vccd1 vccd1 _16872_/B
+ sky130_fd_sc_hd__a31o_1
X_15821_ _16129_/A _16591_/B _15821_/C _15821_/D vssd1 vssd1 vccd1 vccd1 _15821_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_49_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15752_ _16416_/A _16619_/A vssd1 vssd1 vccd1 vccd1 _15853_/A sky130_fd_sc_hd__nor2_2
XTAP_3341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12964_ _12964_/A _12964_/B vssd1 vssd1 vccd1 vccd1 _12966_/A sky130_fd_sc_hd__nor2_1
XTAP_3352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14703_ _14756_/A1 _14700_/Y _14702_/Y _14667_/Y _14668_/X vssd1 vssd1 vccd1 vccd1
+ _17603_/D sky130_fd_sc_hd__a32o_1
XTAP_3374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11915_ _11915_/A _11915_/B _12148_/B _11913_/X vssd1 vssd1 vccd1 vccd1 _11916_/A
+ sky130_fd_sc_hd__or4bb_1
XFILLER_18_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15683_ _15769_/B _15682_/B _15682_/C vssd1 vssd1 vccd1 vccd1 _15690_/B sky130_fd_sc_hd__o21a_1
XTAP_3396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12895_ _12895_/A _12895_/B vssd1 vssd1 vccd1 vccd1 _12897_/B sky130_fd_sc_hd__xnor2_1
XFILLER_45_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17422_ input57/X _17422_/A2 _17421_/X _17422_/C1 vssd1 vssd1 vccd1 vccd1 _17539_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_2673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14634_ _14756_/A1 _14632_/X _14638_/B _14590_/Y _14591_/X vssd1 vssd1 vccd1 vccd1
+ _17601_/D sky130_fd_sc_hd__a32o_1
XTAP_2684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11846_ _12442_/A _14933_/A _14924_/C vssd1 vssd1 vccd1 vccd1 _13626_/B sky130_fd_sc_hd__nor3_2
XTAP_2695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17353_ input56/X _17353_/B _17353_/C vssd1 vssd1 vccd1 vccd1 _17353_/X sky130_fd_sc_hd__or3_1
XTAP_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11777_ _10098_/A _11778_/B _11778_/A vssd1 vssd1 vccd1 vccd1 _11777_/Y sky130_fd_sc_hd__a21boi_1
X_14565_ _14565_/A _14565_/B vssd1 vssd1 vccd1 vccd1 _14566_/B sky130_fd_sc_hd__nor2_1
XTAP_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16304_ _16304_/A _16304_/B _16304_/C vssd1 vssd1 vccd1 vccd1 _16310_/A sky130_fd_sc_hd__or3_1
X_10728_ _10728_/A _10728_/B vssd1 vssd1 vccd1 vccd1 _11212_/A sky130_fd_sc_hd__nand2_1
X_13516_ _12543_/X _12552_/B _13516_/S vssd1 vssd1 vccd1 vccd1 _13516_/X sky130_fd_sc_hd__mux2_2
XFILLER_13_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17284_ _17462_/Q _17293_/A2 _17282_/X _17283_/X _17284_/C1 vssd1 vssd1 vccd1 vccd1
+ _17462_/D sky130_fd_sc_hd__o221a_1
X_14496_ _14497_/A _14497_/B _14497_/C vssd1 vssd1 vccd1 vccd1 _14562_/A sky130_fd_sc_hd__o21ai_1
X_16235_ _16235_/A _16339_/A vssd1 vssd1 vccd1 vccd1 _16238_/A sky130_fd_sc_hd__and2_1
XFILLER_146_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13447_ _13444_/A _13445_/Y _13329_/A _13330_/B vssd1 vssd1 vccd1 vccd1 _13490_/B
+ sky130_fd_sc_hd__o211a_1
X_10659_ _10660_/A _10658_/Y _10993_/C _12054_/B vssd1 vssd1 vccd1 vccd1 _10757_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_173_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_642 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16166_ _15746_/X _16164_/Y _16279_/A vssd1 vssd1 vccd1 vccd1 _16175_/A sky130_fd_sc_hd__a21oi_1
XFILLER_126_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13378_ _13500_/A _13376_/X _13246_/A _13249_/C vssd1 vssd1 vccd1 vccd1 _13378_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_114_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15117_ _15117_/A _15117_/B vssd1 vssd1 vccd1 vccd1 _15119_/A sky130_fd_sc_hd__nand2_1
X_12329_ _12795_/A _12328_/B _12328_/C vssd1 vssd1 vccd1 vccd1 _12330_/B sky130_fd_sc_hd__a21o_1
XFILLER_115_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16097_ _16096_/A _16096_/B _16096_/C vssd1 vssd1 vccd1 vccd1 _16098_/A sky130_fd_sc_hd__o21ai_2
XFILLER_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15048_ _14796_/B _16008_/A2 _15047_/X _14944_/A vssd1 vssd1 vccd1 vccd1 _15048_/Y
+ sky130_fd_sc_hd__a211oi_1
XFILLER_114_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16999_ _17000_/A _17000_/B vssd1 vssd1 vccd1 vccd1 _17052_/B sky130_fd_sc_hd__and2_1
XFILLER_68_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09540_ _09540_/A _09540_/B vssd1 vssd1 vccd1 vccd1 _09674_/A sky130_fd_sc_hd__nor2_1
XFILLER_49_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09471_ _09755_/B _10180_/B _10309_/B _12471_/A vssd1 vssd1 vccd1 vccd1 _09471_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_52_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_776 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_759 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_634 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout200 _11853_/Y vssd1 vssd1 vccd1 vccd1 _15457_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_132_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout211 _17355_/B vssd1 vssd1 vccd1 vccd1 _17353_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_132_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout222 _14938_/X vssd1 vssd1 vccd1 vccd1 _17156_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_8_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout233 _16799_/A2 vssd1 vssd1 vccd1 vccd1 _17162_/A2 sky130_fd_sc_hd__clkbuf_4
Xfanout244 _16731_/B1 vssd1 vssd1 vccd1 vccd1 _17140_/A sky130_fd_sc_hd__buf_2
XFILLER_113_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout255 _14756_/A1 vssd1 vssd1 vccd1 vccd1 _14763_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_8_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout266 fanout266/A vssd1 vssd1 vccd1 vccd1 _17038_/C sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout277 _15523_/A vssd1 vssd1 vccd1 vccd1 _17063_/A sky130_fd_sc_hd__clkbuf_4
X_09807_ _09808_/A _09808_/B vssd1 vssd1 vccd1 vccd1 _09807_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_86_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout288 _12383_/S vssd1 vssd1 vccd1 vccd1 _15096_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_115_77 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout299 _08721_/Y vssd1 vssd1 vccd1 vccd1 fanout299/X sky130_fd_sc_hd__clkbuf_2
XFILLER_86_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09738_ _09732_/X _09868_/A _09724_/X _09725_/Y vssd1 vssd1 vccd1 vccd1 _09740_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_74_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09669_ _09668_/A _09668_/Y _09530_/X _09541_/X vssd1 vssd1 vccd1 vccd1 _09674_/B
+ sky130_fd_sc_hd__a211oi_2
XFILLER_43_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11700_ _11700_/A _11700_/B _11700_/C vssd1 vssd1 vccd1 vccd1 _11700_/Y sky130_fd_sc_hd__nand3_1
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12680_ _12522_/B _12522_/C _12522_/A vssd1 vssd1 vccd1 vccd1 _12682_/B sky130_fd_sc_hd__o21ba_1
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11631_ _11629_/B _15116_/B _11629_/D _11629_/A vssd1 vssd1 vccd1 vccd1 _11632_/B
+ sky130_fd_sc_hd__a22oi_1
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11562_ _11629_/B _11561_/C _11561_/D _11561_/A vssd1 vssd1 vccd1 vccd1 _11562_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_24_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14350_ _14350_/A _14350_/B _14350_/C vssd1 vssd1 vccd1 vccd1 _14351_/B sky130_fd_sc_hd__or3_1
XFILLER_156_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10513_ _10513_/A _10513_/B vssd1 vssd1 vccd1 vccd1 _10613_/B sky130_fd_sc_hd__nor2_1
X_13301_ _13301_/A _13301_/B vssd1 vssd1 vccd1 vccd1 _13303_/A sky130_fd_sc_hd__nor2_1
XFILLER_10_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14281_ _14281_/A _14281_/B vssd1 vssd1 vccd1 vccd1 _14281_/Y sky130_fd_sc_hd__nand2_1
X_11493_ _11496_/B _11493_/B _11493_/C vssd1 vssd1 vccd1 vccd1 _11532_/A sky130_fd_sc_hd__and3_1
XFILLER_155_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16020_ _16021_/A _16054_/B vssd1 vssd1 vccd1 vccd1 _17119_/C sky130_fd_sc_hd__and2_2
XFILLER_137_962 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13232_ _13232_/A _13232_/B vssd1 vssd1 vccd1 vccd1 _13235_/A sky130_fd_sc_hd__xnor2_1
X_10444_ _10321_/B _15003_/B _09502_/B _10321_/A vssd1 vssd1 vccd1 vccd1 _10445_/B
+ sky130_fd_sc_hd__a22oi_1
XFILLER_109_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13163_ _13165_/A _13165_/B _13165_/C vssd1 vssd1 vccd1 vccd1 _13178_/A sky130_fd_sc_hd__a21o_1
XFILLER_123_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10375_ _10390_/A _10375_/B vssd1 vssd1 vccd1 vccd1 _10382_/A sky130_fd_sc_hd__and2_1
XFILLER_124_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12114_ _12115_/A _12115_/B vssd1 vssd1 vccd1 vccd1 _12116_/A sky130_fd_sc_hd__and2_1
XFILLER_123_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13094_ _13578_/A _13968_/B vssd1 vssd1 vccd1 vccd1 _13095_/B sky130_fd_sc_hd__nand2_1
XFILLER_123_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_732 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16922_ _16922_/A _16922_/B vssd1 vssd1 vccd1 vccd1 _16922_/Y sky130_fd_sc_hd__nand2_1
XFILLER_105_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12045_ _12054_/A _15624_/A _11387_/C vssd1 vssd1 vccd1 vccd1 _12046_/B sky130_fd_sc_hd__a21o_1
XFILLER_104_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16853_ _16853_/A _16853_/B _16853_/C vssd1 vssd1 vccd1 vccd1 _16854_/D sky130_fd_sc_hd__and3_1
XFILLER_65_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15804_ _16809_/B _15804_/A2 _15803_/X vssd1 vssd1 vccd1 vccd1 _15804_/Y sky130_fd_sc_hd__a21oi_1
X_16784_ _16784_/A _16784_/B _16784_/C vssd1 vssd1 vccd1 vccd1 _16785_/B sky130_fd_sc_hd__and3_1
XFILLER_18_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13996_ _13997_/A _13997_/B vssd1 vssd1 vccd1 vccd1 _13998_/A sky130_fd_sc_hd__nor2_1
XTAP_3160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15735_ _15735_/A _15735_/B vssd1 vssd1 vccd1 vccd1 _15737_/A sky130_fd_sc_hd__nand2_1
XFILLER_34_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12947_ _12947_/A _12947_/B _12947_/C vssd1 vssd1 vccd1 vccd1 _12949_/A sky130_fd_sc_hd__or3_1
XFILLER_92_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15666_ _15666_/A _15666_/B vssd1 vssd1 vccd1 vccd1 _15668_/A sky130_fd_sc_hd__xnor2_1
XTAP_2470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12878_ _12878_/A _13040_/A vssd1 vssd1 vccd1 vccd1 _12881_/A sky130_fd_sc_hd__or2_1
XTAP_2481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17405_ _17405_/A _17421_/B vssd1 vssd1 vccd1 vccd1 _17405_/X sky130_fd_sc_hd__or2_1
XTAP_2492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14617_ _14618_/A _14618_/B vssd1 vssd1 vccd1 vccd1 _14658_/B sky130_fd_sc_hd__and2_1
X_11829_ _11837_/A _11829_/B vssd1 vssd1 vccd1 vccd1 _11829_/Y sky130_fd_sc_hd__nand2_1
XTAP_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15597_ _15598_/A _15598_/B vssd1 vssd1 vccd1 vccd1 _15599_/A sky130_fd_sc_hd__or2_1
XFILLER_60_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17336_ _09058_/C _17360_/A2 _17335_/X _17406_/C1 vssd1 vssd1 vccd1 vccd1 _17497_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_60_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_80 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14548_ _14548_/A _14601_/A _14548_/C vssd1 vssd1 vccd1 vccd1 _14601_/B sky130_fd_sc_hd__nor3_1
XFILLER_174_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17267_ _17598_/Q _17291_/A2 _17291_/B1 vssd1 vssd1 vccd1 vccd1 _17267_/X sky130_fd_sc_hd__a21o_1
XFILLER_128_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14479_ _14479_/A _14479_/B vssd1 vssd1 vccd1 vccd1 _14479_/Y sky130_fd_sc_hd__nand2_1
XFILLER_128_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16218_ _14778_/X _16799_/A2 _16799_/B1 _14778_/B _16869_/C1 vssd1 vssd1 vccd1 vccd1
+ _16218_/X sky130_fd_sc_hd__a221o_1
XFILLER_174_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17198_ input25/X input28/X _17198_/C _17428_/C vssd1 vssd1 vccd1 vccd1 _17199_/B
+ sky130_fd_sc_hd__and4b_2
X_16149_ _16667_/A _16681_/A _16827_/B _16416_/A vssd1 vssd1 vccd1 vccd1 _16149_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_127_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08971_ _08993_/C _08973_/B _08971_/C vssd1 vssd1 vccd1 vccd1 _09095_/A sky130_fd_sc_hd__nor3_1
XFILLER_114_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_448 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09523_ _09523_/A _09523_/B vssd1 vssd1 vccd1 vccd1 _09524_/B sky130_fd_sc_hd__nor2_1
XFILLER_37_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09454_ _09448_/X _09579_/A _09440_/X _09441_/Y vssd1 vssd1 vccd1 vccd1 _09455_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_51_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09385_ _09385_/A _09385_/B vssd1 vssd1 vccd1 vccd1 _09386_/B sky130_fd_sc_hd__xnor2_1
XFILLER_101_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10160_ _10137_/X _10155_/A _10159_/Y _10054_/B vssd1 vssd1 vccd1 vccd1 _10207_/A
+ sky130_fd_sc_hd__a211oi_2
XFILLER_121_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10091_ _10091_/A _10091_/B _10091_/C vssd1 vssd1 vccd1 vccd1 _10094_/A sky130_fd_sc_hd__nor3_1
XFILLER_126_98 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_58 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_584 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13850_ _13849_/A _13849_/B _13849_/C vssd1 vssd1 vccd1 vccd1 _13958_/A sky130_fd_sc_hd__o21a_1
XFILLER_75_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12801_ _12801_/A _12801_/B vssd1 vssd1 vccd1 vccd1 _12817_/A sky130_fd_sc_hd__xnor2_1
XFILLER_16_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10993_ _11164_/A _10992_/Y _10993_/C _10993_/D vssd1 vssd1 vccd1 vccd1 _11164_/B
+ sky130_fd_sc_hd__and4bb_1
X_13781_ _13781_/A _13781_/B vssd1 vssd1 vccd1 vccd1 _13784_/A sky130_fd_sc_hd__xor2_1
XFILLER_56_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_1012 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15520_ _15520_/A _15520_/B _15520_/C vssd1 vssd1 vccd1 vccd1 _15521_/B sky130_fd_sc_hd__or3_1
XFILLER_15_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12732_ _12566_/A _12568_/B _12566_/B vssd1 vssd1 vccd1 vccd1 _12739_/A sky130_fd_sc_hd__o21ba_1
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_879 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15451_ _15374_/B _15375_/X _15374_/A vssd1 vssd1 vccd1 vccd1 _15453_/C sky130_fd_sc_hd__o21bai_1
X_12663_ _12663_/A _12663_/B vssd1 vssd1 vccd1 vccd1 _12665_/A sky130_fd_sc_hd__nor2_1
XFILLER_31_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14402_ _14296_/X _14404_/C1 _14399_/X _14466_/B vssd1 vssd1 vccd1 vccd1 _14424_/A
+ sky130_fd_sc_hd__o211a_1
X_11614_ _11614_/A _11614_/B _11614_/C vssd1 vssd1 vccd1 vccd1 _11617_/B sky130_fd_sc_hd__and3_1
XFILLER_129_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15382_ _15381_/A _15713_/B1 _14929_/X _14803_/A vssd1 vssd1 vccd1 vccd1 _15382_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_156_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12594_ _13051_/B _13035_/C _13908_/B _13182_/A vssd1 vssd1 vccd1 vccd1 _12596_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_169_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17121_ _17121_/A _17121_/B vssd1 vssd1 vccd1 vccd1 _17124_/A sky130_fd_sc_hd__xnor2_1
XFILLER_7_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14333_ _14333_/A _14333_/B vssd1 vssd1 vccd1 vccd1 _14333_/Y sky130_fd_sc_hd__nand2_1
X_11545_ _11502_/B _11543_/A _11544_/Y _11461_/B vssd1 vssd1 vccd1 vccd1 _11705_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_156_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17052_ _17052_/A _17052_/B _17050_/X vssd1 vssd1 vccd1 vccd1 _17053_/B sky130_fd_sc_hd__or3b_1
X_11476_ _11433_/A _11433_/C _11433_/B vssd1 vssd1 vccd1 vccd1 _11477_/C sky130_fd_sc_hd__a21o_1
XFILLER_156_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14264_ _14190_/A _14190_/B _14151_/A vssd1 vssd1 vccd1 vccd1 _14266_/B sky130_fd_sc_hd__a21o_1
XFILLER_137_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16003_ _16004_/A _16004_/B vssd1 vssd1 vccd1 vccd1 _16003_/X sky130_fd_sc_hd__or2_1
X_10427_ _10427_/A _10427_/B _10427_/C vssd1 vssd1 vccd1 vccd1 _10437_/B sky130_fd_sc_hd__nand3_1
X_13215_ _13215_/A _13346_/A vssd1 vssd1 vccd1 vccd1 _13216_/C sky130_fd_sc_hd__and2_1
XFILLER_109_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14195_ _14195_/A _14195_/B vssd1 vssd1 vccd1 vccd1 _14197_/C sky130_fd_sc_hd__xor2_1
XFILLER_152_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13146_ _13625_/A _14735_/A1 _12037_/A _13145_/Y _14636_/A vssd1 vssd1 vccd1 vccd1
+ _13146_/X sky130_fd_sc_hd__a311o_1
X_10358_ _10358_/A _10358_/B vssd1 vssd1 vccd1 vccd1 _10383_/A sky130_fd_sc_hd__xnor2_1
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13077_ _13074_/X _13075_/Y _12933_/B _12935_/A vssd1 vssd1 vccd1 vccd1 _13121_/B
+ sky130_fd_sc_hd__a211oi_2
XFILLER_111_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10289_ _10289_/A _10289_/B vssd1 vssd1 vccd1 vccd1 _10305_/A sky130_fd_sc_hd__nand2_1
X_16905_ _16905_/A _16905_/B vssd1 vssd1 vccd1 vccd1 _16908_/A sky130_fd_sc_hd__xnor2_1
X_12028_ _12020_/Y _12022_/Y _12024_/Y _12026_/Y _14948_/A _15384_/S vssd1 vssd1 vccd1
+ vccd1 _12028_/X sky130_fd_sc_hd__mux4_1
XFILLER_78_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16836_ _16836_/A _16836_/B vssd1 vssd1 vccd1 vccd1 _16838_/A sky130_fd_sc_hd__nor2_1
XFILLER_66_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16767_ _16767_/A _16767_/B vssd1 vssd1 vccd1 vccd1 _16835_/B sky130_fd_sc_hd__nor2_1
XFILLER_19_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13979_ _14155_/A _14063_/C vssd1 vssd1 vccd1 vccd1 _13980_/B sky130_fd_sc_hd__nand2_1
XFILLER_65_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15718_ _16485_/A _15707_/Y _15708_/X _15717_/Y vssd1 vssd1 vccd1 vccd1 _15718_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_18_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16698_ _16698_/A _16698_/B vssd1 vssd1 vccd1 vccd1 _16699_/B sky130_fd_sc_hd__and2_1
XFILLER_80_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15649_ _16226_/B _16152_/A _15557_/A _15554_/Y vssd1 vssd1 vccd1 vccd1 _15651_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_22_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09170_ _09170_/A _09170_/B vssd1 vssd1 vccd1 vccd1 _09178_/C sky130_fd_sc_hd__xor2_1
XFILLER_159_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17319_ input38/X _17359_/B _17359_/C vssd1 vssd1 vccd1 vccd1 _17319_/X sky130_fd_sc_hd__or3_1
XFILLER_174_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08954_ _09755_/A _11930_/B _11895_/D _12275_/D vssd1 vssd1 vccd1 vccd1 _08958_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_130_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08885_ _17395_/A _11859_/D _09030_/C _17397_/A vssd1 vssd1 vccd1 vccd1 _08887_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_56_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09506_ _09499_/Y _09658_/A _09500_/X vssd1 vssd1 vccd1 vccd1 _09508_/B sky130_fd_sc_hd__a21boi_1
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09437_ _09437_/A _09437_/B _09456_/B vssd1 vssd1 vccd1 vccd1 _09437_/X sky130_fd_sc_hd__and3_1
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09368_ _09498_/A _09489_/B vssd1 vssd1 vccd1 vccd1 _09370_/C sky130_fd_sc_hd__nand2_1
XFILLER_123_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_882 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09299_ _17385_/A _09299_/B _09446_/D _11867_/D vssd1 vssd1 vccd1 vccd1 _09302_/A
+ sky130_fd_sc_hd__and4_1
XANTENNA_60 _10743_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_71 _15151_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11330_ _11331_/B _11331_/C _11331_/A vssd1 vssd1 vccd1 vccd1 _11341_/A sky130_fd_sc_hd__a21o_1
XANTENNA_82 _17496_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_93 _10743_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_31 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11261_ _11261_/A _11304_/A vssd1 vssd1 vccd1 vccd1 _11270_/A sky130_fd_sc_hd__nor2_1
XFILLER_153_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13000_ _13001_/A _13001_/B _13001_/C vssd1 vssd1 vccd1 vccd1 _13002_/A sky130_fd_sc_hd__a21oi_1
X_10212_ _10212_/A _10212_/B vssd1 vssd1 vccd1 vccd1 _10214_/B sky130_fd_sc_hd__xnor2_1
XFILLER_106_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11192_ _11067_/Y _11069_/X _11222_/B _11191_/X vssd1 vssd1 vccd1 vccd1 _11194_/A
+ sky130_fd_sc_hd__a211oi_1
XFILLER_121_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10143_ _10145_/A _15707_/A vssd1 vssd1 vccd1 vccd1 _10148_/B sky130_fd_sc_hd__nor2_1
XFILLER_122_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10074_ _10074_/A _10074_/B vssd1 vssd1 vccd1 vccd1 _10075_/B sky130_fd_sc_hd__nand2_1
X_14951_ _15180_/B _14950_/X _15103_/S vssd1 vssd1 vccd1 vccd1 _15460_/B sky130_fd_sc_hd__mux2_1
XFILLER_94_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_521 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13902_ _13902_/A _13902_/B vssd1 vssd1 vccd1 vccd1 _13904_/A sky130_fd_sc_hd__nand2_1
XFILLER_47_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14882_ _15262_/A _15262_/C _15262_/D vssd1 vssd1 vccd1 vccd1 _14882_/X sky130_fd_sc_hd__or3_1
X_16621_ _16622_/A _16622_/B _16622_/C vssd1 vssd1 vccd1 vccd1 _16699_/A sky130_fd_sc_hd__o21a_1
X_13833_ _12845_/X _12849_/B _13833_/S vssd1 vssd1 vccd1 vccd1 _13834_/A sky130_fd_sc_hd__mux2_1
XFILLER_46_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16552_ _16455_/A _16455_/B _16456_/Y vssd1 vssd1 vccd1 vccd1 _16554_/B sky130_fd_sc_hd__a21bo_1
X_13764_ _13966_/A _14213_/B _13866_/D _13764_/D vssd1 vssd1 vccd1 vccd1 _13765_/B
+ sky130_fd_sc_hd__and4_1
X_10976_ _10976_/A _10976_/B vssd1 vssd1 vccd1 vccd1 _10978_/B sky130_fd_sc_hd__xnor2_1
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15503_ _15504_/A _15504_/B vssd1 vssd1 vccd1 vccd1 _15590_/B sky130_fd_sc_hd__nand2_1
X_12715_ _12715_/A _12715_/B vssd1 vssd1 vccd1 vccd1 _12717_/A sky130_fd_sc_hd__nor2_1
X_16483_ _16390_/Y _16395_/Y _16481_/X _16482_/Y _16917_/A vssd1 vssd1 vccd1 vccd1
+ _16483_/X sky130_fd_sc_hd__o311a_1
X_13695_ _13695_/A _13695_/B _13695_/C vssd1 vssd1 vccd1 vccd1 _13697_/A sky130_fd_sc_hd__or3_1
XFILLER_148_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15434_ _15359_/A _15359_/B _15351_/X vssd1 vssd1 vccd1 vccd1 _15436_/B sky130_fd_sc_hd__o21ai_1
X_12646_ _12795_/A _14778_/B _12645_/C vssd1 vssd1 vccd1 vccd1 _12647_/B sky130_fd_sc_hd__a21o_1
XFILLER_169_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_1015 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15365_ _15366_/B _15365_/B vssd1 vssd1 vccd1 vccd1 _15365_/X sky130_fd_sc_hd__and2b_1
XFILLER_168_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12577_ _12577_/A _12577_/B vssd1 vssd1 vccd1 vccd1 _12579_/A sky130_fd_sc_hd__nor2_1
XFILLER_50_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17104_ _14597_/B _14827_/Y _14826_/X _14492_/A vssd1 vssd1 vccd1 vccd1 _17104_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_172_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14316_ _14316_/A _14316_/B vssd1 vssd1 vccd1 vccd1 _14333_/A sky130_fd_sc_hd__nand2_1
X_11528_ _11527_/A _11527_/B _11526_/Y vssd1 vssd1 vccd1 vccd1 _11530_/B sky130_fd_sc_hd__o21bai_1
XFILLER_117_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15296_ _15296_/A _15296_/B vssd1 vssd1 vccd1 vccd1 _15299_/A sky130_fd_sc_hd__xnor2_1
XFILLER_144_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17035_ _17035_/A _17035_/B _17035_/C vssd1 vssd1 vccd1 vccd1 _17035_/X sky130_fd_sc_hd__and3_1
X_14247_ _14247_/A _14330_/A vssd1 vssd1 vccd1 vccd1 _14248_/C sky130_fd_sc_hd__and2_1
XFILLER_171_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11459_ _11458_/A _11458_/B _11458_/C vssd1 vssd1 vccd1 vccd1 _11460_/C sky130_fd_sc_hd__a21oi_1
XFILLER_139_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14178_ _14090_/A _14090_/B _14088_/B vssd1 vssd1 vccd1 vccd1 _14180_/B sky130_fd_sc_hd__o21ai_1
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13129_ _12987_/X _12993_/A _13127_/X _13128_/Y vssd1 vssd1 vccd1 vccd1 _13264_/A
+ sky130_fd_sc_hd__o211a_1
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_860 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_885 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16819_ _16819_/A _16888_/B vssd1 vssd1 vccd1 vccd1 _16822_/A sky130_fd_sc_hd__nand2_1
XFILLER_26_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09222_ _09221_/A _09221_/B _09221_/C vssd1 vssd1 vccd1 vccd1 _09223_/B sky130_fd_sc_hd__o21a_1
XFILLER_22_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09153_ _09153_/A _09153_/B _09153_/C vssd1 vssd1 vccd1 vccd1 _09153_/X sky130_fd_sc_hd__or3_1
XFILLER_21_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09084_ _09084_/A _09088_/A _09084_/C vssd1 vssd1 vccd1 vccd1 _09091_/B sky130_fd_sc_hd__or3_1
XFILLER_107_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_635 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_957 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09986_ _09986_/A _09986_/B vssd1 vssd1 vccd1 vccd1 _09988_/A sky130_fd_sc_hd__nor2_1
XFILLER_130_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08937_ _08937_/A _08953_/A vssd1 vssd1 vccd1 vccd1 _08946_/A sky130_fd_sc_hd__or2_1
XFILLER_97_690 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08868_ _08869_/A _08869_/B _08869_/C vssd1 vssd1 vccd1 vccd1 _08868_/X sky130_fd_sc_hd__a21o_2
XFILLER_57_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_77 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08799_ _11911_/B _08799_/B vssd1 vssd1 vccd1 vccd1 _08801_/C sky130_fd_sc_hd__and2_1
X_10830_ _11092_/A _11092_/B vssd1 vssd1 vccd1 vccd1 _11072_/C sky130_fd_sc_hd__nand2_1
XFILLER_16_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10761_ _10761_/A vssd1 vssd1 vccd1 vccd1 _10761_/Y sky130_fd_sc_hd__inv_2
XFILLER_40_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_618 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12500_ _17405_/A _12500_/B vssd1 vssd1 vccd1 vccd1 _12501_/B sky130_fd_sc_hd__nand2_1
X_10692_ _10667_/A _10667_/C _10667_/B vssd1 vssd1 vccd1 vccd1 _10692_/X sky130_fd_sc_hd__o21a_1
XFILLER_9_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13480_ _13595_/A _13480_/B vssd1 vssd1 vccd1 vccd1 _13482_/B sky130_fd_sc_hd__and2_1
XFILLER_160_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12431_ _12432_/A _12432_/B vssd1 vssd1 vccd1 vccd1 _12607_/B sky130_fd_sc_hd__and2b_1
XFILLER_8_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15150_ _15208_/C _15208_/D _14905_/C _15149_/X _08731_/A vssd1 vssd1 vccd1 vccd1
+ _15152_/B sky130_fd_sc_hd__o32a_1
XFILLER_32_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12362_ _12526_/B _12361_/B _12361_/C vssd1 vssd1 vccd1 vccd1 _12364_/B sky130_fd_sc_hd__a21o_1
XFILLER_165_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14101_ _14188_/B _14101_/B _14102_/B vssd1 vssd1 vccd1 vccd1 _14195_/A sky130_fd_sc_hd__and3_1
X_11313_ _11313_/A _11313_/B vssd1 vssd1 vccd1 vccd1 _11331_/A sky130_fd_sc_hd__xnor2_1
X_12293_ _12143_/A _12143_/B _12146_/A vssd1 vssd1 vccd1 vccd1 _12311_/A sky130_fd_sc_hd__o21ai_1
X_15081_ _15081_/A _16315_/C vssd1 vssd1 vccd1 vccd1 _15342_/A sky130_fd_sc_hd__nor2_1
XFILLER_153_367 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11244_ _11306_/A _11244_/B vssd1 vssd1 vccd1 vccd1 _11308_/A sky130_fd_sc_hd__xnor2_1
X_14032_ _14032_/A _14032_/B vssd1 vssd1 vccd1 vccd1 _14034_/B sky130_fd_sc_hd__nor2_1
XFILLER_106_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11175_ _11176_/A _11176_/B _11176_/C vssd1 vssd1 vccd1 vccd1 _11175_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_80_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10126_ _14873_/B _10126_/B _10255_/B _10920_/B vssd1 vssd1 vccd1 vccd1 _10128_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15983_ _15983_/A _15983_/B vssd1 vssd1 vccd1 vccd1 _15984_/B sky130_fd_sc_hd__xnor2_1
XFILLER_67_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_543 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10057_ _10057_/A _10057_/B _10057_/C vssd1 vssd1 vccd1 vccd1 _10194_/A sky130_fd_sc_hd__and3_1
X_14934_ _12054_/A _15108_/A _14932_/Y _16799_/B1 _15553_/A vssd1 vssd1 vccd1 vccd1
+ _14934_/X sky130_fd_sc_hd__a2111o_1
XFILLER_169_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14865_ _16974_/A _14865_/B _16868_/A vssd1 vssd1 vccd1 vccd1 _17028_/B sky130_fd_sc_hd__and3_1
XFILLER_36_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16604_ _16745_/A _16604_/B _16758_/B _16743_/B vssd1 vssd1 vccd1 vccd1 _16604_/X
+ sky130_fd_sc_hd__and4_1
X_13816_ _13817_/A _13817_/B vssd1 vssd1 vccd1 vccd1 _13925_/B sky130_fd_sc_hd__nand2_1
X_17584_ fanout938/X _17584_/D vssd1 vssd1 vccd1 vccd1 _17584_/Q sky130_fd_sc_hd__dfxtp_1
X_14796_ _14796_/A _14796_/B _14796_/C _14796_/D vssd1 vssd1 vccd1 vccd1 _15051_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_91_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16535_ _16536_/A _16695_/B vssd1 vssd1 vccd1 vccd1 _16537_/B sky130_fd_sc_hd__nand2_1
X_13747_ _13747_/A vssd1 vssd1 vccd1 vccd1 _13748_/B sky130_fd_sc_hd__inv_2
X_10959_ _11010_/B _10961_/B vssd1 vssd1 vccd1 vccd1 _11043_/A sky130_fd_sc_hd__nor2_1
XFILLER_16_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16466_ _16466_/A _16466_/B vssd1 vssd1 vccd1 vccd1 _16469_/A sky130_fd_sc_hd__xnor2_2
XFILLER_149_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13678_ _13678_/A _13678_/B vssd1 vssd1 vccd1 vccd1 _13680_/C sky130_fd_sc_hd__xnor2_1
XFILLER_32_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15417_ _15417_/A _15417_/B vssd1 vssd1 vccd1 vccd1 _15419_/B sky130_fd_sc_hd__xor2_1
X_12629_ _12629_/A _12629_/B vssd1 vssd1 vccd1 vccd1 _12631_/C sky130_fd_sc_hd__xor2_1
X_16397_ _12235_/C _16397_/B vssd1 vssd1 vccd1 vccd1 _16398_/B sky130_fd_sc_hd__nand2b_1
XFILLER_129_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15348_ _15428_/A _15428_/B vssd1 vssd1 vccd1 vccd1 _15350_/B sky130_fd_sc_hd__xnor2_1
XFILLER_117_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15279_ _15279_/A _15279_/B vssd1 vssd1 vccd1 vccd1 _15281_/B sky130_fd_sc_hd__xor2_1
XFILLER_137_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17018_ _17018_/A vssd1 vssd1 vccd1 vccd1 _17018_/Y sky130_fd_sc_hd__inv_2
XFILLER_104_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout607 _15058_/S0 vssd1 vssd1 vccd1 vccd1 _14942_/A sky130_fd_sc_hd__clkbuf_4
X_09840_ _09841_/A _09839_/Y _10111_/C _09979_/C vssd1 vssd1 vccd1 vccd1 _09983_/A
+ sky130_fd_sc_hd__and4bb_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout618 _14450_/B vssd1 vssd1 vccd1 vccd1 _14738_/B sky130_fd_sc_hd__buf_2
XFILLER_99_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout629 _17508_/Q vssd1 vssd1 vccd1 vccd1 _14829_/B sky130_fd_sc_hd__buf_4
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09771_ _09812_/B _09812_/C vssd1 vssd1 vccd1 vccd1 _09773_/C sky130_fd_sc_hd__nor2_1
XFILLER_86_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08722_ _10993_/C vssd1 vssd1 vccd1 vccd1 _15036_/S sky130_fd_sc_hd__inv_2
XFILLER_39_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_708 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09205_ _09206_/A _09204_/Y _09639_/C _09843_/D vssd1 vssd1 vccd1 vccd1 _09375_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_136_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09136_ _17536_/Q _12127_/D _09176_/B _09135_/A vssd1 vssd1 vccd1 vccd1 _09170_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_108_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09067_ _09076_/A _09055_/Y _09062_/X _09294_/A vssd1 vssd1 vccd1 vccd1 _09069_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_135_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09969_ _09969_/A _09969_/B _09969_/C vssd1 vssd1 vccd1 vccd1 _09970_/B sky130_fd_sc_hd__nor3_1
XFILLER_89_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12980_ _12981_/A _12981_/B vssd1 vssd1 vccd1 vccd1 _12980_/X sky130_fd_sc_hd__or2_1
XTAP_3501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11931_ _11931_/A _11931_/B vssd1 vssd1 vccd1 vccd1 _11933_/A sky130_fd_sc_hd__nor2_1
XFILLER_40_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14650_ _14651_/B vssd1 vssd1 vccd1 vccd1 _14710_/B sky130_fd_sc_hd__inv_2
XTAP_3589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11862_ _11862_/A _11862_/B vssd1 vssd1 vccd1 vccd1 _11865_/A sky130_fd_sc_hd__xnor2_1
XTAP_2855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13601_ _13601_/A _13601_/B vssd1 vssd1 vccd1 vccd1 _13603_/C sky130_fd_sc_hd__or2_1
X_10813_ _10814_/B _10814_/A vssd1 vssd1 vccd1 vccd1 _11057_/A sky130_fd_sc_hd__nand2b_1
XFILLER_150_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14581_ _14583_/A _14583_/B _14583_/C vssd1 vssd1 vccd1 vccd1 _14582_/A sky130_fd_sc_hd__a21o_1
XFILLER_72_398 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11793_ _15262_/B _15472_/A vssd1 vssd1 vccd1 vccd1 _14876_/C sky130_fd_sc_hd__or2_1
XFILLER_25_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16320_ _16321_/A _16321_/B vssd1 vssd1 vccd1 vccd1 _16425_/A sky130_fd_sc_hd__and2b_1
XFILLER_41_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13532_ _13532_/A _13532_/B vssd1 vssd1 vccd1 vccd1 _13534_/A sky130_fd_sc_hd__nor2_1
XFILLER_14_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10744_ _10851_/B _10786_/B _10933_/C _11122_/A vssd1 vssd1 vccd1 vccd1 _10744_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_9_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16251_ _16251_/A _16251_/B vssd1 vssd1 vccd1 vccd1 _16252_/B sky130_fd_sc_hd__nor2_1
X_13463_ _13463_/A _13463_/B vssd1 vssd1 vccd1 vccd1 _13465_/A sky130_fd_sc_hd__nor2_1
X_10675_ _10769_/A _10675_/B vssd1 vssd1 vccd1 vccd1 _10677_/B sky130_fd_sc_hd__xor2_1
X_15202_ _14899_/X _14968_/X _15493_/A _11675_/B vssd1 vssd1 vccd1 vccd1 _15214_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_139_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12414_ _12722_/A _12722_/B _12871_/B _13450_/C vssd1 vssd1 vccd1 vccd1 _12415_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_173_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16182_ _16183_/A _16183_/B _16183_/C vssd1 vssd1 vccd1 vccd1 _16184_/A sky130_fd_sc_hd__o21a_1
XFILLER_126_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13394_ _13625_/A _14735_/A1 _12394_/A _13393_/Y _14636_/A vssd1 vssd1 vccd1 vccd1
+ _13394_/X sky130_fd_sc_hd__a311o_1
XFILLER_64_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15133_ _17063_/A _15094_/X _15114_/X _15132_/X vssd1 vssd1 vccd1 vccd1 _15133_/X
+ sky130_fd_sc_hd__o211a_1
X_12345_ _12175_/A _12177_/B _12175_/B vssd1 vssd1 vccd1 vccd1 _12346_/B sky130_fd_sc_hd__o21ba_1
XFILLER_142_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15064_ _15057_/X _15059_/Y _15061_/Y _15063_/Y _15312_/S _17369_/A vssd1 vssd1 vccd1
+ vccd1 _15064_/X sky130_fd_sc_hd__mux4_1
X_12276_ _12276_/A _12276_/B vssd1 vssd1 vccd1 vccd1 _12278_/A sky130_fd_sc_hd__nor2_1
XFILLER_141_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14015_ _14016_/A _14015_/B _14015_/C vssd1 vssd1 vccd1 vccd1 _14015_/X sky130_fd_sc_hd__or3_1
X_11227_ _11228_/A _11228_/B vssd1 vssd1 vccd1 vccd1 _11756_/A sky130_fd_sc_hd__and2_1
XFILLER_136_1042 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11158_ _11159_/A _11159_/B vssd1 vssd1 vccd1 vccd1 _11225_/A sky130_fd_sc_hd__or2_1
XFILLER_68_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10109_ _10236_/A _10109_/B _10594_/B _17479_/Q vssd1 vssd1 vccd1 vccd1 _10112_/A
+ sky130_fd_sc_hd__and4_1
X_11089_ _11084_/A _11084_/C _11084_/B vssd1 vssd1 vccd1 vccd1 _11090_/B sky130_fd_sc_hd__o21a_1
X_15966_ _15966_/A _15966_/B _15966_/C vssd1 vssd1 vccd1 vccd1 _15967_/B sky130_fd_sc_hd__and3_1
X_14917_ _10920_/B _10255_/B _10270_/B _10142_/B _14914_/S _14958_/A vssd1 vssd1 vccd1
+ vccd1 _14918_/B sky130_fd_sc_hd__mux4_1
XFILLER_63_310 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15897_ _16007_/A _15897_/B _15897_/C vssd1 vssd1 vccd1 vccd1 _15897_/X sky130_fd_sc_hd__or3_1
XFILLER_64_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14848_ _14906_/B _15175_/B _14848_/C vssd1 vssd1 vccd1 vccd1 _15314_/B sky130_fd_sc_hd__and3_1
XFILLER_51_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17567_ fanout934/X _17567_/D vssd1 vssd1 vccd1 vccd1 _17567_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14779_ _16108_/C _16114_/A vssd1 vssd1 vccd1 vccd1 _16112_/B sky130_fd_sc_hd__or2_1
XFILLER_32_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16518_ _16519_/A _16519_/B _16519_/C vssd1 vssd1 vccd1 vccd1 _16625_/A sky130_fd_sc_hd__a21oi_1
XFILLER_32_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17498_ fanout945/X _17498_/D vssd1 vssd1 vccd1 vccd1 _17498_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_20_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16449_ _16536_/A _16533_/B vssd1 vssd1 vccd1 vccd1 _16450_/B sky130_fd_sc_hd__nand2_1
XFILLER_143_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout404 _13735_/A vssd1 vssd1 vccd1 vccd1 _13632_/A sky130_fd_sc_hd__buf_2
XFILLER_113_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout415 _14775_/A vssd1 vssd1 vccd1 vccd1 _12871_/A sky130_fd_sc_hd__clkbuf_4
Xfanout426 _12068_/B vssd1 vssd1 vccd1 vccd1 _17399_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_86_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09823_ _09827_/A _09822_/B _09822_/A vssd1 vssd1 vccd1 vccd1 _09825_/B sky130_fd_sc_hd__o21ba_1
Xfanout437 _17527_/Q vssd1 vssd1 vccd1 vccd1 _10694_/A sky130_fd_sc_hd__clkbuf_4
Xfanout448 _13028_/A vssd1 vssd1 vccd1 vccd1 _13643_/A sky130_fd_sc_hd__buf_2
XFILLER_58_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout459 _17524_/Q vssd1 vssd1 vccd1 vccd1 _08791_/A sky130_fd_sc_hd__buf_2
XFILLER_59_649 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_958 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09754_ _09754_/A _09758_/A _09754_/C vssd1 vssd1 vccd1 vccd1 _09762_/B sky130_fd_sc_hd__or3_1
XFILLER_74_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09685_ _09773_/A _09773_/B vssd1 vssd1 vccd1 vccd1 _09812_/A sky130_fd_sc_hd__nor2_1
XFILLER_54_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_398 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_763 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_802 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_982 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10460_ _10459_/A _10459_/Y _10336_/Y _10353_/X vssd1 vssd1 vccd1 vccd1 _10463_/A
+ sky130_fd_sc_hd__a211oi_2
XFILLER_109_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09119_ _09119_/A _09119_/B _09119_/C _09119_/D vssd1 vssd1 vccd1 vccd1 _09119_/Y
+ sky130_fd_sc_hd__nand4_1
X_10391_ _10391_/A _10391_/B vssd1 vssd1 vccd1 vccd1 _10397_/A sky130_fd_sc_hd__xnor2_1
XFILLER_108_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12130_ _12131_/A _12131_/B vssd1 vssd1 vccd1 vccd1 _12343_/B sky130_fd_sc_hd__nor2_1
XFILLER_123_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12061_ _14912_/B _12061_/B vssd1 vssd1 vccd1 vccd1 _12061_/Y sky130_fd_sc_hd__nand2_1
XFILLER_78_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11012_ _11097_/C _10920_/B _10720_/A _10718_/Y vssd1 vssd1 vccd1 vccd1 _11013_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_150_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15820_ _15820_/A _16025_/A _16662_/C _16662_/D vssd1 vssd1 vccd1 vccd1 _15821_/D
+ sky130_fd_sc_hd__or4_1
XFILLER_77_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15751_ _15751_/A _15751_/B vssd1 vssd1 vccd1 vccd1 _15760_/A sky130_fd_sc_hd__xor2_1
X_12963_ _13227_/A _13352_/B _13434_/D _13321_/D vssd1 vssd1 vccd1 vccd1 _12964_/B
+ sky130_fd_sc_hd__and4_1
XTAP_3331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14702_ _14729_/B vssd1 vssd1 vccd1 vccd1 _14702_/Y sky130_fd_sc_hd__inv_2
XTAP_3364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11914_ _11915_/A _11915_/B _12148_/B _11913_/X vssd1 vssd1 vccd1 vccd1 _11914_/X
+ sky130_fd_sc_hd__a2bb2o_1
XTAP_2630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15682_ _15769_/B _15682_/B _15682_/C vssd1 vssd1 vccd1 vccd1 _15690_/A sky130_fd_sc_hd__nor3_1
XTAP_3375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12894_ _12895_/A _12895_/B vssd1 vssd1 vccd1 vccd1 _13057_/A sky130_fd_sc_hd__and2b_1
XFILLER_33_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17421_ _17421_/A _17421_/B vssd1 vssd1 vccd1 vccd1 _17421_/X sky130_fd_sc_hd__or2_1
XTAP_2663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14633_ _14633_/A _14633_/B vssd1 vssd1 vccd1 vccd1 _14638_/B sky130_fd_sc_hd__nand2_1
XFILLER_166_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11845_ _11822_/X _11844_/X _16012_/S vssd1 vssd1 vccd1 vccd1 _11845_/X sky130_fd_sc_hd__mux2_1
XTAP_2685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17352_ _11895_/C _17356_/A2 _17351_/X _17406_/C1 vssd1 vssd1 vccd1 vccd1 _17505_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14564_ _14565_/A _14612_/A _14564_/C vssd1 vssd1 vccd1 vccd1 _14566_/A sky130_fd_sc_hd__and3_1
XTAP_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11776_ _11775_/A _11773_/A _11773_/B _11774_/Y vssd1 vssd1 vccd1 vccd1 _17138_/B
+ sky130_fd_sc_hd__a31o_1
XTAP_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16303_ _16302_/A _16302_/B _16302_/C vssd1 vssd1 vccd1 vccd1 _16304_/C sky130_fd_sc_hd__a21oi_1
X_13515_ _16106_/A _13513_/Y _13619_/B _13391_/Y _13394_/X vssd1 vssd1 vccd1 vccd1
+ _17587_/D sky130_fd_sc_hd__a32o_1
X_10727_ _10721_/X _10725_/X _10714_/X _10715_/Y vssd1 vssd1 vccd1 vccd1 _10728_/B
+ sky130_fd_sc_hd__o211ai_2
X_17283_ _17571_/Q _17292_/B vssd1 vssd1 vccd1 vccd1 _17283_/X sky130_fd_sc_hd__and2_1
XFILLER_9_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14495_ _14495_/A _14495_/B vssd1 vssd1 vccd1 vccd1 _14497_/C sky130_fd_sc_hd__nor2_1
XFILLER_174_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16234_ _16410_/A _16662_/D _16234_/C vssd1 vssd1 vccd1 vccd1 _16339_/A sky130_fd_sc_hd__or3_1
XFILLER_146_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13446_ _13329_/A _13330_/B _13444_/A _13445_/Y vssd1 vssd1 vccd1 vccd1 _13607_/A
+ sky130_fd_sc_hd__a211oi_2
X_10658_ _15126_/A _11841_/B _14956_/A vssd1 vssd1 vccd1 vccd1 _10658_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_139_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16165_ _16165_/A _16165_/B _16454_/A vssd1 vssd1 vccd1 vccd1 _16279_/A sky130_fd_sc_hd__and3_1
X_13377_ _13246_/A _13249_/C _13500_/A _13376_/X vssd1 vssd1 vccd1 vccd1 _13500_/B
+ sky130_fd_sc_hd__a211oi_2
X_10589_ _10589_/A _10589_/B vssd1 vssd1 vccd1 vccd1 _10589_/X sky130_fd_sc_hd__and2_1
XFILLER_126_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15116_ _15116_/A _15116_/B _15450_/B vssd1 vssd1 vccd1 vccd1 _15117_/B sky130_fd_sc_hd__or3_1
X_12328_ _12795_/A _12328_/B _12328_/C vssd1 vssd1 vccd1 vccd1 _12498_/B sky130_fd_sc_hd__nand3_1
XFILLER_114_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16096_ _16096_/A _16096_/B _16096_/C vssd1 vssd1 vccd1 vccd1 _16203_/A sky130_fd_sc_hd__nor3_1
XFILLER_108_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15047_ _11595_/B _15804_/A2 _15713_/B1 _15042_/B vssd1 vssd1 vccd1 vccd1 _15047_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_130_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12259_ _12259_/A _12259_/B vssd1 vssd1 vccd1 vccd1 _12261_/B sky130_fd_sc_hd__xnor2_1
XFILLER_141_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_788 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16998_ _16880_/A _09424_/X _15724_/X _16937_/A vssd1 vssd1 vccd1 vccd1 _17000_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_77_980 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15949_ _16055_/A _16938_/B _16533_/B _16056_/A vssd1 vssd1 vccd1 vccd1 _15949_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_83_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_332 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09470_ _12471_/A _09755_/B _10180_/B _10309_/B vssd1 vssd1 vccd1 vccd1 _09602_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_110_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_560 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_788 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_646 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout201 _16735_/A vssd1 vssd1 vccd1 vccd1 _16653_/A sky130_fd_sc_hd__buf_2
XFILLER_160_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout212 _17359_/B vssd1 vssd1 vccd1 vccd1 _17355_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_99_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout223 _15454_/A vssd1 vssd1 vccd1 vccd1 _16917_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_86_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout234 _16008_/A2 vssd1 vssd1 vccd1 vccd1 _16799_/A2 sky130_fd_sc_hd__buf_2
XFILLER_101_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_690 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout245 _16731_/B1 vssd1 vssd1 vccd1 vccd1 _16579_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout256 _16106_/A vssd1 vssd1 vccd1 vccd1 _14756_/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_115_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_906 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09806_ _09806_/A _09806_/B vssd1 vssd1 vccd1 vccd1 _09808_/B sky130_fd_sc_hd__and2_1
Xfanout278 _08733_/Y vssd1 vssd1 vccd1 vccd1 _15523_/A sky130_fd_sc_hd__buf_4
XFILLER_28_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout289 _12212_/S vssd1 vssd1 vccd1 vccd1 _12383_/S sky130_fd_sc_hd__buf_2
XFILLER_46_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_89 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09737_ _09724_/X _09725_/Y _09732_/X _09868_/A vssd1 vssd1 vccd1 vccd1 _09740_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_55_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09668_ _09668_/A _09668_/B _09668_/C vssd1 vssd1 vccd1 vccd1 _09668_/Y sky130_fd_sc_hd__nand3_2
XFILLER_27_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_26 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09599_ _09480_/A _09480_/B _09480_/C vssd1 vssd1 vccd1 vccd1 _09599_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11630_ _11630_/A _15042_/B vssd1 vssd1 vccd1 vccd1 _11649_/A sky130_fd_sc_hd__nand2_1
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_571 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11561_ _11561_/A _11629_/B _11561_/C _11561_/D vssd1 vssd1 vccd1 vccd1 _11564_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_23_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13300_ _13658_/A _13414_/B _14181_/B _14094_/B vssd1 vssd1 vccd1 vccd1 _13301_/B
+ sky130_fd_sc_hd__and4_1
X_10512_ _14788_/A _10745_/D _10415_/A _10413_/Y vssd1 vssd1 vccd1 vccd1 _10513_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_7_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14280_ _14121_/X _14281_/B _14279_/Y _14204_/A vssd1 vssd1 vccd1 vccd1 _14280_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_11492_ _11492_/A _11492_/B vssd1 vssd1 vccd1 vccd1 _11493_/C sky130_fd_sc_hd__xnor2_1
XFILLER_10_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13231_ _13232_/A _13232_/B vssd1 vssd1 vccd1 vccd1 _13361_/A sky130_fd_sc_hd__and2b_1
XFILLER_109_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10443_ _10407_/Y _10442_/Y _10319_/Y _10354_/X vssd1 vssd1 vccd1 vccd1 _10459_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_137_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13162_ _13295_/B _13162_/B vssd1 vssd1 vccd1 vccd1 _13165_/C sky130_fd_sc_hd__nand2_1
XFILLER_40_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10374_ _10374_/A _10374_/B _10374_/C vssd1 vssd1 vccd1 vccd1 _10375_/B sky130_fd_sc_hd__or3_1
XFILLER_163_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12113_ _12113_/A _12113_/B vssd1 vssd1 vccd1 vccd1 _12115_/B sky130_fd_sc_hd__xnor2_1
XFILLER_3_976 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13093_ _13093_/A _13093_/B vssd1 vssd1 vccd1 vccd1 _13095_/A sky130_fd_sc_hd__nor2_1
X_12044_ _14912_/B _12044_/B vssd1 vssd1 vccd1 vccd1 _12044_/Y sky130_fd_sc_hd__nand2_1
X_16921_ _16921_/A _16921_/B vssd1 vssd1 vccd1 vccd1 _16922_/B sky130_fd_sc_hd__xnor2_1
XFILLER_111_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16852_ _16786_/A _16853_/A _16786_/B vssd1 vssd1 vccd1 vccd1 _16852_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_65_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_939 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout790 _15811_/A vssd1 vssd1 vccd1 vccd1 _11132_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_93_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15803_ _15801_/B _16008_/A2 _16008_/B1 _15811_/A _14944_/A vssd1 vssd1 vccd1 vccd1
+ _15803_/X sky130_fd_sc_hd__a221o_1
X_16783_ _16784_/A _16784_/B _16784_/C vssd1 vssd1 vccd1 vccd1 _16850_/A sky130_fd_sc_hd__a21oi_1
XFILLER_1_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13995_ _14387_/A _14301_/C vssd1 vssd1 vccd1 vccd1 _13997_/B sky130_fd_sc_hd__and2_1
XFILLER_65_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15734_ _15734_/A _15734_/B _16827_/A _16514_/A vssd1 vssd1 vccd1 vccd1 _15735_/B
+ sky130_fd_sc_hd__or4_1
XTAP_3150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12946_ _12946_/A _13085_/B vssd1 vssd1 vccd1 vccd1 _12947_/C sky130_fd_sc_hd__nor2_1
XTAP_3161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15665_ _15666_/A _15666_/B vssd1 vssd1 vccd1 vccd1 _15665_/Y sky130_fd_sc_hd__nand2_1
X_12877_ _13641_/A _13156_/B _12877_/C _13464_/B vssd1 vssd1 vccd1 vccd1 _13040_/A
+ sky130_fd_sc_hd__and4_1
XTAP_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17404_ input48/X _17422_/A2 _17403_/X _17406_/C1 vssd1 vssd1 vccd1 vccd1 _17530_/D
+ sky130_fd_sc_hd__o211a_1
X_14616_ _14658_/A _14616_/B vssd1 vssd1 vccd1 vccd1 _14618_/B sky130_fd_sc_hd__nor2_1
XTAP_2493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11828_ _12618_/D _12463_/D _12050_/S vssd1 vssd1 vccd1 vccd1 _11829_/B sky130_fd_sc_hd__mux2_1
XFILLER_33_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15596_ _16281_/A _16812_/A vssd1 vssd1 vccd1 vccd1 _15598_/B sky130_fd_sc_hd__nand2_1
XTAP_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17335_ input46/X _17353_/B _17353_/C vssd1 vssd1 vccd1 vccd1 _17335_/X sky130_fd_sc_hd__or3_1
XFILLER_53_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14547_ _14548_/A _14601_/A _14548_/C vssd1 vssd1 vccd1 vccd1 _14549_/A sky130_fd_sc_hd__o21a_1
X_11759_ _11759_/A _11762_/A vssd1 vssd1 vccd1 vccd1 _16641_/A sky130_fd_sc_hd__xor2_4
XFILLER_41_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17266_ _17456_/Q _17290_/A2 _17264_/X _17265_/X _17293_/C1 vssd1 vssd1 vccd1 vccd1
+ _17456_/D sky130_fd_sc_hd__o221a_1
XFILLER_146_226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14478_ _14479_/A _14479_/B vssd1 vssd1 vccd1 vccd1 _14478_/X sky130_fd_sc_hd__or2_1
XFILLER_140_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16217_ _14778_/B _16115_/B _16216_/Y vssd1 vssd1 vccd1 vccd1 _16221_/B sky130_fd_sc_hd__o21a_1
X_13429_ _13428_/A _13428_/B _13427_/X vssd1 vssd1 vccd1 vccd1 _13430_/B sky130_fd_sc_hd__o21bai_1
X_17197_ _17198_/C _17185_/X _17187_/Y _17575_/Q _17172_/Y vssd1 vssd1 vccd1 vccd1
+ _17197_/X sky130_fd_sc_hd__a221o_1
XFILLER_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16148_ _16032_/A _16034_/B _16032_/B vssd1 vssd1 vccd1 vccd1 _16155_/A sky130_fd_sc_hd__o21ba_1
XFILLER_143_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16079_ _16080_/A _16080_/B _16080_/C vssd1 vssd1 vccd1 vccd1 _16081_/A sky130_fd_sc_hd__o21ai_1
X_08970_ _12845_/S _11815_/B _12700_/C vssd1 vssd1 vccd1 vccd1 _08971_/C sky130_fd_sc_hd__a21oi_1
XFILLER_115_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_498 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_863 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput1 buttons vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__buf_4
XFILLER_65_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09522_ _09522_/A _09522_/B _09634_/A vssd1 vssd1 vccd1 vccd1 _09523_/B sky130_fd_sc_hd__nor3_1
XFILLER_71_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09453_ _09440_/X _09441_/Y _09448_/X _09579_/A vssd1 vssd1 vccd1 vccd1 _09455_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_51_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_677 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09384_ _09385_/B _09385_/A vssd1 vssd1 vccd1 vccd1 _09384_/X sky130_fd_sc_hd__and2b_1
XFILLER_20_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_524 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10090_ _10090_/A _10101_/A vssd1 vssd1 vccd1 vccd1 _10091_/C sky130_fd_sc_hd__nor2_1
XFILLER_86_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_75 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12800_ _17405_/A _13208_/C vssd1 vssd1 vccd1 vccd1 _12801_/B sky130_fd_sc_hd__nand2_1
XFILLER_27_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13780_ _13676_/A _13678_/B _13676_/B vssd1 vssd1 vccd1 vccd1 _13781_/B sky130_fd_sc_hd__o21ba_1
X_10992_ _10753_/A _10899_/D _10657_/C vssd1 vssd1 vccd1 vccd1 _10992_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_16_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_847 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12731_ _12577_/A _12579_/B _12577_/B vssd1 vssd1 vccd1 vccd1 _12741_/A sky130_fd_sc_hd__o21ba_1
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15450_ _15463_/A _15450_/B _15396_/A vssd1 vssd1 vccd1 vccd1 _15453_/B sky130_fd_sc_hd__or3b_1
X_12662_ _12662_/A _12662_/B _12662_/C vssd1 vssd1 vccd1 vccd1 _12663_/B sky130_fd_sc_hd__nor3_1
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14401_ _14401_/A vssd1 vssd1 vccd1 vccd1 _14466_/B sky130_fd_sc_hd__inv_2
X_11613_ _11613_/A _11646_/A vssd1 vssd1 vccd1 vccd1 _11614_/C sky130_fd_sc_hd__nand2_1
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15381_ _15381_/A _15381_/B vssd1 vssd1 vccd1 vccd1 _15381_/Y sky130_fd_sc_hd__nor2_1
X_12593_ _12593_/A _12775_/A vssd1 vssd1 vccd1 vccd1 _12605_/A sky130_fd_sc_hd__or2_1
X_17120_ _17119_/A _17081_/A _17038_/B _17038_/C _17086_/A vssd1 vssd1 vccd1 vccd1
+ _17121_/B sky130_fd_sc_hd__o41a_1
X_14332_ _14333_/A _14333_/B vssd1 vssd1 vccd1 vccd1 _14332_/X sky130_fd_sc_hd__or2_1
X_11544_ _11460_/B _11460_/C _11460_/A vssd1 vssd1 vccd1 vccd1 _11544_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_51_73 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17051_ _17052_/A _17052_/B _17050_/X vssd1 vssd1 vccd1 vccd1 _17091_/A sky130_fd_sc_hd__o21ba_1
XFILLER_7_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14263_ _14265_/A _14265_/B vssd1 vssd1 vccd1 vccd1 _14266_/A sky130_fd_sc_hd__nand2_1
XFILLER_171_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11475_ _11475_/A _11475_/B _11475_/C vssd1 vssd1 vccd1 vccd1 _11514_/A sky130_fd_sc_hd__and3_1
XFILLER_171_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16002_ _15891_/X _15892_/Y _15890_/X vssd1 vssd1 vccd1 vccd1 _16004_/B sky130_fd_sc_hd__a21boi_1
X_13214_ _13213_/A _13213_/B _13213_/C vssd1 vssd1 vccd1 vccd1 _13346_/A sky130_fd_sc_hd__o21ai_1
XFILLER_137_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10426_ _10427_/B _10427_/C _10427_/A vssd1 vssd1 vccd1 vccd1 _10437_/A sky130_fd_sc_hd__a21o_1
XFILLER_124_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14194_ _14194_/A _14195_/B _14102_/B vssd1 vssd1 vccd1 vccd1 _14270_/B sky130_fd_sc_hd__or3b_1
XFILLER_125_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13145_ _13625_/A _13145_/B vssd1 vssd1 vccd1 vccd1 _13145_/Y sky130_fd_sc_hd__nor2_1
X_10357_ _10262_/A _10262_/C _10262_/B vssd1 vssd1 vccd1 vccd1 _10357_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_151_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_796 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13076_ _12933_/B _12935_/A _13074_/X _13075_/Y vssd1 vssd1 vccd1 vccd1 _13121_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_78_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10288_ _10288_/A _10296_/A _10288_/C vssd1 vssd1 vccd1 vccd1 _10289_/B sky130_fd_sc_hd__or3_1
XFILLER_111_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16904_ _16905_/A _16905_/B vssd1 vssd1 vccd1 vccd1 _17008_/A sky130_fd_sc_hd__nand2_1
X_12027_ _12024_/Y _12026_/Y _15096_/S vssd1 vssd1 vccd1 vccd1 _12027_/X sky130_fd_sc_hd__mux2_1
XFILLER_66_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16835_ _16835_/A _16835_/B _16835_/C vssd1 vssd1 vccd1 vccd1 _16836_/B sky130_fd_sc_hd__nor3_1
XFILLER_66_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16766_ _16767_/A _16767_/B vssd1 vssd1 vccd1 vccd1 _16768_/A sky130_fd_sc_hd__and2_1
X_13978_ _13978_/A _13978_/B vssd1 vssd1 vccd1 vccd1 _13980_/A sky130_fd_sc_hd__nor2_1
XFILLER_80_216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12929_ _13117_/A _12929_/B vssd1 vssd1 vccd1 vccd1 _12931_/B sky130_fd_sc_hd__and2_1
X_15717_ _14924_/A _15457_/B _13273_/X _15716_/X vssd1 vssd1 vccd1 vccd1 _15717_/Y
+ sky130_fd_sc_hd__o31ai_1
X_16697_ _16697_/A _16697_/B _16697_/C vssd1 vssd1 vccd1 vccd1 _16698_/B sky130_fd_sc_hd__or3_1
XFILLER_80_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15648_ _15648_/A _15648_/B vssd1 vssd1 vccd1 vccd1 _15651_/A sky130_fd_sc_hd__xnor2_1
XFILLER_33_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_474 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_91 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15579_ _16056_/A _16065_/B _15578_/B vssd1 vssd1 vccd1 vccd1 _15580_/B sky130_fd_sc_hd__a21oi_1
X_17318_ _12340_/B _17322_/A2 _17317_/X _17388_/C1 vssd1 vssd1 vccd1 vccd1 _17488_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_174_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_568 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17249_ _17592_/Q _17291_/A2 _17291_/B1 vssd1 vssd1 vccd1 vccd1 _17249_/X sky130_fd_sc_hd__a21o_1
XFILLER_174_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08953_ _08953_/A _08959_/A _08953_/C vssd1 vssd1 vccd1 vccd1 _08962_/B sky130_fd_sc_hd__or3_1
XFILLER_102_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08884_ _11027_/B _10899_/D vssd1 vssd1 vccd1 vccd1 _16315_/A sky130_fd_sc_hd__nand2_8
XFILLER_97_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_622 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09505_ _09786_/A _09657_/B vssd1 vssd1 vccd1 vccd1 _09658_/A sky130_fd_sc_hd__and2_1
XFILLER_112_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09436_ _09436_/A _09577_/A vssd1 vssd1 vccd1 vccd1 _09456_/B sky130_fd_sc_hd__nand2_1
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09367_ _09370_/B _09367_/B vssd1 vssd1 vccd1 vccd1 _09489_/B sky130_fd_sc_hd__and2_1
XFILLER_8_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09298_ _09298_/A _09298_/B vssd1 vssd1 vccd1 vccd1 _09304_/A sky130_fd_sc_hd__nor2_1
XANTENNA_50 _14889_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_61 fanout795/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_72 _10479_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_83 _17452_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_94 _12340_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11260_ _11261_/A _11259_/Y _11423_/B _11563_/D vssd1 vssd1 vccd1 vccd1 _11304_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_4_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10211_ _10212_/A _10212_/B vssd1 vssd1 vccd1 vccd1 _10211_/Y sky130_fd_sc_hd__nand2_1
XFILLER_106_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11191_ _11222_/A _11190_/C _11190_/A vssd1 vssd1 vccd1 vccd1 _11191_/X sky130_fd_sc_hd__o21a_1
XFILLER_122_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10142_ _10142_/A _10142_/B vssd1 vssd1 vccd1 vccd1 _15707_/A sky130_fd_sc_hd__nand2_2
XFILLER_121_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_31 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14950_ _15096_/S _14949_/Y _14948_/Y _15097_/A vssd1 vssd1 vccd1 vccd1 _14950_/X
+ sky130_fd_sc_hd__a211o_1
X_10073_ _10073_/A _10073_/B vssd1 vssd1 vccd1 vccd1 _10208_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13901_ _13900_/B _13901_/B vssd1 vssd1 vccd1 vccd1 _13902_/B sky130_fd_sc_hd__nand2b_1
XFILLER_75_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14881_ _14876_/X _14880_/X _15147_/D vssd1 vssd1 vccd1 vccd1 _14881_/X sky130_fd_sc_hd__a21o_1
XFILLER_130_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16620_ _16620_/A _16774_/A vssd1 vssd1 vccd1 vccd1 _16622_/C sky130_fd_sc_hd__and2_1
X_13832_ _14421_/S _13832_/B vssd1 vssd1 vccd1 vccd1 _13832_/Y sky130_fd_sc_hd__nor2_1
XFILLER_75_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_780 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16551_ _16636_/A _16551_/B vssd1 vssd1 vccd1 vccd1 _16554_/A sky130_fd_sc_hd__nand2_1
X_13763_ _14213_/B _13866_/D _13764_/D _13966_/A vssd1 vssd1 vccd1 vccd1 _13765_/A
+ sky130_fd_sc_hd__a22oi_1
X_10975_ _10976_/A _10976_/B vssd1 vssd1 vccd1 vccd1 _11024_/B sky130_fd_sc_hd__and2_1
XFILLER_15_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12714_ _12714_/A _12869_/A _12871_/B _13334_/C vssd1 vssd1 vccd1 vccd1 _12715_/B
+ sky130_fd_sc_hd__and4_1
X_15502_ _15594_/A _15502_/B vssd1 vssd1 vccd1 vccd1 _15504_/B sky130_fd_sc_hd__nor2_1
X_16482_ _16390_/Y _16395_/Y _16481_/X vssd1 vssd1 vccd1 vccd1 _16482_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_15_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13694_ _13694_/A _13793_/B vssd1 vssd1 vccd1 vccd1 _13695_/C sky130_fd_sc_hd__nor2_1
XFILLER_30_102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15433_ _15433_/A _15433_/B vssd1 vssd1 vccd1 vccd1 _15436_/A sky130_fd_sc_hd__xor2_1
X_12645_ _12795_/A _14778_/B _12645_/C vssd1 vssd1 vccd1 vccd1 _12798_/B sky130_fd_sc_hd__nand3_1
XFILLER_157_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15364_ _15296_/A _15296_/B _15294_/Y vssd1 vssd1 vccd1 vccd1 _15365_/B sky130_fd_sc_hd__o21ai_1
X_12576_ _13035_/A _12734_/B _13704_/B _12877_/C vssd1 vssd1 vccd1 vccd1 _12577_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_7_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14315_ _14315_/A _14315_/B vssd1 vssd1 vccd1 vccd1 _14316_/B sky130_fd_sc_hd__nand2_1
X_17103_ _17156_/B _17103_/B _17102_/X vssd1 vssd1 vccd1 vccd1 _17103_/X sky130_fd_sc_hd__or3b_1
X_11527_ _11527_/A _11527_/B _11526_/Y vssd1 vssd1 vccd1 vccd1 _11534_/B sky130_fd_sc_hd__or3b_1
XFILLER_11_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15295_ _15295_/A _15295_/B vssd1 vssd1 vccd1 vccd1 _15296_/B sky130_fd_sc_hd__xor2_1
XFILLER_172_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17034_ _17021_/Y _17022_/X _17024_/X _16304_/A vssd1 vssd1 vccd1 vccd1 _17035_/C
+ sky130_fd_sc_hd__o22a_1
X_14246_ _14245_/A _14245_/B _14245_/C vssd1 vssd1 vccd1 vccd1 _14330_/A sky130_fd_sc_hd__o21ai_1
X_11458_ _11458_/A _11458_/B _11458_/C vssd1 vssd1 vccd1 vccd1 _11460_/B sky130_fd_sc_hd__and3_1
XFILLER_172_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10409_ _10402_/A _10402_/Y _10408_/Y _10315_/X vssd1 vssd1 vccd1 vccd1 _10453_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_171_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14177_ _14177_/A _14177_/B vssd1 vssd1 vccd1 vccd1 _14180_/A sky130_fd_sc_hd__xor2_1
X_11389_ _11561_/A _14850_/A vssd1 vssd1 vccd1 vccd1 _11389_/X sky130_fd_sc_hd__and2_1
XFILLER_125_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13128_ _13258_/A _13125_/X _12980_/X _12984_/A vssd1 vssd1 vccd1 vccd1 _13128_/Y
+ sky130_fd_sc_hd__o211ai_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13059_ _13060_/A _13060_/B vssd1 vssd1 vccd1 vccd1 _13199_/B sky130_fd_sc_hd__and2b_1
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_872 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16818_ _16818_/A _16818_/B vssd1 vssd1 vccd1 vccd1 _16888_/B sky130_fd_sc_hd__nand2_1
XFILLER_94_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16749_ _16883_/C _16749_/B vssd1 vssd1 vccd1 vccd1 _16750_/B sky130_fd_sc_hd__xnor2_1
XFILLER_35_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1000 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09221_ _09221_/A _09221_/B _09221_/C vssd1 vssd1 vccd1 vccd1 _09223_/A sky130_fd_sc_hd__nor3_1
XFILLER_107_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09152_ _09152_/A vssd1 vssd1 vccd1 vccd1 _09152_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_888 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09083_ _09084_/A _09084_/C vssd1 vssd1 vccd1 vccd1 _09088_/B sky130_fd_sc_hd__nor2_1
Xinput70 reset vssd1 vssd1 vccd1 vccd1 input70/X sky130_fd_sc_hd__clkbuf_2
XFILLER_174_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_390 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09985_ _10694_/A _10241_/B _10799_/B _09985_/D vssd1 vssd1 vccd1 vccd1 _09986_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_103_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08936_ _09327_/C _09350_/B _08936_/C _08936_/D vssd1 vssd1 vccd1 vccd1 _08953_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_130_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08867_ _08867_/A _08867_/B vssd1 vssd1 vccd1 vccd1 _08869_/C sky130_fd_sc_hd__or2_1
XFILLER_85_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08798_ _08798_/A _08821_/A _08798_/C vssd1 vssd1 vccd1 vccd1 _08799_/B sky130_fd_sc_hd__or3_1
XFILLER_123_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_942 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_750 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10760_ _10760_/A _10760_/B _10760_/C vssd1 vssd1 vccd1 vccd1 _10761_/A sky130_fd_sc_hd__and3_1
XFILLER_13_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09419_ _09434_/B _09434_/C _09434_/A vssd1 vssd1 vccd1 vccd1 _09436_/A sky130_fd_sc_hd__a21o_1
XFILLER_52_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10691_ _10678_/A _10677_/C _10677_/B vssd1 vssd1 vccd1 vccd1 _10691_/X sky130_fd_sc_hd__a21o_1
XFILLER_40_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12430_ _12607_/A _12430_/B vssd1 vssd1 vccd1 vccd1 _12432_/B sky130_fd_sc_hd__nor2_1
XFILLER_32_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12361_ _12526_/B _12361_/B _12361_/C vssd1 vssd1 vccd1 vccd1 _12364_/A sky130_fd_sc_hd__nand3_1
XFILLER_138_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_836 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14100_ _14011_/A _14115_/B _14010_/B _13990_/B _13990_/A vssd1 vssd1 vccd1 vccd1
+ _14102_/B sky130_fd_sc_hd__a32o_1
X_11312_ _11311_/A _11311_/C _11311_/B vssd1 vssd1 vccd1 vccd1 _11312_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_153_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15080_ _15278_/A _15647_/A vssd1 vssd1 vccd1 vccd1 _15157_/A sky130_fd_sc_hd__nand2_1
XFILLER_165_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12292_ _12289_/Y _12290_/X _12122_/A _12122_/Y vssd1 vssd1 vccd1 vccd1 _12312_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_154_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14031_ _14029_/Y _14031_/B vssd1 vssd1 vccd1 vccd1 _14122_/B sky130_fd_sc_hd__nand2b_1
X_11243_ _11306_/A _11244_/B vssd1 vssd1 vccd1 vccd1 _11249_/B sky130_fd_sc_hd__and2_1
XFILLER_153_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_711 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11174_ _11174_/A _11174_/B vssd1 vssd1 vccd1 vccd1 _11176_/C sky130_fd_sc_hd__xor2_1
XFILLER_122_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10125_ _10125_/A _10125_/B vssd1 vssd1 vccd1 vccd1 _10132_/A sky130_fd_sc_hd__xnor2_1
X_15982_ _16086_/A _16165_/B vssd1 vssd1 vccd1 vccd1 _15983_/B sky130_fd_sc_hd__nand2_1
XFILLER_48_511 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10056_ _10029_/A _10029_/B _10029_/C vssd1 vssd1 vccd1 vccd1 _10057_/C sky130_fd_sc_hd__o21ai_1
X_14933_ _14933_/A _14933_/B vssd1 vssd1 vccd1 vccd1 _14933_/Y sky130_fd_sc_hd__nor2_1
XFILLER_48_555 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14864_ _14864_/A _14864_/B vssd1 vssd1 vccd1 vccd1 _16868_/A sky130_fd_sc_hd__and2_1
XFILLER_91_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16603_ _16758_/B _16809_/C _16165_/B _16604_/B vssd1 vssd1 vccd1 vccd1 _16603_/X
+ sky130_fd_sc_hd__a22o_1
X_13815_ _13925_/A _13815_/B vssd1 vssd1 vccd1 vccd1 _13817_/B sky130_fd_sc_hd__and2_1
X_14795_ _14794_/A _15008_/A _15008_/B _11651_/A vssd1 vssd1 vccd1 vccd1 _14796_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_17_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17583_ fanout939/X _17583_/D vssd1 vssd1 vccd1 vccd1 _17583_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_901 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16534_ _16534_/A _16622_/A vssd1 vssd1 vccd1 vccd1 _16537_/A sky130_fd_sc_hd__nor2_1
X_13746_ _13746_/A _13858_/A vssd1 vssd1 vccd1 vccd1 _13747_/A sky130_fd_sc_hd__or2_1
X_10958_ _11005_/A _17469_/D _10955_/Y _10957_/B vssd1 vssd1 vccd1 vccd1 _10961_/B
+ sky130_fd_sc_hd__a22oi_1
XFILLER_32_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_945 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16465_ _16466_/A _16466_/B vssd1 vssd1 vccd1 vccd1 _16557_/B sky130_fd_sc_hd__nor2_1
X_13677_ _14155_/A _14141_/D vssd1 vssd1 vccd1 vccd1 _13678_/B sky130_fd_sc_hd__nand2_1
X_10889_ _11281_/A _10933_/C _11131_/B vssd1 vssd1 vccd1 vccd1 _10891_/C sky130_fd_sc_hd__and3_1
X_12628_ _12629_/B _12629_/A vssd1 vssd1 vccd1 vccd1 _12820_/B sky130_fd_sc_hd__nand2b_1
X_15416_ _15417_/A _15417_/B vssd1 vssd1 vccd1 vccd1 _15416_/Y sky130_fd_sc_hd__nor2_1
X_16396_ _16396_/A _16396_/B vssd1 vssd1 vccd1 vccd1 _16396_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_157_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15347_ _15428_/A _15428_/B vssd1 vssd1 vccd1 vccd1 _15429_/A sky130_fd_sc_hd__nand2_1
X_12559_ _12235_/C _12869_/C _12557_/X vssd1 vssd1 vccd1 vccd1 _12560_/B sky130_fd_sc_hd__a21bo_1
XFILLER_117_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15278_ _15278_/A _15397_/A vssd1 vssd1 vccd1 vccd1 _15279_/B sky130_fd_sc_hd__nand2_1
XFILLER_117_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14229_ _14229_/A _14229_/B _14229_/C vssd1 vssd1 vccd1 vccd1 _14230_/B sky130_fd_sc_hd__nor3_1
X_17017_ _14766_/A _16965_/B _17028_/A vssd1 vssd1 vccd1 vccd1 _17018_/A sky130_fd_sc_hd__a21bo_1
XFILLER_172_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout608 _15058_/S0 vssd1 vssd1 vccd1 vccd1 _09925_/A sky130_fd_sc_hd__clkbuf_4
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout619 _17153_/A vssd1 vssd1 vccd1 vccd1 _14450_/B sky130_fd_sc_hd__buf_2
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09770_ _09812_/C vssd1 vssd1 vccd1 vccd1 _09770_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08721_ _12845_/S vssd1 vssd1 vccd1 vccd1 _08721_/Y sky130_fd_sc_hd__inv_2
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09204_ _09514_/B _09937_/B _12127_/C _09942_/A vssd1 vssd1 vccd1 vccd1 _09204_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_22_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_1022 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09135_ _09135_/A _09135_/B vssd1 vssd1 vccd1 vccd1 _09176_/B sky130_fd_sc_hd__nor2_1
XFILLER_135_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09066_ _09293_/A _09293_/B vssd1 vssd1 vccd1 vccd1 _09294_/A sky130_fd_sc_hd__and2_1
XFILLER_136_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_655 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09968_ _09968_/A _09968_/B _09970_/A vssd1 vssd1 vccd1 vccd1 _11778_/A sky130_fd_sc_hd__or3_1
X_08919_ _09321_/C _11902_/B vssd1 vssd1 vccd1 vccd1 _08923_/A sky130_fd_sc_hd__nand2_1
XFILLER_76_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_1004 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09899_ _09899_/A _09899_/B _10308_/B _10657_/B vssd1 vssd1 vccd1 vccd1 _10034_/A
+ sky130_fd_sc_hd__and4_1
XTAP_3502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_20 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11930_ _17373_/A _11930_/B _12592_/D _12439_/D vssd1 vssd1 vccd1 vccd1 _11931_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_73_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_160 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11861_ _12070_/A _11861_/B vssd1 vssd1 vccd1 vccd1 _11862_/B sky130_fd_sc_hd__nand2_1
XTAP_3579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13600_ _13600_/A _13600_/B vssd1 vssd1 vccd1 vccd1 _13601_/B sky130_fd_sc_hd__and2_1
X_10812_ _10812_/A _10823_/A vssd1 vssd1 vccd1 vccd1 _10814_/B sky130_fd_sc_hd__nor2_1
XTAP_2867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14580_ _14627_/B _14580_/B vssd1 vssd1 vccd1 vccd1 _14583_/C sky130_fd_sc_hd__or2_1
XFILLER_13_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11792_ _16809_/A _16136_/A _15262_/A vssd1 vssd1 vccd1 vccd1 _14888_/C sky130_fd_sc_hd__or3_2
XTAP_2889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13531_ _13852_/A _13745_/B _13846_/B _13738_/B vssd1 vssd1 vccd1 vccd1 _13532_/B
+ sky130_fd_sc_hd__and4_1
X_10743_ _11122_/A _10851_/B _10743_/C _10743_/D vssd1 vssd1 vccd1 vccd1 _10746_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_25_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16250_ _16250_/A _16250_/B _16250_/C vssd1 vssd1 vccd1 vccd1 _16251_/B sky130_fd_sc_hd__nor3_1
X_13462_ _13462_/A _13462_/B _13462_/C vssd1 vssd1 vccd1 vccd1 _13463_/B sky130_fd_sc_hd__and3_1
XFILLER_174_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10674_ _10769_/A _10675_/B vssd1 vssd1 vccd1 vccd1 _10674_/Y sky130_fd_sc_hd__nor2_1
XFILLER_41_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15201_ _15726_/A _16536_/A vssd1 vssd1 vccd1 vccd1 _15218_/A sky130_fd_sc_hd__nand2_1
X_12413_ _12722_/B _12871_/B _13450_/C _12722_/A vssd1 vssd1 vccd1 vccd1 _12415_/A
+ sky130_fd_sc_hd__a22oi_1
X_16181_ _16181_/A _16181_/B vssd1 vssd1 vccd1 vccd1 _16183_/C sky130_fd_sc_hd__xnor2_1
XFILLER_154_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13393_ _13625_/A _13393_/B vssd1 vssd1 vccd1 vccd1 _13393_/Y sky130_fd_sc_hd__nor2_1
XFILLER_154_611 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15132_ _15119_/Y _15120_/X _15106_/Y vssd1 vssd1 vccd1 vccd1 _15132_/X sky130_fd_sc_hd__o21a_1
X_12344_ _12344_/A _12344_/B vssd1 vssd1 vccd1 vccd1 _12346_/A sky130_fd_sc_hd__nor2_1
XFILLER_153_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15063_ _15131_/A _15063_/B vssd1 vssd1 vccd1 vccd1 _15063_/Y sky130_fd_sc_hd__nand2_1
X_12275_ _12275_/A _12275_/B _12445_/D _12275_/D vssd1 vssd1 vccd1 vccd1 _12276_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_154_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14014_ _14015_/B _14015_/C vssd1 vssd1 vccd1 vccd1 _14016_/B sky130_fd_sc_hd__nor2_1
X_11226_ _11195_/A _11194_/B _11194_/A vssd1 vssd1 vccd1 vccd1 _11228_/B sky130_fd_sc_hd__o21bai_1
XFILLER_141_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11157_ _11157_/A _11157_/B vssd1 vssd1 vccd1 vccd1 _11159_/B sky130_fd_sc_hd__and2_1
XFILLER_0_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10108_ _10113_/A _10113_/B vssd1 vssd1 vccd1 vccd1 _10119_/A sky130_fd_sc_hd__nor2_1
X_15965_ _15966_/A _15966_/B _15966_/C vssd1 vssd1 vccd1 vccd1 _16084_/A sky130_fd_sc_hd__a21oi_1
X_11088_ _11088_/A _11088_/B vssd1 vssd1 vccd1 vccd1 _11232_/A sky130_fd_sc_hd__xnor2_1
XFILLER_48_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14916_ _14958_/A _14913_/Y _14915_/Y _15097_/A vssd1 vssd1 vccd1 vccd1 _14916_/X
+ sky130_fd_sc_hd__a211o_1
X_10039_ _10039_/A _10151_/A vssd1 vssd1 vccd1 vccd1 _10046_/A sky130_fd_sc_hd__nor2_1
XFILLER_63_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15896_ _16933_/A _15895_/B _15895_/C vssd1 vssd1 vccd1 vccd1 _15897_/C sky130_fd_sc_hd__a21oi_1
XFILLER_63_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14847_ _15116_/B _15110_/B vssd1 vssd1 vccd1 vccd1 _14848_/C sky130_fd_sc_hd__and2_1
XFILLER_36_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17566_ fanout952/X _17566_/D vssd1 vssd1 vccd1 vccd1 _17566_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14778_ _16209_/C _14778_/B vssd1 vssd1 vccd1 vccd1 _14778_/X sky130_fd_sc_hd__or2_1
X_16517_ _16517_/A _16517_/B vssd1 vssd1 vccd1 vccd1 _16519_/C sky130_fd_sc_hd__xnor2_1
XFILLER_149_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13729_ _13514_/A _13729_/B vssd1 vssd1 vccd1 vccd1 _13935_/A sky130_fd_sc_hd__nand2b_1
XFILLER_90_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17497_ fanout945/X _17497_/D vssd1 vssd1 vccd1 vccd1 _17497_/Q sky130_fd_sc_hd__dfxtp_4
X_16448_ _16533_/A _16165_/B _16533_/C _16447_/Y vssd1 vssd1 vccd1 vccd1 _16450_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_149_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16379_ _16285_/A _16285_/B _16287_/Y vssd1 vssd1 vccd1 vccd1 _16381_/B sky130_fd_sc_hd__a21bo_1
XFILLER_9_982 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_633 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout405 _13948_/A vssd1 vssd1 vccd1 vccd1 _13735_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_63_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout416 _17529_/Q vssd1 vssd1 vccd1 vccd1 _14775_/A sky130_fd_sc_hd__clkbuf_4
Xfanout427 _17528_/Q vssd1 vssd1 vccd1 vccd1 _12068_/B sky130_fd_sc_hd__buf_4
XFILLER_59_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09822_ _09822_/A _09822_/B vssd1 vssd1 vccd1 vccd1 _09827_/B sky130_fd_sc_hd__nor2_1
XFILLER_63_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_274 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout438 _17527_/Q vssd1 vssd1 vccd1 vccd1 _10591_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_141_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout449 _09412_/A vssd1 vssd1 vccd1 vccd1 _13028_/A sky130_fd_sc_hd__buf_4
XFILLER_150_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09753_ _09754_/A _09754_/C vssd1 vssd1 vccd1 vccd1 _09758_/B sky130_fd_sc_hd__nor2_1
XFILLER_100_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09684_ _09626_/A _09629_/B _09626_/C vssd1 vssd1 vccd1 vccd1 _09773_/B sky130_fd_sc_hd__a21oi_1
XTAP_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_994 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_77 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09118_ _09119_/A _09119_/D vssd1 vssd1 vccd1 vccd1 _09257_/B sky130_fd_sc_hd__nand2_1
XFILLER_159_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10390_ _10390_/A _10390_/B _10390_/C vssd1 vssd1 vccd1 vccd1 _10402_/B sky130_fd_sc_hd__nand3_1
XFILLER_124_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09049_ _09050_/A _09049_/B _09049_/C vssd1 vssd1 vccd1 vccd1 _09261_/A sky130_fd_sc_hd__nand3_2
XFILLER_2_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_647 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12060_ _17302_/A1 _15003_/B _14942_/A vssd1 vssd1 vccd1 vccd1 _12061_/B sky130_fd_sc_hd__mux2_1
XFILLER_104_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11011_ _11025_/B _11025_/A vssd1 vssd1 vccd1 vccd1 _11022_/A sky130_fd_sc_hd__nand2b_1
XFILLER_131_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout950 fanout957/X vssd1 vssd1 vccd1 vccd1 fanout950/X sky130_fd_sc_hd__clkbuf_2
XFILLER_131_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15750_ _15750_/A _16259_/B _15751_/A vssd1 vssd1 vccd1 vccd1 _15750_/X sky130_fd_sc_hd__and3_1
X_12962_ _13352_/B _13434_/D _13321_/D _14153_/A vssd1 vssd1 vccd1 vccd1 _12964_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_38_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_992 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11913_ _12148_/A _11911_/Y _08863_/X _08867_/A vssd1 vssd1 vccd1 vccd1 _11913_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_45_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14701_ _14701_/A _14701_/B vssd1 vssd1 vccd1 vccd1 _14729_/B sky130_fd_sc_hd__nor2_1
XTAP_3354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12893_ _13043_/B _12893_/B vssd1 vssd1 vccd1 vccd1 _12895_/B sky130_fd_sc_hd__nor2_1
XFILLER_46_878 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_804 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15681_ _15588_/A _15588_/B _15563_/Y vssd1 vssd1 vccd1 vccd1 _15682_/C sky130_fd_sc_hd__a21oi_1
XTAP_3376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17420_ input56/X _17424_/A2 _17419_/X _17420_/C1 vssd1 vssd1 vccd1 vccd1 _17538_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_33_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11844_ _11827_/X _11832_/X _11838_/X _11843_/X _17367_/A _13833_/S vssd1 vssd1 vccd1
+ vccd1 _11844_/X sky130_fd_sc_hd__mux4_1
X_14632_ _14633_/A _14633_/B vssd1 vssd1 vccd1 vccd1 _14632_/X sky130_fd_sc_hd__or2_1
XFILLER_127_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_51 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17351_ input55/X _17353_/B _17353_/C vssd1 vssd1 vccd1 vccd1 _17351_/X sky130_fd_sc_hd__or3_1
X_14563_ _14612_/A _14564_/C vssd1 vssd1 vccd1 vccd1 _14565_/B sky130_fd_sc_hd__and2_1
XTAP_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11775_ _11775_/A _11775_/B vssd1 vssd1 vccd1 vccd1 _11775_/Y sky130_fd_sc_hd__nand2_1
XFILLER_159_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16302_ _16302_/A _16302_/B _16302_/C vssd1 vssd1 vccd1 vccd1 _16304_/B sky130_fd_sc_hd__and3_1
X_10726_ _10714_/X _10715_/Y _10721_/X _10725_/X vssd1 vssd1 vccd1 vccd1 _10728_/A
+ sky130_fd_sc_hd__a211o_1
X_13514_ _13514_/A _13514_/B vssd1 vssd1 vccd1 vccd1 _13619_/B sky130_fd_sc_hd__or2_1
XFILLER_147_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17282_ _17603_/Q _17282_/A2 _17282_/B1 vssd1 vssd1 vccd1 vccd1 _17282_/X sky130_fd_sc_hd__a21o_1
X_14494_ _14554_/A _14708_/D _14493_/C vssd1 vssd1 vccd1 vccd1 _14495_/B sky130_fd_sc_hd__a21oi_1
XFILLER_158_279 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16233_ _16809_/A _16317_/B _15397_/A _16743_/C vssd1 vssd1 vccd1 vccd1 _16235_/A
+ sky130_fd_sc_hd__a22o_1
X_13445_ _13443_/A _13443_/B _13443_/C vssd1 vssd1 vccd1 vccd1 _13445_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_127_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10657_ _10753_/A _10657_/B _10657_/C vssd1 vssd1 vccd1 vccd1 _10660_/A sky130_fd_sc_hd__and3_1
XFILLER_155_931 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_110 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16164_ _16165_/A _16695_/B vssd1 vssd1 vccd1 vccd1 _16164_/Y sky130_fd_sc_hd__nand2_1
X_13376_ _13376_/A1 _13374_/X _13249_/A _13249_/Y vssd1 vssd1 vccd1 vccd1 _13376_/X
+ sky130_fd_sc_hd__o211a_1
X_10588_ _10519_/A _10519_/C _10519_/B vssd1 vssd1 vccd1 vccd1 _10588_/X sky130_fd_sc_hd__o21a_1
XFILLER_6_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_817 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12327_ _12327_/A _12498_/A vssd1 vssd1 vccd1 vccd1 _12328_/C sky130_fd_sc_hd__and2_1
XFILLER_86_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15115_ _15116_/A _15450_/B _15116_/B vssd1 vssd1 vccd1 vccd1 _15117_/A sky130_fd_sc_hd__o21ai_1
XFILLER_170_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16095_ _16095_/A _16095_/B vssd1 vssd1 vccd1 vccd1 _16096_/C sky130_fd_sc_hd__xnor2_2
XFILLER_142_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_327 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15046_ _15008_/A _15008_/B _15042_/B vssd1 vssd1 vccd1 vccd1 _15046_/Y sky130_fd_sc_hd__a21oi_1
X_12258_ _13302_/A _12258_/B vssd1 vssd1 vccd1 vccd1 _12259_/B sky130_fd_sc_hd__nand2_1
XFILLER_79_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11209_ _11168_/A _11168_/Y _11719_/A _11208_/Y vssd1 vssd1 vccd1 vccd1 _11719_/B
+ sky130_fd_sc_hd__o211ai_1
X_12189_ _12189_/A _12189_/B vssd1 vssd1 vccd1 vccd1 _12190_/B sky130_fd_sc_hd__nand2_1
XFILLER_69_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16997_ _16997_/A _17052_/A vssd1 vssd1 vccd1 vccd1 _17000_/A sky130_fd_sc_hd__nor2_1
XFILLER_23_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15948_ _16055_/A _16827_/C vssd1 vssd1 vccd1 vccd1 _16361_/A sky130_fd_sc_hd__or2_2
XFILLER_77_992 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15879_ _15773_/B _15775_/B _15773_/A vssd1 vssd1 vccd1 vccd1 _15881_/B sky130_fd_sc_hd__o21ba_1
XFILLER_63_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17549_ fanout939/X _17549_/D vssd1 vssd1 vccd1 vccd1 _17549_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout202 _11849_/Y vssd1 vssd1 vccd1 vccd1 _16735_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_99_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout213 _17362_/C vssd1 vssd1 vccd1 vccd1 _17359_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_59_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout224 _16799_/B1 vssd1 vssd1 vccd1 vccd1 _16974_/B sky130_fd_sc_hd__clkbuf_4
Xfanout235 _14928_/Y vssd1 vssd1 vccd1 vccd1 _16008_/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_87_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout246 _16731_/B1 vssd1 vssd1 vccd1 vccd1 _16015_/A sky130_fd_sc_hd__buf_2
XFILLER_59_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09805_ _09805_/A _09805_/B _09939_/A vssd1 vssd1 vccd1 vccd1 _09806_/B sky130_fd_sc_hd__or3_1
XFILLER_101_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout257 _16106_/A vssd1 vssd1 vccd1 vccd1 _16922_/A sky130_fd_sc_hd__buf_4
XFILLER_115_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout268 _17153_/B vssd1 vssd1 vccd1 vccd1 _16571_/B sky130_fd_sc_hd__buf_2
Xfanout279 _16911_/A vssd1 vssd1 vccd1 vccd1 _17131_/A sky130_fd_sc_hd__buf_4
XFILLER_75_918 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_823 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09736_ _09867_/A _09867_/B vssd1 vssd1 vccd1 vccd1 _09868_/A sky130_fd_sc_hd__and2_1
XFILLER_83_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09667_ _09628_/A _09628_/B _09628_/C vssd1 vssd1 vccd1 vccd1 _09668_/C sky130_fd_sc_hd__o21ai_1
XFILLER_131_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_78 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09598_ _09624_/B _09624_/C _09624_/A vssd1 vssd1 vccd1 vccd1 _09627_/A sky130_fd_sc_hd__o21a_1
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_336 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11560_ _11565_/A _11565_/B vssd1 vssd1 vccd1 vccd1 _11566_/A sky130_fd_sc_hd__nor2_1
XFILLER_24_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10511_ _10511_/A _10511_/B vssd1 vssd1 vccd1 vccd1 _10613_/A sky130_fd_sc_hd__xnor2_1
XFILLER_128_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11491_ _11444_/Y _11466_/X _11487_/A _11527_/A vssd1 vssd1 vccd1 vccd1 _11493_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_149_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13230_ _13230_/A _13230_/B vssd1 vssd1 vccd1 vccd1 _13232_/B sky130_fd_sc_hd__xnor2_1
XFILLER_137_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10442_ _10473_/A _10473_/B vssd1 vssd1 vccd1 vccd1 _10442_/Y sky130_fd_sc_hd__nor2_1
XFILLER_164_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13161_ _13161_/A _13161_/B vssd1 vssd1 vccd1 vccd1 _13162_/B sky130_fd_sc_hd__or2_1
XFILLER_156_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10373_ _10374_/A _10374_/B _10374_/C vssd1 vssd1 vccd1 vccd1 _10390_/A sky130_fd_sc_hd__o21ai_1
XFILLER_136_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12112_ _12113_/B _12113_/A vssd1 vssd1 vccd1 vccd1 _12112_/X sky130_fd_sc_hd__and2b_1
XFILLER_2_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13092_ _13092_/A _13092_/B _13092_/C vssd1 vssd1 vccd1 vccd1 _13093_/B sky130_fd_sc_hd__and3_1
XFILLER_97_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_988 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12043_ _12770_/D _12618_/D _14942_/A vssd1 vssd1 vccd1 vccd1 _12044_/B sky130_fd_sc_hd__mux2_1
X_16920_ _10784_/A _10784_/B _11766_/X vssd1 vssd1 vccd1 vccd1 _16921_/B sky130_fd_sc_hd__o21ai_1
XFILLER_133_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16851_ _16851_/A _16851_/B vssd1 vssd1 vccd1 vccd1 _16931_/A sky130_fd_sc_hd__nand2_1
XFILLER_131_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_907 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout780 _10786_/B vssd1 vssd1 vccd1 vccd1 _10932_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_92_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout791 fanout795/X vssd1 vssd1 vccd1 vccd1 _15811_/A sky130_fd_sc_hd__clkbuf_4
X_15802_ _15802_/A _15802_/B vssd1 vssd1 vccd1 vccd1 _15802_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_65_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16782_ _16846_/B _16782_/B vssd1 vssd1 vccd1 vccd1 _16784_/C sky130_fd_sc_hd__or2_1
XFILLER_18_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13994_ _16864_/A _16918_/A _13991_/X vssd1 vssd1 vccd1 vccd1 _13997_/A sky130_fd_sc_hd__o21a_1
XFILLER_1_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15733_ _15647_/A _16604_/B _16758_/B _16129_/A vssd1 vssd1 vccd1 vccd1 _15735_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_74_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12945_ _12945_/A _13085_/A _12945_/C vssd1 vssd1 vccd1 vccd1 _13085_/B sky130_fd_sc_hd__nor3_1
XTAP_3162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15664_ _16410_/A _16446_/A vssd1 vssd1 vccd1 vccd1 _15666_/B sky130_fd_sc_hd__nor2_1
XFILLER_73_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12876_ _13156_/B _12877_/C _13464_/B _13641_/A vssd1 vssd1 vccd1 vccd1 _12878_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_73_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17403_ _17403_/A _17421_/B vssd1 vssd1 vccd1 vccd1 _17403_/X sky130_fd_sc_hd__or2_1
X_14615_ _14614_/B _14615_/B vssd1 vssd1 vccd1 vccd1 _14616_/B sky130_fd_sc_hd__and2b_1
XTAP_2483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11827_ _11824_/Y _11826_/Y _17365_/A vssd1 vssd1 vccd1 vccd1 _11827_/X sky130_fd_sc_hd__mux2_1
XTAP_2494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15595_ _15595_/A _15595_/B vssd1 vssd1 vccd1 vccd1 _15598_/A sky130_fd_sc_hd__nand2_1
XTAP_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17334_ _09446_/D _17356_/A2 _17333_/X _17422_/C1 vssd1 vssd1 vccd1 vccd1 _17496_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_42_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11758_ _11758_/A _11758_/B vssd1 vssd1 vccd1 vccd1 _11762_/A sky130_fd_sc_hd__nor2_2
X_14546_ _14676_/A _14641_/D vssd1 vssd1 vccd1 vccd1 _14548_/C sky130_fd_sc_hd__nand2_1
XFILLER_159_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10709_ _10709_/A _10709_/B vssd1 vssd1 vccd1 vccd1 _11180_/B sky130_fd_sc_hd__xor2_2
X_17265_ _17565_/Q _17289_/B vssd1 vssd1 vccd1 vccd1 _17265_/X sky130_fd_sc_hd__and2_1
X_11689_ _15302_/A _15302_/B vssd1 vssd1 vccd1 vccd1 _15303_/A sky130_fd_sc_hd__nand2_1
X_14477_ _14533_/A _14419_/B _14414_/A vssd1 vssd1 vccd1 vccd1 _14479_/B sky130_fd_sc_hd__a21oi_1
XFILLER_146_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16216_ _14859_/B _16115_/B _16579_/A vssd1 vssd1 vccd1 vccd1 _16216_/Y sky130_fd_sc_hd__a21oi_1
X_13428_ _13428_/A _13428_/B _13427_/X vssd1 vssd1 vccd1 vccd1 _13430_/A sky130_fd_sc_hd__or3b_1
X_17196_ input29/X _17196_/B _17196_/C vssd1 vssd1 vccd1 vccd1 _17196_/X sky130_fd_sc_hd__or3_1
XFILLER_115_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16147_ _16040_/A _16040_/B _16043_/A vssd1 vssd1 vccd1 vccd1 _16157_/A sky130_fd_sc_hd__a21bo_1
X_13359_ _13360_/B _13360_/A vssd1 vssd1 vccd1 vccd1 _13477_/B sky130_fd_sc_hd__and2b_1
XFILLER_142_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16078_ _16183_/B _16078_/B vssd1 vssd1 vccd1 vccd1 _16080_/C sky130_fd_sc_hd__nor2_1
XFILLER_142_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15029_ _15820_/A _15687_/A _15028_/A vssd1 vssd1 vccd1 vccd1 _15030_/D sky130_fd_sc_hd__o21ai_1
XFILLER_123_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput2 clk vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__clkbuf_1
XFILLER_84_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09521_ _09522_/B _09634_/A _09522_/A vssd1 vssd1 vccd1 vccd1 _09523_/A sky130_fd_sc_hd__o21a_1
XFILLER_36_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09452_ _09578_/A _09578_/B vssd1 vssd1 vccd1 vccd1 _09579_/A sky130_fd_sc_hd__and2_1
XFILLER_80_932 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09383_ _09383_/A _09511_/A vssd1 vssd1 vccd1 vccd1 _09385_/B sky130_fd_sc_hd__nor2_1
XFILLER_51_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_199 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_536 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_975 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_912 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_200 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09719_ _09720_/A _09719_/B _09719_/C vssd1 vssd1 vccd1 vccd1 _09866_/A sky130_fd_sc_hd__nand3_1
X_10991_ _10991_/A _11841_/B _10991_/C vssd1 vssd1 vccd1 vccd1 _11164_/A sky130_fd_sc_hd__and3_1
XFILLER_56_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12730_ _12730_/A _12730_/B _12730_/C vssd1 vssd1 vccd1 vccd1 _12743_/B sky130_fd_sc_hd__nand3_1
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12661_ _12662_/A _12662_/B _12662_/C vssd1 vssd1 vccd1 vccd1 _12663_/A sky130_fd_sc_hd__o21a_1
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_818 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11612_ _11613_/A _11612_/B _11612_/C vssd1 vssd1 vccd1 vccd1 _11646_/A sky130_fd_sc_hd__nand3_1
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14400_ _14400_/A _14466_/A _14400_/C vssd1 vssd1 vccd1 vccd1 _14401_/A sky130_fd_sc_hd__and3_1
XFILLER_169_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12592_ _12592_/A _12592_/B _12592_/C _12592_/D vssd1 vssd1 vccd1 vccd1 _12775_/A
+ sky130_fd_sc_hd__and4_1
X_15380_ _15102_/Y _15123_/Y _15125_/Y _15131_/Y _15312_/S _15116_/A vssd1 vssd1 vccd1
+ vccd1 _15380_/X sky130_fd_sc_hd__mux4_1
XFILLER_23_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_531 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11543_ _11543_/A _11543_/B _11542_/X vssd1 vssd1 vccd1 vccd1 _11586_/A sky130_fd_sc_hd__or3b_1
XFILLER_156_514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14331_ _14409_/A _14331_/B vssd1 vssd1 vccd1 vccd1 _14333_/B sky130_fd_sc_hd__or2_1
XFILLER_7_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17050_ _17088_/B _17050_/B vssd1 vssd1 vccd1 vccd1 _17050_/X sky130_fd_sc_hd__or2_1
XFILLER_51_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14262_ _14262_/A _14340_/A _14262_/C vssd1 vssd1 vccd1 vccd1 _14265_/B sky130_fd_sc_hd__or3_1
X_11474_ _11430_/A _11430_/C _11430_/B vssd1 vssd1 vccd1 vccd1 _11475_/C sky130_fd_sc_hd__o21ai_1
XFILLER_109_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_761 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13213_ _13213_/A _13213_/B _13213_/C vssd1 vssd1 vccd1 vccd1 _13215_/A sky130_fd_sc_hd__or3_1
XFILLER_100_1012 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16001_ _16001_/A _16001_/B vssd1 vssd1 vccd1 vccd1 _16004_/A sky130_fd_sc_hd__nand2_1
XFILLER_171_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10425_ _10427_/B _10427_/C _10427_/A vssd1 vssd1 vccd1 vccd1 _10425_/Y sky130_fd_sc_hd__a21oi_1
X_14193_ _14270_/A _14193_/B vssd1 vssd1 vccd1 vccd1 _14195_/B sky130_fd_sc_hd__nand2_1
XFILLER_136_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13144_ _12028_/X _12056_/X _13516_/S vssd1 vssd1 vccd1 vccd1 _13145_/B sky130_fd_sc_hd__mux2_1
X_10356_ _10283_/X _10356_/B vssd1 vssd1 vccd1 vccd1 _10441_/A sky130_fd_sc_hd__nand2b_1
XFILLER_152_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13075_ _13075_/A _13075_/B _13075_/C vssd1 vssd1 vccd1 vccd1 _13075_/Y sky130_fd_sc_hd__nand3_2
XFILLER_3_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10287_ _10187_/X _10285_/Y _10283_/C _10266_/X vssd1 vssd1 vccd1 vccd1 _10287_/Y
+ sky130_fd_sc_hd__o211ai_2
X_16903_ _16838_/A _16838_/B _16836_/A vssd1 vssd1 vccd1 vccd1 _16905_/B sky130_fd_sc_hd__a21o_1
XFILLER_2_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12026_ _14949_/A _14948_/C _14911_/B vssd1 vssd1 vccd1 vccd1 _12026_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_78_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16834_ _16835_/A _16835_/B _16835_/C vssd1 vssd1 vccd1 vccd1 _16836_/A sky130_fd_sc_hd__o21a_1
XFILLER_65_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16765_ _16765_/A _16765_/B vssd1 vssd1 vccd1 vccd1 _16767_/B sky130_fd_sc_hd__or2_1
XFILLER_20_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13977_ _13977_/A _13977_/B _14213_/C _14213_/D vssd1 vssd1 vccd1 vccd1 _13978_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_46_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15716_ _14963_/X _15715_/X _15714_/Y _15712_/X _15710_/X vssd1 vssd1 vccd1 vccd1
+ _15716_/X sky130_fd_sc_hd__o2111a_1
X_12928_ _12928_/A _12928_/B _12928_/C vssd1 vssd1 vccd1 vccd1 _12929_/B sky130_fd_sc_hd__or3_1
XFILLER_80_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16696_ _16697_/A _16697_/B _16697_/C vssd1 vssd1 vccd1 vccd1 _16698_/A sky130_fd_sc_hd__o21ai_1
XFILLER_33_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15647_ _15647_/A _16152_/A vssd1 vssd1 vccd1 vccd1 _15648_/B sky130_fd_sc_hd__nand2_1
XFILLER_33_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12859_ _17164_/A _12857_/X _12858_/Y _13837_/C vssd1 vssd1 vccd1 vccd1 _15457_/C
+ sky130_fd_sc_hd__o22a_1
XTAP_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15578_ _16056_/A _15578_/B _16065_/B vssd1 vssd1 vccd1 vccd1 _15580_/A sky130_fd_sc_hd__and3_1
X_17317_ input37/X _17321_/B _17321_/C vssd1 vssd1 vccd1 vccd1 _17317_/X sky130_fd_sc_hd__or3_1
XFILLER_30_851 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14529_ _14583_/B _14529_/B vssd1 vssd1 vccd1 vccd1 _14531_/C sky130_fd_sc_hd__and2_1
XFILLER_147_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17248_ _17450_/Q _17293_/A2 _17246_/X _17247_/X _17284_/C1 vssd1 vssd1 vccd1 vccd1
+ _17450_/D sky130_fd_sc_hd__o221a_1
X_17179_ input10/X input13/X input12/X input16/X vssd1 vssd1 vccd1 vccd1 _17180_/D
+ sky130_fd_sc_hd__or4_1
XFILLER_103_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_274 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08952_ _08953_/A _08953_/C vssd1 vssd1 vccd1 vccd1 _08959_/B sky130_fd_sc_hd__nor2_1
XFILLER_130_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08883_ _08883_/A _08883_/B _08889_/B vssd1 vssd1 vccd1 vccd1 _08904_/B sky130_fd_sc_hd__or3_1
XFILLER_96_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09504_ _09504_/A _09504_/B vssd1 vssd1 vccd1 vccd1 _09657_/B sky130_fd_sc_hd__nor2_1
XFILLER_72_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09435_ _09436_/A _09435_/B _09435_/C vssd1 vssd1 vccd1 vccd1 _09577_/A sky130_fd_sc_hd__nand3_1
XFILLER_169_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09366_ _09366_/A _09366_/B _09366_/C vssd1 vssd1 vccd1 vccd1 _09367_/B sky130_fd_sc_hd__nand3_1
XFILLER_21_851 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09297_ _17381_/A _09319_/D _09061_/A _09059_/Y vssd1 vssd1 vccd1 vccd1 _09298_/B
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA_40 fanout380/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_51 _17153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_62 _10525_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_73 _09981_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_84 _17464_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_95 _09979_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10210_ _10210_/A _10210_/B vssd1 vssd1 vccd1 vccd1 _10212_/B sky130_fd_sc_hd__xnor2_1
XFILLER_97_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11190_ _11190_/A _11222_/A _11190_/C vssd1 vssd1 vccd1 vccd1 _11222_/B sky130_fd_sc_hd__nor3_1
XFILLER_106_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10141_ _10142_/A _10142_/B vssd1 vssd1 vccd1 vccd1 _10145_/B sky130_fd_sc_hd__and2_2
XFILLER_106_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10072_ _10560_/B _10072_/B _10073_/A vssd1 vssd1 vccd1 vccd1 _10072_/Y sky130_fd_sc_hd__nand3_1
XFILLER_94_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_726 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13900_ _13901_/B _13900_/B vssd1 vssd1 vccd1 vccd1 _13902_/A sky130_fd_sc_hd__nand2b_1
XFILLER_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14880_ _15147_/C _15262_/D _14877_/Y vssd1 vssd1 vccd1 vccd1 _14880_/X sky130_fd_sc_hd__a21o_1
XFILLER_47_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13831_ _12844_/X _12852_/B _13831_/S vssd1 vssd1 vccd1 vccd1 _13832_/B sky130_fd_sc_hd__mux2_1
XFILLER_75_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16550_ _16550_/A _16550_/B _16550_/C vssd1 vssd1 vccd1 vccd1 _16551_/B sky130_fd_sc_hd__nand3_1
XFILLER_15_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10974_ _10974_/A _10974_/B vssd1 vssd1 vccd1 vccd1 _10976_/B sky130_fd_sc_hd__xnor2_1
X_13762_ _13762_/A _13762_/B vssd1 vssd1 vccd1 vccd1 _13768_/A sky130_fd_sc_hd__nor2_1
XFILLER_44_943 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15501_ _15501_/A _15501_/B _15501_/C vssd1 vssd1 vccd1 vccd1 _15502_/B sky130_fd_sc_hd__nor3_1
X_12713_ _12869_/A _12871_/B _13334_/C _12714_/A vssd1 vssd1 vccd1 vccd1 _12715_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_31_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16481_ _16481_/A _16481_/B vssd1 vssd1 vccd1 vccd1 _16481_/X sky130_fd_sc_hd__and2_1
X_13693_ _16796_/A _13693_/B _13793_/A vssd1 vssd1 vccd1 vccd1 _13793_/B sky130_fd_sc_hd__nor3_1
XFILLER_15_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_114 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15432_ _15433_/A _15433_/B vssd1 vssd1 vccd1 vccd1 _15514_/B sky130_fd_sc_hd__nand2_1
X_12644_ _12644_/A _12798_/A vssd1 vssd1 vccd1 vccd1 _12645_/C sky130_fd_sc_hd__and2_1
XFILLER_62_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12575_ _12734_/B _13704_/B _12877_/C _17524_/Q vssd1 vssd1 vccd1 vccd1 _12577_/A
+ sky130_fd_sc_hd__a22oi_1
X_15363_ _15363_/A _15363_/B vssd1 vssd1 vccd1 vccd1 _15366_/B sky130_fd_sc_hd__xnor2_1
XFILLER_11_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17102_ _17064_/X _17067_/Y _17099_/A _17100_/X vssd1 vssd1 vccd1 vccd1 _17102_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_129_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14314_ _14315_/A _14315_/B vssd1 vssd1 vccd1 vccd1 _14316_/A sky130_fd_sc_hd__or2_1
X_11526_ _11526_/A _11526_/B vssd1 vssd1 vccd1 vccd1 _11526_/Y sky130_fd_sc_hd__nand2_1
XFILLER_117_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15294_ _15295_/A _15295_/B vssd1 vssd1 vccd1 vccd1 _15294_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17033_ _17033_/A _17033_/B _17033_/C _17033_/D vssd1 vssd1 vccd1 vccd1 _17035_/B
+ sky130_fd_sc_hd__and4_1
X_11457_ _11456_/B _11456_/C _11456_/A vssd1 vssd1 vccd1 vccd1 _11458_/C sky130_fd_sc_hd__o21bai_1
XFILLER_156_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14245_ _14245_/A _14245_/B _14245_/C vssd1 vssd1 vccd1 vccd1 _14247_/A sky130_fd_sc_hd__or3_1
XFILLER_109_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10408_ _10315_/A _10315_/B _10315_/C vssd1 vssd1 vccd1 vccd1 _10408_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_171_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14176_ _14176_/A _14385_/B _14177_/A vssd1 vssd1 vccd1 vccd1 _14252_/B sky130_fd_sc_hd__nand3_1
X_11388_ _11520_/C _14895_/B vssd1 vssd1 vccd1 vccd1 _11436_/A sky130_fd_sc_hd__nand2_1
XFILLER_140_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_571 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13127_ _12980_/X _12984_/A _13258_/A _13125_/X vssd1 vssd1 vccd1 vccd1 _13127_/X
+ sky130_fd_sc_hd__a211o_1
X_10339_ _10215_/B _10228_/Y _10336_/A _10336_/Y vssd1 vssd1 vccd1 vccd1 _10340_/B
+ sky130_fd_sc_hd__a211o_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13058_ _13199_/A _13058_/B vssd1 vssd1 vccd1 vccd1 _13060_/B sky130_fd_sc_hd__nor2_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12009_ _12009_/A vssd1 vssd1 vccd1 vccd1 _12010_/B sky130_fd_sc_hd__inv_2
XFILLER_39_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_854 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16817_ _16818_/A _16818_/B vssd1 vssd1 vccd1 vccd1 _16819_/A sky130_fd_sc_hd__or2_1
XFILLER_54_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16748_ _16814_/A _16938_/D _16748_/C vssd1 vssd1 vccd1 vccd1 _16749_/B sky130_fd_sc_hd__or3_1
XFILLER_19_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1012 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16679_ _16807_/A _16760_/B _16603_/X _16604_/X vssd1 vssd1 vccd1 vccd1 _16688_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_34_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09220_ _09220_/A _11958_/B vssd1 vssd1 vccd1 vccd1 _09221_/C sky130_fd_sc_hd__nor2_1
XFILLER_107_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09151_ _09153_/A _09153_/B _09153_/C vssd1 vssd1 vccd1 vccd1 _09152_/A sky130_fd_sc_hd__o21ai_1
XFILLER_21_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09082_ _11932_/A _11895_/C _08957_/C _08957_/D vssd1 vssd1 vccd1 vccd1 _09084_/C
+ sky130_fd_sc_hd__a22oi_1
XFILLER_174_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput60 i_wb_data[31] vssd1 vssd1 vccd1 vccd1 input60/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09984_ _10241_/B _10799_/B _14788_/B _10694_/A vssd1 vssd1 vccd1 vccd1 _09986_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_88_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_767 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08935_ _09325_/B _11895_/C _12445_/D _09755_/A vssd1 vssd1 vccd1 vccd1 _08936_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_76_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08866_ _08866_/A _08866_/B vssd1 vssd1 vccd1 vccd1 _08867_/B sky130_fd_sc_hd__nor2_1
XFILLER_85_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08797_ _08798_/A _08821_/A _08798_/C vssd1 vssd1 vccd1 vccd1 _11911_/B sky130_fd_sc_hd__o21ai_1
XFILLER_45_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_902 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09418_ _09546_/A _09546_/B vssd1 vssd1 vccd1 vccd1 _09434_/C sky130_fd_sc_hd__nand2_1
XFILLER_12_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10690_ _10690_/A _10690_/B vssd1 vssd1 vccd1 vccd1 _10779_/A sky130_fd_sc_hd__xor2_1
XFILLER_12_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09349_ _11839_/S _12025_/B vssd1 vssd1 vccd1 vccd1 _14982_/B sky130_fd_sc_hd__and2_1
XFILLER_8_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12360_ _12360_/A _12360_/B vssd1 vssd1 vccd1 vccd1 _12361_/C sky130_fd_sc_hd__nand2_1
XFILLER_120_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11311_ _11311_/A _11311_/B _11311_/C vssd1 vssd1 vccd1 vccd1 _11343_/A sky130_fd_sc_hd__or3_1
XFILLER_154_848 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12291_ _12122_/A _12122_/Y _12289_/Y _12290_/X vssd1 vssd1 vccd1 vccd1 _12312_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_10_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14030_ _14030_/A _14030_/B _14030_/C vssd1 vssd1 vccd1 vccd1 _14031_/B sky130_fd_sc_hd__nand3_1
X_11242_ _11242_/A _11242_/B vssd1 vssd1 vccd1 vccd1 _11244_/B sky130_fd_sc_hd__nor2_1
XFILLER_106_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_723 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_200 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11173_ _11202_/A _11171_/Y _10988_/Y _10999_/X vssd1 vssd1 vccd1 vccd1 _11186_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_164_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10124_ _10125_/A _10125_/B vssd1 vssd1 vccd1 vccd1 _10138_/A sky130_fd_sc_hd__nand2b_1
XFILLER_79_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15981_ _15981_/A _15981_/B vssd1 vssd1 vccd1 vccd1 _15983_/A sky130_fd_sc_hd__nor2_1
XFILLER_79_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10055_ _10055_/A _10055_/B vssd1 vssd1 vccd1 vccd1 _10057_/B sky130_fd_sc_hd__xnor2_1
X_14932_ _17070_/B _14931_/X _12054_/A vssd1 vssd1 vccd1 vccd1 _14932_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14863_ _14863_/A _14863_/B _16652_/B vssd1 vssd1 vccd1 vccd1 _14864_/B sky130_fd_sc_hd__and3_1
XFILLER_48_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16602_ _16517_/A _16517_/B _16515_/B vssd1 vssd1 vccd1 vccd1 _16611_/B sky130_fd_sc_hd__o21ai_1
X_13814_ _13814_/A wire118/X _13814_/C vssd1 vssd1 vccd1 vccd1 _13815_/B sky130_fd_sc_hd__or3_1
XFILLER_35_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17582_ fanout937/X _17582_/D vssd1 vssd1 vccd1 vccd1 _17582_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_857 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14794_ _14794_/A _15008_/A vssd1 vssd1 vccd1 vccd1 _14796_/C sky130_fd_sc_hd__or2_1
XFILLER_113_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16533_ _16533_/A _16533_/B _16533_/C vssd1 vssd1 vccd1 vccd1 _16622_/A sky130_fd_sc_hd__and3_1
XFILLER_17_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13745_ _13852_/A _13745_/B _13852_/B _13844_/C vssd1 vssd1 vccd1 vccd1 _13858_/A
+ sky130_fd_sc_hd__and4_1
X_10957_ _11010_/A _10957_/B _11005_/A _17469_/D vssd1 vssd1 vccd1 vccd1 _11010_/B
+ sky130_fd_sc_hd__and4b_1
XFILLER_43_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_83 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16464_ _16362_/A _16362_/B _16365_/A vssd1 vssd1 vccd1 vccd1 _16466_/B sky130_fd_sc_hd__a21oi_2
X_13676_ _13676_/A _13676_/B vssd1 vssd1 vccd1 vccd1 _13678_/A sky130_fd_sc_hd__nor2_1
X_10888_ _10891_/B _10888_/B vssd1 vssd1 vccd1 vccd1 _11131_/B sky130_fd_sc_hd__nor2_1
X_15415_ _15415_/A _15755_/B vssd1 vssd1 vccd1 vccd1 _15417_/B sky130_fd_sc_hd__or2_1
X_12627_ _12820_/A _12627_/B vssd1 vssd1 vccd1 vccd1 _12629_/B sky130_fd_sc_hd__nand2_1
X_16395_ _16394_/A _16394_/B _16396_/A vssd1 vssd1 vccd1 vccd1 _16395_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_169_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15346_ _15346_/A _15346_/B vssd1 vssd1 vccd1 vccd1 _15428_/B sky130_fd_sc_hd__xnor2_1
XFILLER_156_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12558_ _12714_/A _13450_/C vssd1 vssd1 vccd1 vccd1 _12869_/C sky130_fd_sc_hd__and2_4
XFILLER_157_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11509_ _11506_/X _11509_/B _11553_/B _15042_/B vssd1 vssd1 vccd1 vccd1 _11555_/A
+ sky130_fd_sc_hd__and4b_1
XFILLER_129_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15277_ _15277_/A _15277_/B vssd1 vssd1 vccd1 vccd1 _15279_/A sky130_fd_sc_hd__xor2_1
XFILLER_172_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12489_ _12490_/A _12642_/A _12490_/C vssd1 vssd1 vccd1 vccd1 _12491_/A sky130_fd_sc_hd__o21a_1
X_17016_ _17063_/A _17016_/B _17016_/C vssd1 vssd1 vccd1 vccd1 _17035_/A sky130_fd_sc_hd__or3_2
XFILLER_172_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14228_ _14229_/A _14229_/B _14229_/C vssd1 vssd1 vccd1 vccd1 _14230_/A sky130_fd_sc_hd__o21a_1
XFILLER_99_913 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14159_ _14159_/A _14159_/B vssd1 vssd1 vccd1 vccd1 _14161_/A sky130_fd_sc_hd__nor2_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout609 _15058_/S0 vssd1 vssd1 vccd1 vccd1 _14914_/S sky130_fd_sc_hd__buf_2
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08720_ _11470_/A vssd1 vssd1 vccd1 vccd1 _08720_/Y sky130_fd_sc_hd__inv_2
XFILLER_79_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_386 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09203_ _09942_/A _09514_/B _09937_/B _12127_/C vssd1 vssd1 vccd1 vccd1 _09206_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_33_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_787 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09134_ _09172_/A _11920_/D _09362_/D _09360_/A vssd1 vssd1 vccd1 vccd1 _09135_/B
+ sky130_fd_sc_hd__a22oi_1
XFILLER_136_826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09065_ _09065_/A _09065_/B vssd1 vssd1 vccd1 vccd1 _09293_/B sky130_fd_sc_hd__nor2_1
XFILLER_120_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_255 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09967_ _09969_/A _09969_/B _09969_/C vssd1 vssd1 vccd1 vccd1 _09970_/A sky130_fd_sc_hd__o21a_1
X_08918_ _08918_/A _08918_/B vssd1 vssd1 vccd1 vccd1 _09052_/A sky130_fd_sc_hd__xnor2_1
XFILLER_69_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1016 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09898_ _09898_/A _09902_/A _09898_/C vssd1 vssd1 vccd1 vccd1 _09906_/B sky130_fd_sc_hd__or3_1
XTAP_3503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08849_ _09321_/C _11895_/D _08846_/Y _08996_/A vssd1 vssd1 vccd1 vccd1 _08850_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_85_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_32 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11860_ _11860_/A _11860_/B vssd1 vssd1 vccd1 vccd1 _11862_/A sky130_fd_sc_hd__nor2_1
XTAP_2835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10811_ _10812_/A _10810_/Y _11097_/C _11115_/C vssd1 vssd1 vccd1 vccd1 _10823_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_14_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_773 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11791_ _16021_/A _16317_/A _16809_/A _16136_/A vssd1 vssd1 vccd1 vccd1 _15262_/D
+ sky130_fd_sc_hd__or4_1
XTAP_2879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13530_ _13745_/B _13846_/B _13738_/B _13852_/A vssd1 vssd1 vccd1 vccd1 _13532_/A
+ sky130_fd_sc_hd__a22oi_1
X_10742_ _10742_/A _10747_/A _10742_/C vssd1 vssd1 vccd1 vccd1 _10750_/B sky130_fd_sc_hd__or3_1
XFILLER_13_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_20 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10673_ _10673_/A _10673_/B vssd1 vssd1 vccd1 vccd1 _10675_/B sky130_fd_sc_hd__xnor2_1
XFILLER_43_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13461_ _13462_/A _13462_/B _13462_/C vssd1 vssd1 vccd1 vccd1 _13463_/A sky130_fd_sc_hd__a21oi_1
XFILLER_9_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15200_ _14887_/B _15198_/X _14924_/A vssd1 vssd1 vccd1 vccd1 _16262_/A sky130_fd_sc_hd__a21bo_2
XFILLER_40_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12412_ _12412_/A _12412_/B vssd1 vssd1 vccd1 vccd1 _12419_/A sky130_fd_sc_hd__xor2_1
X_16180_ _16279_/C _16180_/B vssd1 vssd1 vccd1 vccd1 _16181_/B sky130_fd_sc_hd__nor2_1
XFILLER_138_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13392_ _12387_/X _12391_/X _13840_/S vssd1 vssd1 vccd1 vccd1 _13393_/B sky130_fd_sc_hd__mux2_1
XFILLER_154_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15131_ _15131_/A _15131_/B vssd1 vssd1 vccd1 vccd1 _15131_/Y sky130_fd_sc_hd__nand2_1
X_12343_ _12343_/A _12343_/B _12343_/C vssd1 vssd1 vccd1 vccd1 _12344_/B sky130_fd_sc_hd__nor3_1
XFILLER_154_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12274_ _12275_/B _12445_/D _12275_/D _12275_/A vssd1 vssd1 vccd1 vccd1 _12276_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_4_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15062_ _17302_/A1 _15116_/B _15175_/B _14906_/B _14942_/A _15095_/B vssd1 vssd1
+ vccd1 vccd1 _15063_/B sky130_fd_sc_hd__mux4_1
XFILLER_153_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_188 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11225_ _11225_/A _11225_/B vssd1 vssd1 vccd1 vccd1 _11228_/A sky130_fd_sc_hd__xnor2_1
X_14013_ _14013_/A _14013_/B _14013_/C vssd1 vssd1 vccd1 vccd1 _14015_/C sky130_fd_sc_hd__and3_1
XFILLER_136_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11156_ _11155_/A _11234_/A _11232_/A vssd1 vssd1 vccd1 vccd1 _11201_/A sky130_fd_sc_hd__o21ai_1
X_10107_ _10111_/C _09981_/D _09982_/A _09980_/Y vssd1 vssd1 vccd1 vccd1 _10113_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_1_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15964_ _15964_/A _15964_/B vssd1 vssd1 vccd1 vccd1 _15966_/C sky130_fd_sc_hd__xnor2_1
X_11087_ _11087_/A _11087_/B vssd1 vssd1 vccd1 vccd1 _11088_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14915_ _14958_/A _14915_/B vssd1 vssd1 vccd1 vccd1 _14915_/Y sky130_fd_sc_hd__nor2_1
X_10038_ _10039_/A _10037_/Y _10970_/A _11841_/B vssd1 vssd1 vccd1 vccd1 _10151_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_64_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15895_ _16933_/A _15895_/B _15895_/C vssd1 vssd1 vccd1 vccd1 _15897_/B sky130_fd_sc_hd__and3_1
XFILLER_91_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14846_ _15274_/A _14846_/B vssd1 vssd1 vccd1 vccd1 _15110_/B sky130_fd_sc_hd__nor2_1
XFILLER_63_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17565_ fanout953/X _17565_/D vssd1 vssd1 vccd1 vccd1 _17565_/Q sky130_fd_sc_hd__dfxtp_1
X_14777_ _14777_/A _16298_/A vssd1 vssd1 vccd1 vccd1 _16302_/B sky130_fd_sc_hd__or2_1
XFILLER_32_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11989_ _11990_/A _11990_/B _11990_/C vssd1 vssd1 vccd1 vccd1 _12155_/A sky130_fd_sc_hd__a21oi_1
XFILLER_16_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_721 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16516_ _16745_/A _16760_/B vssd1 vssd1 vccd1 vccd1 _16517_/B sky130_fd_sc_hd__nand2_1
XFILLER_90_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13728_ _13619_/A _13616_/Y _13617_/X vssd1 vssd1 vccd1 vccd1 _13728_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_56_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17496_ fanout945/X _17496_/D vssd1 vssd1 vccd1 vccd1 _17496_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_149_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16447_ _16533_/A _16355_/B _16352_/C vssd1 vssd1 vccd1 vccd1 _16447_/Y sky130_fd_sc_hd__a21oi_1
X_13659_ _13659_/A _13659_/B vssd1 vssd1 vccd1 vccd1 _13662_/C sky130_fd_sc_hd__xnor2_1
XFILLER_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16378_ _16378_/A _16378_/B vssd1 vssd1 vccd1 vccd1 _16381_/A sky130_fd_sc_hd__xnor2_2
XFILLER_157_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_994 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15329_ _15553_/A _15553_/B _16619_/A vssd1 vssd1 vccd1 vccd1 _15331_/B sky130_fd_sc_hd__or3_1
XFILLER_129_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout406 _12714_/A vssd1 vssd1 vccd1 vccd1 _13948_/A sky130_fd_sc_hd__buf_2
Xfanout417 _12070_/A vssd1 vssd1 vccd1 vccd1 _17401_/A sky130_fd_sc_hd__clkbuf_4
X_09821_ _09819_/A _09819_/B _09819_/C vssd1 vssd1 vccd1 vccd1 _09822_/B sky130_fd_sc_hd__o21a_1
XFILLER_87_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout428 _17528_/Q vssd1 vssd1 vccd1 vccd1 _10236_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_141_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout439 _12722_/B vssd1 vssd1 vccd1 vccd1 _13745_/B sky130_fd_sc_hd__buf_2
XFILLER_140_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09752_ _15538_/A _10180_/B _09746_/A _09612_/Y vssd1 vssd1 vccd1 vccd1 _09754_/C
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_100_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09683_ _09668_/A _09668_/C _09668_/B vssd1 vssd1 vccd1 vccd1 _09683_/X sky130_fd_sc_hd__a21o_1
XFILLER_67_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_838 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_89 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09117_ _08930_/X _09018_/Y _09071_/A _09259_/A vssd1 vssd1 vccd1 vccd1 _09119_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_108_325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09048_ _09048_/A _09048_/B _09048_/C vssd1 vssd1 vccd1 vccd1 _09049_/C sky130_fd_sc_hd__nand3_1
XFILLER_163_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11010_ _11010_/A _11010_/B vssd1 vssd1 vccd1 vccd1 _11025_/B sky130_fd_sc_hd__nor2_1
XFILLER_145_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout940 fanout941/X vssd1 vssd1 vccd1 vccd1 fanout940/X sky130_fd_sc_hd__buf_2
XFILLER_104_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_139 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout951 fanout952/X vssd1 vssd1 vccd1 vccd1 fanout951/X sky130_fd_sc_hd__clkbuf_2
XFILLER_92_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12961_ _12771_/A _12773_/B _12771_/B vssd1 vssd1 vccd1 vccd1 _12968_/A sky130_fd_sc_hd__o21ba_1
XFILLER_46_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14700_ _14701_/A _14701_/B vssd1 vssd1 vccd1 vccd1 _14700_/Y sky130_fd_sc_hd__nand2_1
XTAP_3344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11912_ _08863_/X _08867_/A _12148_/A _11911_/Y vssd1 vssd1 vccd1 vccd1 _12148_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_46_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15680_ _15772_/B _15679_/C _15679_/A vssd1 vssd1 vccd1 vccd1 _15682_/B sky130_fd_sc_hd__a21oi_1
XTAP_2621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12892_ _13302_/A _13035_/C _12889_/Y _13043_/A vssd1 vssd1 vccd1 vccd1 _12893_/B
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_3366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_816 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14631_ _14631_/A _14631_/B vssd1 vssd1 vccd1 vccd1 _14633_/B sky130_fd_sc_hd__or2_1
XTAP_3399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11843_ _11840_/Y _11842_/Y _17365_/A vssd1 vssd1 vccd1 vccd1 _11843_/X sky130_fd_sc_hd__mux2_1
XTAP_2665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17350_ _11895_/D _17356_/A2 _17349_/X _17406_/C1 vssd1 vssd1 vccd1 vccd1 _17504_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_72_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14562_ _14562_/A _14562_/B _14562_/C vssd1 vssd1 vccd1 vccd1 _14564_/C sky130_fd_sc_hd__nand3_1
XTAP_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11774_ _10347_/X _11775_/B _11775_/A vssd1 vssd1 vccd1 vccd1 _11774_/Y sky130_fd_sc_hd__a21boi_1
XTAP_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16301_ _16301_/A _16301_/B vssd1 vssd1 vccd1 vccd1 _16301_/Y sky130_fd_sc_hd__xnor2_1
X_13513_ _13514_/A _13514_/B vssd1 vssd1 vccd1 vccd1 _13513_/Y sky130_fd_sc_hd__nand2_1
XFILLER_158_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10725_ _11174_/A _11174_/B vssd1 vssd1 vccd1 vccd1 _10725_/X sky130_fd_sc_hd__and2_1
XFILLER_14_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17281_ _17461_/Q _17293_/A2 _17279_/X _17280_/X _17284_/C1 vssd1 vssd1 vccd1 vccd1
+ _17461_/D sky130_fd_sc_hd__o221a_1
XTAP_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14493_ _14554_/A _14708_/D _14493_/C vssd1 vssd1 vccd1 vccd1 _14495_/A sky130_fd_sc_hd__and3_1
XFILLER_174_707 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16232_ _16232_/A _16232_/B vssd1 vssd1 vccd1 vccd1 _16239_/A sky130_fd_sc_hd__xor2_1
X_13444_ _13444_/A vssd1 vssd1 vccd1 vccd1 _13444_/Y sky130_fd_sc_hd__inv_2
XFILLER_174_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10656_ _11651_/A _11841_/B vssd1 vssd1 vccd1 vccd1 _10657_/C sky130_fd_sc_hd__and2_2
XFILLER_127_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16163_ _16044_/A _16044_/B _16045_/X vssd1 vssd1 vccd1 vccd1 _16177_/A sky130_fd_sc_hd__a21oi_1
XFILLER_70_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10587_ _10555_/A _10555_/C _10555_/B vssd1 vssd1 vccd1 vccd1 _10587_/Y sky130_fd_sc_hd__o21ai_1
X_13375_ _13249_/A _13249_/Y _13376_/A1 _13374_/X vssd1 vssd1 vccd1 vccd1 _13500_/A
+ sky130_fd_sc_hd__a211oi_2
XFILLER_155_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15114_ _15628_/A _16219_/A1 _12230_/B _15113_/X vssd1 vssd1 vccd1 vccd1 _15114_/X
+ sky130_fd_sc_hd__o31a_1
X_12326_ _12325_/A _12325_/B _12325_/C vssd1 vssd1 vccd1 vccd1 _12498_/A sky130_fd_sc_hd__o21ai_1
X_16094_ _16095_/B _16095_/A vssd1 vssd1 vccd1 vccd1 _16200_/B sky130_fd_sc_hd__nand2b_1
XFILLER_115_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15045_ _15041_/X _15042_/X _15043_/X _14938_/X vssd1 vssd1 vccd1 vccd1 _15045_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_114_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12257_ _12257_/A _12257_/B vssd1 vssd1 vccd1 vccd1 _12259_/A sky130_fd_sc_hd__nor2_1
XFILLER_170_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11208_ _10761_/A _11206_/Y _11178_/Y _11175_/Y vssd1 vssd1 vccd1 vccd1 _11208_/Y
+ sky130_fd_sc_hd__o211ai_1
X_12188_ _12188_/A _12188_/B vssd1 vssd1 vccd1 vccd1 _12189_/B sky130_fd_sc_hd__or2_1
XFILLER_123_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11139_ _11139_/A _11139_/B _11139_/C vssd1 vssd1 vccd1 vccd1 _11255_/A sky130_fd_sc_hd__and3_1
XFILLER_68_448 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16996_ _16995_/B _16996_/B vssd1 vssd1 vccd1 vccd1 _17052_/A sky130_fd_sc_hd__and2b_1
XFILLER_96_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15947_ _16880_/A _16021_/B vssd1 vssd1 vccd1 vccd1 _16827_/C sky130_fd_sc_hd__nand2_1
XFILLER_49_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15878_ _15992_/A _15878_/B vssd1 vssd1 vccd1 vccd1 _15881_/A sky130_fd_sc_hd__nand2b_1
XFILLER_24_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14829_ _17134_/A _14829_/B vssd1 vssd1 vccd1 vccd1 _14829_/X sky130_fd_sc_hd__or2_1
XFILLER_36_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17548_ fanout937/X _17548_/D vssd1 vssd1 vccd1 vccd1 _17548_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17479_ fanout949/X _17479_/D vssd1 vssd1 vccd1 vccd1 _17479_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_32_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_751 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout203 _16219_/A1 vssd1 vssd1 vccd1 vccd1 _17143_/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_8_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout214 _17196_/X vssd1 vssd1 vccd1 vccd1 _17362_/C sky130_fd_sc_hd__buf_4
XFILLER_141_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout225 _16799_/B1 vssd1 vssd1 vccd1 vccd1 _16580_/B1 sky130_fd_sc_hd__clkbuf_2
Xfanout236 _14962_/B vssd1 vssd1 vccd1 vccd1 _15808_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_113_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09804_ _09805_/B _09939_/A _09805_/A vssd1 vssd1 vccd1 vccd1 _09806_/A sky130_fd_sc_hd__o21ai_1
Xfanout247 _14844_/X vssd1 vssd1 vccd1 vccd1 _16731_/B1 sky130_fd_sc_hd__clkbuf_2
Xfanout258 _16106_/A vssd1 vssd1 vccd1 vccd1 _16389_/A sky130_fd_sc_hd__clkbuf_2
Xfanout269 _17153_/B vssd1 vssd1 vccd1 vccd1 _15450_/B sky130_fd_sc_hd__buf_2
XFILLER_86_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09735_ _09735_/A _09735_/B vssd1 vssd1 vccd1 vccd1 _09867_/B sky130_fd_sc_hd__nor2_1
XFILLER_74_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09666_ _09666_/A _09666_/B vssd1 vssd1 vccd1 vccd1 _09668_/B sky130_fd_sc_hd__and2_1
XFILLER_27_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_985 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09597_ _09597_/A _09597_/B _09686_/B vssd1 vssd1 vccd1 vccd1 _09624_/C sky130_fd_sc_hd__and3_1
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10510_ _10511_/B _10511_/A vssd1 vssd1 vccd1 vccd1 _10510_/X sky130_fd_sc_hd__and2b_1
X_11490_ _11456_/A _11456_/C _11456_/B vssd1 vssd1 vccd1 vccd1 _11490_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_168_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_910 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10441_ _10441_/A _10441_/B vssd1 vssd1 vccd1 vccd1 _10473_/B sky130_fd_sc_hd__xnor2_1
XFILLER_148_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13160_ _13161_/A _13161_/B vssd1 vssd1 vccd1 vccd1 _13295_/B sky130_fd_sc_hd__nand2_1
X_10372_ _10372_/A _10372_/B vssd1 vssd1 vccd1 vccd1 _10374_/C sky130_fd_sc_hd__xnor2_1
XFILLER_108_166 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12111_ _11901_/A _11903_/B _11901_/B vssd1 vssd1 vccd1 vccd1 _12113_/B sky130_fd_sc_hd__o21ba_1
XFILLER_123_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13091_ _13092_/A _13092_/B _13092_/C vssd1 vssd1 vccd1 vccd1 _13093_/A sky130_fd_sc_hd__a21oi_1
XFILLER_151_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_1011 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12042_ _14912_/B _12042_/B vssd1 vssd1 vccd1 vccd1 _12042_/Y sky130_fd_sc_hd__nand2_1
XFILLER_123_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16850_ _16850_/A _16850_/B vssd1 vssd1 vccd1 vccd1 _16851_/B sky130_fd_sc_hd__or2_1
XFILLER_78_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_854 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15801_ _15801_/A _15801_/B vssd1 vssd1 vccd1 vccd1 _15802_/B sky130_fd_sc_hd__and2_1
Xfanout770 _10532_/D vssd1 vssd1 vccd1 vccd1 _10897_/B sky130_fd_sc_hd__buf_4
Xfanout781 _10146_/B vssd1 vssd1 vccd1 vccd1 _10786_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_172_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16781_ _16781_/A _16781_/B vssd1 vssd1 vccd1 vccd1 _16782_/B sky130_fd_sc_hd__and2_1
Xfanout792 fanout795/X vssd1 vssd1 vccd1 vccd1 _10933_/C sky130_fd_sc_hd__buf_4
XFILLER_19_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13993_ _14167_/A _13993_/B vssd1 vssd1 vccd1 vccd1 _16918_/A sky130_fd_sc_hd__nand2_2
XTAP_3130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15732_ _15732_/A _15732_/B vssd1 vssd1 vccd1 vccd1 _15741_/A sky130_fd_sc_hd__xnor2_2
XFILLER_46_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12944_ _12945_/A _13085_/A _12945_/C vssd1 vssd1 vccd1 vccd1 _12946_/A sky130_fd_sc_hd__o21a_1
XTAP_3141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15663_ _15663_/A _15663_/B vssd1 vssd1 vccd1 vccd1 _15673_/A sky130_fd_sc_hd__xnor2_1
XTAP_3185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12875_ _12875_/A _12875_/B vssd1 vssd1 vccd1 vccd1 _12884_/A sky130_fd_sc_hd__xor2_1
XFILLER_61_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17402_ input46/X _17422_/A2 _17401_/X _17422_/C1 vssd1 vssd1 vccd1 vccd1 _17529_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_33_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14614_ _14615_/B _14614_/B vssd1 vssd1 vccd1 vccd1 _14658_/A sky130_fd_sc_hd__and2b_1
XTAP_2473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11826_ _12046_/A _11826_/B vssd1 vssd1 vccd1 vccd1 _11826_/Y sky130_fd_sc_hd__nand2_1
XTAP_2484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15594_ _15594_/A _15594_/B vssd1 vssd1 vccd1 vccd1 _15595_/B sky130_fd_sc_hd__or2_1
XTAP_2495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17333_ input45/X _17355_/B _17355_/C vssd1 vssd1 vccd1 vccd1 _17333_/X sky130_fd_sc_hd__or3_1
XFILLER_60_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14545_ _14641_/A _14641_/B _14593_/D _14545_/D vssd1 vssd1 vccd1 vccd1 _14601_/A
+ sky130_fd_sc_hd__and4_1
X_11757_ _11732_/Y _11733_/X _11737_/Y _11753_/A vssd1 vssd1 vccd1 vccd1 _11758_/B
+ sky130_fd_sc_hd__o211a_1
XTAP_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10708_ _10708_/A _10708_/B vssd1 vssd1 vccd1 vccd1 _11180_/A sky130_fd_sc_hd__xnor2_2
X_17264_ _17597_/Q _17282_/A2 _17282_/B1 vssd1 vssd1 vccd1 vccd1 _17264_/X sky130_fd_sc_hd__a21o_1
XFILLER_147_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14476_ _14533_/B _14533_/C vssd1 vssd1 vccd1 vccd1 _14479_/A sky130_fd_sc_hd__nand2_1
X_11688_ _11688_/A _11688_/B vssd1 vssd1 vccd1 vccd1 _15302_/B sky130_fd_sc_hd__xor2_1
X_16215_ _08760_/Y _14778_/X _14813_/X _15456_/B _16214_/Y vssd1 vssd1 vccd1 vccd1
+ _16215_/X sky130_fd_sc_hd__a311o_1
X_13427_ _13304_/A _13304_/B _13305_/Y vssd1 vssd1 vccd1 vccd1 _13427_/X sky130_fd_sc_hd__a21bo_1
X_10639_ _10638_/B _10933_/D _10970_/B _10638_/A vssd1 vssd1 vccd1 vccd1 _10639_/Y
+ sky130_fd_sc_hd__a22oi_1
X_17195_ _17195_/A _17195_/B _17195_/C vssd1 vssd1 vccd1 vccd1 _17196_/C sky130_fd_sc_hd__or3_1
XFILLER_10_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16146_ _16146_/A _16146_/B vssd1 vssd1 vccd1 vccd1 _16158_/A sky130_fd_sc_hd__xnor2_1
X_13358_ _13228_/A _13230_/B _13228_/B vssd1 vssd1 vccd1 vccd1 _13360_/B sky130_fd_sc_hd__o21ba_1
XFILLER_170_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12309_ _12309_/A _12309_/B _12309_/C vssd1 vssd1 vccd1 vccd1 _12310_/B sky130_fd_sc_hd__and3_1
XFILLER_5_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16077_ _16077_/A _16077_/B vssd1 vssd1 vccd1 vccd1 _16078_/B sky130_fd_sc_hd__nor2_1
XFILLER_114_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13289_ _13643_/A _13738_/B _13286_/Y _13417_/A vssd1 vssd1 vccd1 vccd1 _13290_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15028_ _15028_/A _15687_/A vssd1 vssd1 vccd1 vccd1 _15093_/A sky130_fd_sc_hd__or2_1
XFILLER_130_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_908 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput3 i_wb_addr[0] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__clkbuf_1
X_16979_ _16304_/A _16971_/Y _16972_/Y _17070_/B _16978_/X vssd1 vssd1 vccd1 vccd1
+ _16979_/X sky130_fd_sc_hd__o221a_1
XFILLER_49_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09520_ _10560_/A _09843_/D _09520_/C vssd1 vssd1 vccd1 vccd1 _09634_/A sky130_fd_sc_hd__and3_1
XFILLER_83_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_900 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09451_ _09451_/A _09451_/B vssd1 vssd1 vccd1 vccd1 _09578_/B sky130_fd_sc_hd__nor2_1
XFILLER_64_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_944 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09382_ _10560_/A _09843_/C _09382_/C vssd1 vssd1 vccd1 vccd1 _09511_/A sky130_fd_sc_hd__and3_1
XFILLER_33_860 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_910 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_621 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09718_ _09718_/A _09718_/B _09718_/C vssd1 vssd1 vccd1 vccd1 _09719_/C sky130_fd_sc_hd__nand3_1
X_10990_ _10990_/A _10990_/B _10990_/C vssd1 vssd1 vccd1 vccd1 _10999_/B sky130_fd_sc_hd__nand3_1
XFILLER_90_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09649_ _09969_/B _09649_/B vssd1 vssd1 vccd1 vccd1 _09774_/A sky130_fd_sc_hd__nor2_1
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12660_ _12660_/A _12660_/B vssd1 vssd1 vccd1 vccd1 _12662_/C sky130_fd_sc_hd__xnor2_1
XFILLER_150_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11611_ _11617_/A _11611_/B vssd1 vssd1 vccd1 vccd1 _11612_/C sky130_fd_sc_hd__and2_1
XFILLER_30_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12591_ _12592_/A _12592_/C vssd1 vssd1 vccd1 vccd1 _12759_/A sky130_fd_sc_hd__nand2_1
XFILLER_169_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14330_ _14330_/A _14330_/B _14330_/C vssd1 vssd1 vccd1 vccd1 _14331_/B sky130_fd_sc_hd__and3_1
X_11542_ _11542_/A _11584_/A vssd1 vssd1 vccd1 vccd1 _11542_/X sky130_fd_sc_hd__or2_1
XFILLER_129_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_543 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14261_ _14340_/A _14262_/C _14262_/A vssd1 vssd1 vccd1 vccd1 _14265_/A sky130_fd_sc_hd__o21ai_1
X_11473_ _11469_/X _11471_/X _11472_/A vssd1 vssd1 vccd1 vccd1 _11475_/B sky130_fd_sc_hd__a21o_1
XFILLER_51_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16000_ _16014_/A _16571_/B _16317_/A vssd1 vssd1 vccd1 vccd1 _16001_/B sky130_fd_sc_hd__or3b_1
X_13212_ _13212_/A _13339_/B vssd1 vssd1 vccd1 vccd1 _13213_/C sky130_fd_sc_hd__nor2_1
XFILLER_137_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10424_ _10524_/A _10524_/B vssd1 vssd1 vccd1 vccd1 _10427_/C sky130_fd_sc_hd__nand2_1
X_14192_ _14192_/A _14192_/B _14192_/C vssd1 vssd1 vccd1 vccd1 _14193_/B sky130_fd_sc_hd__nand3_1
XFILLER_100_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13143_ _12710_/A _13142_/X _16653_/A vssd1 vssd1 vccd1 vccd1 _13143_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_124_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10355_ _10283_/B _10283_/C _10283_/D _10283_/A vssd1 vssd1 vccd1 vccd1 _10356_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_124_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13074_ _13075_/A _13075_/B _13075_/C vssd1 vssd1 vccd1 vccd1 _13074_/X sky130_fd_sc_hd__a21o_1
X_10286_ _10266_/X _10283_/C _10285_/Y _10187_/X vssd1 vssd1 vccd1 vccd1 _10330_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_32_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16902_ _16902_/A _16902_/B vssd1 vssd1 vccd1 vccd1 _16905_/A sky130_fd_sc_hd__nor2_1
X_12025_ _12025_/A _12025_/B vssd1 vssd1 vccd1 vccd1 _14948_/C sky130_fd_sc_hd__and2_1
XFILLER_76_50 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16833_ _16833_/A _16897_/B vssd1 vssd1 vccd1 vccd1 _16835_/C sky130_fd_sc_hd__nor2_1
XFILLER_120_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_524 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16764_ _16763_/B _16764_/B vssd1 vssd1 vccd1 vccd1 _16765_/B sky130_fd_sc_hd__and2b_1
XFILLER_18_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13976_ _13977_/B _14213_/C _14213_/D _13977_/A vssd1 vssd1 vccd1 vccd1 _13978_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_18_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15715_ _15715_/A _15715_/B vssd1 vssd1 vccd1 vccd1 _15715_/X sky130_fd_sc_hd__or2_2
X_12927_ _12928_/A _12928_/B _12928_/C vssd1 vssd1 vccd1 vccd1 _13117_/A sky130_fd_sc_hd__o21ai_1
XFILLER_47_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16695_ _16695_/A _16695_/B _16695_/C vssd1 vssd1 vccd1 vccd1 _16697_/C sky130_fd_sc_hd__and3_1
XFILLER_62_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15646_ _15734_/A _15645_/B _16514_/A _15644_/X vssd1 vssd1 vccd1 vccd1 _15648_/A
+ sky130_fd_sc_hd__o31a_1
XFILLER_34_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12858_ _13516_/S _17367_/A vssd1 vssd1 vccd1 vccd1 _12858_/Y sky130_fd_sc_hd__nand2_4
XTAP_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_819 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11809_ _09652_/C _14982_/C _14911_/B vssd1 vssd1 vccd1 vccd1 _11809_/Y sky130_fd_sc_hd__o21ai_1
X_15577_ _15846_/A _16065_/B vssd1 vssd1 vccd1 vccd1 _15577_/Y sky130_fd_sc_hd__nand2_1
XFILLER_61_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12789_ _12790_/A _12947_/A _12790_/C vssd1 vssd1 vccd1 vccd1 _12791_/A sky130_fd_sc_hd__o21a_1
XTAP_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17316_ _12338_/C _17322_/A2 _17315_/X _17388_/C1 vssd1 vssd1 vccd1 vccd1 _17487_/D
+ sky130_fd_sc_hd__o211a_1
X_14528_ _14528_/A _14528_/B vssd1 vssd1 vccd1 vccd1 _14529_/B sky130_fd_sc_hd__nand2_1
XFILLER_30_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17247_ _17559_/Q _17289_/B vssd1 vssd1 vccd1 vccd1 _17247_/X sky130_fd_sc_hd__and2_1
X_14459_ _14518_/A _14459_/B _14459_/C vssd1 vssd1 vccd1 vccd1 _14518_/B sky130_fd_sc_hd__nand3_1
XFILLER_162_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17178_ input6/X input9/X input8/X input11/X vssd1 vssd1 vccd1 vccd1 _17180_/C sky130_fd_sc_hd__or4_1
X_16129_ _16129_/A _16129_/B vssd1 vssd1 vccd1 vccd1 _16130_/B sky130_fd_sc_hd__nand2_1
XFILLER_116_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08951_ _09327_/C _12447_/B _08936_/C _08936_/D vssd1 vssd1 vccd1 vccd1 _08953_/C
+ sky130_fd_sc_hd__a22oi_1
XFILLER_103_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08882_ _08882_/A _09027_/A vssd1 vssd1 vccd1 vccd1 _08889_/B sky130_fd_sc_hd__nor2_1
XFILLER_29_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_760 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09503_ _09502_/A _09362_/D _09497_/A _09361_/Y vssd1 vssd1 vccd1 vccd1 _09504_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_37_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_59 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09434_ _09434_/A _09434_/B _09434_/C vssd1 vssd1 vccd1 vccd1 _09435_/C sky130_fd_sc_hd__nand3_1
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09365_ _09497_/A _09504_/A _09497_/C vssd1 vssd1 vccd1 vccd1 _09498_/A sky130_fd_sc_hd__o21a_1
XFILLER_166_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_30 _17543_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09296_ _09296_/A _09296_/B _09296_/C vssd1 vssd1 vccd1 vccd1 _09296_/Y sky130_fd_sc_hd__nand3_1
XFILLER_123_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_41 _14772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_52 _08967_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_63 _10508_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_559 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_74 _17480_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_85 _12077_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_96 _09979_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_732 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10140_ _10140_/A _10140_/B vssd1 vssd1 vccd1 vccd1 _10148_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10071_ _10560_/B _10072_/B vssd1 vssd1 vccd1 vccd1 _10073_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13830_ _13936_/B _13830_/B vssd1 vssd1 vccd1 vccd1 _13830_/X sky130_fd_sc_hd__or2_1
XFILLER_29_974 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_911 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13761_ _13761_/A _13761_/B vssd1 vssd1 vccd1 vccd1 _13762_/B sky130_fd_sc_hd__and2_1
X_10973_ _10973_/A _10973_/B vssd1 vssd1 vccd1 vccd1 _10974_/B sky130_fd_sc_hd__nor2_1
XFILLER_16_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_955 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15500_ _15501_/A _15501_/B _15501_/C vssd1 vssd1 vccd1 vccd1 _15594_/A sky130_fd_sc_hd__o21a_1
XFILLER_16_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12712_ _12698_/Y _12699_/X _12711_/X vssd1 vssd1 vccd1 vccd1 _17581_/D sky130_fd_sc_hd__o21ai_1
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16480_ _16480_/A _16571_/B _14775_/A vssd1 vssd1 vccd1 vccd1 _16481_/B sky130_fd_sc_hd__or3b_1
X_13692_ _13693_/B _13793_/A _16796_/A vssd1 vssd1 vccd1 vccd1 _13694_/A sky130_fd_sc_hd__o21a_1
XFILLER_43_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15431_ _15431_/A _15431_/B vssd1 vssd1 vccd1 vccd1 _15433_/B sky130_fd_sc_hd__xnor2_1
X_12643_ _12642_/A _12642_/B _12642_/C vssd1 vssd1 vccd1 vccd1 _12798_/A sky130_fd_sc_hd__o21ai_1
XFILLER_15_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15362_ _15362_/A _15362_/B vssd1 vssd1 vccd1 vccd1 _15363_/B sky130_fd_sc_hd__xnor2_1
X_12574_ _12415_/A _12417_/B _12415_/B vssd1 vssd1 vccd1 vccd1 _12581_/A sky130_fd_sc_hd__o21ba_1
XFILLER_30_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17101_ _17099_/A _17100_/X _17064_/X _17067_/Y vssd1 vssd1 vccd1 vccd1 _17103_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_11_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14313_ _14381_/A _14313_/B vssd1 vssd1 vccd1 vccd1 _14315_/B sky130_fd_sc_hd__or2_1
X_11525_ _11526_/A _11525_/B _11525_/C vssd1 vssd1 vccd1 vccd1 _11526_/B sky130_fd_sc_hd__nand3_1
XFILLER_12_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_868 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15293_ _15159_/A _15159_/B _15221_/B _15226_/A _15226_/B vssd1 vssd1 vccd1 vccd1
+ _15295_/B sky130_fd_sc_hd__a32o_1
XFILLER_172_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17032_ _16735_/A _14636_/B _17164_/C _15715_/X vssd1 vssd1 vccd1 vccd1 _17033_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_116_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14244_ _14244_/A _14244_/B vssd1 vssd1 vccd1 vccd1 _14245_/C sky130_fd_sc_hd__xnor2_1
XFILLER_109_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11456_ _11456_/A _11456_/B _11456_/C vssd1 vssd1 vccd1 vccd1 _11456_/X sky130_fd_sc_hd__or3_1
XFILLER_109_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10407_ _10441_/A _10441_/B vssd1 vssd1 vccd1 vccd1 _10407_/Y sky130_fd_sc_hd__nor2_1
X_14175_ _14176_/A _14385_/B vssd1 vssd1 vccd1 vccd1 _14177_/B sky130_fd_sc_hd__nand2_1
X_11387_ _11561_/A _11387_/B _11387_/C vssd1 vssd1 vccd1 vccd1 _11393_/B sky130_fd_sc_hd__and3_1
XFILLER_125_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_927 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13126_ _12980_/X _12984_/A _13258_/A _13125_/X vssd1 vssd1 vccd1 vccd1 _13258_/B
+ sky130_fd_sc_hd__a211oi_1
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10338_ _10451_/A _10334_/B _10332_/X vssd1 vssd1 vccd1 vccd1 _10352_/A sky130_fd_sc_hd__a21o_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13057_ _13057_/A _13057_/B _13057_/C vssd1 vssd1 vccd1 vccd1 _13058_/B sky130_fd_sc_hd__nor3_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10269_ _14784_/A _10270_/B vssd1 vssd1 vccd1 vccd1 _10269_/X sky130_fd_sc_hd__and2_1
XFILLER_78_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_971 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12008_ _17405_/A _09229_/B _09230_/A _09228_/A vssd1 vssd1 vccd1 vccd1 _12009_/A
+ sky130_fd_sc_hd__a31oi_1
XFILLER_94_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16816_ _16816_/A _16888_/A _16816_/C vssd1 vssd1 vccd1 vccd1 _16818_/B sky130_fd_sc_hd__and3_1
XFILLER_94_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16747_ _16747_/A _16813_/B vssd1 vssd1 vccd1 vccd1 _16883_/C sky130_fd_sc_hd__nor2_2
X_13959_ _14044_/B _13959_/B vssd1 vssd1 vccd1 vccd1 _13961_/C sky130_fd_sc_hd__nor2_1
XFILLER_34_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16678_ _16770_/A _16678_/B vssd1 vssd1 vccd1 vccd1 _16690_/A sky130_fd_sc_hd__or2_1
XFILLER_35_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_796 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15629_ _15037_/X _15039_/X _15057_/X _15059_/Y _15312_/S _15901_/S vssd1 vssd1 vccd1
+ vccd1 _15629_/X sky130_fd_sc_hd__mux4_1
XFILLER_148_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09150_ _09150_/A _09150_/B vssd1 vssd1 vccd1 vccd1 _09153_/C sky130_fd_sc_hd__xnor2_1
XFILLER_147_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09081_ _09081_/A _09306_/A vssd1 vssd1 vccd1 vccd1 _09088_/A sky130_fd_sc_hd__nor2_1
XFILLER_163_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput50 i_wb_data[22] vssd1 vssd1 vccd1 vccd1 input50/X sky130_fd_sc_hd__clkbuf_1
XFILLER_162_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput61 i_wb_data[3] vssd1 vssd1 vccd1 vccd1 input61/X sky130_fd_sc_hd__clkbuf_2
XFILLER_174_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1003 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09983_ _09983_/A _09983_/B _09989_/B vssd1 vssd1 vccd1 vccd1 _10004_/B sky130_fd_sc_hd__or3_1
XFILLER_130_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08934_ _08937_/A vssd1 vssd1 vccd1 vccd1 _08936_/C sky130_fd_sc_hd__inv_2
XFILLER_131_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08865_ _08866_/A _08866_/B vssd1 vssd1 vccd1 vccd1 _08867_/A sky130_fd_sc_hd__and2_1
XFILLER_57_524 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08796_ _08796_/A _08796_/B vssd1 vssd1 vccd1 vccd1 _08798_/C sky130_fd_sc_hd__xor2_1
XFILLER_84_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_914 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09417_ _09417_/A _09417_/B vssd1 vssd1 vccd1 vccd1 _09546_/B sky130_fd_sc_hd__xnor2_1
XFILLER_41_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09348_ _09354_/A _09354_/B vssd1 vssd1 vccd1 vccd1 _09355_/A sky130_fd_sc_hd__nor2_1
XFILLER_166_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_170 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09279_ _09279_/A _09279_/B vssd1 vssd1 vccd1 vccd1 _09281_/B sky130_fd_sc_hd__xnor2_1
XFILLER_166_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11310_ _11285_/A _11285_/B _11285_/C vssd1 vssd1 vccd1 vccd1 _11311_/C sky130_fd_sc_hd__a21oi_1
X_12290_ _12267_/Y _12268_/X _12476_/B _12290_/D vssd1 vssd1 vccd1 vccd1 _12290_/X
+ sky130_fd_sc_hd__and4bb_2
XFILLER_113_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11241_ _11097_/C _17468_/D _11098_/A _11096_/Y vssd1 vssd1 vccd1 vccd1 _11242_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_10_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11172_ _10988_/Y _10999_/X _11202_/A _11171_/Y vssd1 vssd1 vccd1 vccd1 _11202_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_122_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10123_ _10123_/A _10123_/B vssd1 vssd1 vccd1 vccd1 _10125_/B sky130_fd_sc_hd__xnor2_1
X_15980_ _15980_/A _15980_/B _15980_/C vssd1 vssd1 vccd1 vccd1 _15981_/B sky130_fd_sc_hd__nor3_1
XFILLER_121_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14931_ _17476_/D _17477_/D _14836_/B vssd1 vssd1 vccd1 vccd1 _14931_/X sky130_fd_sc_hd__or3b_4
X_10054_ _10054_/A _10054_/B vssd1 vssd1 vccd1 vccd1 _10055_/B sky130_fd_sc_hd__nor2_1
XFILLER_121_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_844 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14862_ _16651_/A _16651_/B vssd1 vssd1 vccd1 vccd1 _16652_/B sky130_fd_sc_hd__and2_1
XFILLER_48_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_911 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16601_ _16601_/A _16601_/B vssd1 vssd1 vccd1 vccd1 _16614_/A sky130_fd_sc_hd__nand2_1
X_13813_ _13814_/A wire118/X _13814_/C vssd1 vssd1 vccd1 vccd1 _13925_/A sky130_fd_sc_hd__o21ai_1
XFILLER_63_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17581_ fanout949/X _17581_/D vssd1 vssd1 vccd1 vccd1 _17581_/Q sky130_fd_sc_hd__dfxtp_1
X_14793_ _14794_/A _15008_/A vssd1 vssd1 vccd1 vccd1 _14793_/Y sky130_fd_sc_hd__nor2_1
XFILLER_29_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16532_ _16533_/C _16695_/C vssd1 vssd1 vccd1 vccd1 _16534_/A sky130_fd_sc_hd__and2b_1
XFILLER_73_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13744_ _13852_/A _13852_/B vssd1 vssd1 vccd1 vccd1 _13853_/A sky130_fd_sc_hd__nand2_1
X_10956_ _11006_/B _17468_/D _10954_/D _10954_/A vssd1 vssd1 vccd1 vccd1 _10957_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_90_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16463_ _16557_/A _16463_/B vssd1 vssd1 vccd1 vccd1 _16466_/A sky130_fd_sc_hd__nand2b_1
XFILLER_73_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13675_ _13977_/A _13977_/B _14050_/D _13966_/D vssd1 vssd1 vccd1 vccd1 _13676_/B
+ sky130_fd_sc_hd__and4_1
X_10887_ _11651_/A _10932_/B _15206_/A _15130_/S vssd1 vssd1 vccd1 vccd1 _10888_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_31_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15414_ _15414_/A _15414_/B vssd1 vssd1 vccd1 vccd1 _15417_/A sky130_fd_sc_hd__xor2_1
X_12626_ _12626_/A _12626_/B _12626_/C vssd1 vssd1 vccd1 vccd1 _12627_/B sky130_fd_sc_hd__nand3_1
X_16394_ _16394_/A _16394_/B vssd1 vssd1 vccd1 vccd1 _16396_/B sky130_fd_sc_hd__and2_1
XFILLER_12_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15345_ _15345_/A _15345_/B vssd1 vssd1 vccd1 vccd1 _15346_/B sky130_fd_sc_hd__xnor2_1
XFILLER_8_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12557_ _12869_/A _13450_/C _13208_/C _12714_/A vssd1 vssd1 vccd1 vccd1 _12557_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_172_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11508_ _11553_/A _11629_/D _11605_/B _11427_/A vssd1 vssd1 vccd1 vccd1 _11509_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_145_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15276_ _15277_/A _15277_/B vssd1 vssd1 vccd1 vccd1 _15276_/Y sky130_fd_sc_hd__nor2_1
X_12488_ _17409_/A _12787_/D vssd1 vssd1 vccd1 vccd1 _12490_/C sky130_fd_sc_hd__nand2_1
XFILLER_156_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17015_ _17014_/A _17014_/C _17014_/B vssd1 vssd1 vccd1 vccd1 _17016_/C sky130_fd_sc_hd__a21oi_1
XFILLER_7_196 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14227_ _14227_/A _16970_/A vssd1 vssd1 vccd1 vccd1 _14229_/C sky130_fd_sc_hd__xnor2_1
X_11439_ _11440_/A _11438_/Y _11520_/C _14850_/A vssd1 vssd1 vccd1 vccd1 _11479_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_144_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14158_ _14158_/A _14158_/B _14158_/C vssd1 vssd1 vccd1 vccd1 _14159_/B sky130_fd_sc_hd__nor3_1
XFILLER_99_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13109_ _13109_/A _13109_/B vssd1 vssd1 vccd1 vccd1 _13110_/B sky130_fd_sc_hd__nand2_1
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14089_ _14176_/A _14433_/B vssd1 vssd1 vccd1 vccd1 _14090_/B sky130_fd_sc_hd__nand2_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09202_ _09202_/A _09202_/B vssd1 vssd1 vccd1 vccd1 _09208_/A sky130_fd_sc_hd__nor2_1
XFILLER_148_621 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09133_ _17536_/Q _12127_/D vssd1 vssd1 vccd1 vccd1 _09176_/A sky130_fd_sc_hd__nand2_1
XFILLER_33_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1016 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09064_ _17375_/A _12258_/B _08950_/A _08948_/Y vssd1 vssd1 vccd1 vccd1 _09065_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_162_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09966_ _09966_/A _09966_/B vssd1 vssd1 vccd1 vccd1 _09969_/C sky130_fd_sc_hd__xnor2_1
XFILLER_103_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08917_ _08918_/B _08918_/A vssd1 vssd1 vccd1 vccd1 _08917_/X sky130_fd_sc_hd__and2b_1
XFILLER_98_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09897_ _09898_/A _09898_/C vssd1 vssd1 vccd1 vccd1 _09902_/B sky130_fd_sc_hd__nor2_1
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_952 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08848_ _08846_/Y _08996_/A _09321_/C _11895_/D vssd1 vssd1 vccd1 vccd1 _08996_/B
+ sky130_fd_sc_hd__and4bb_1
XFILLER_73_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08779_ _08779_/A _08779_/B vssd1 vssd1 vccd1 vccd1 _08802_/A sky130_fd_sc_hd__xor2_1
XFILLER_84_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_77 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10810_ _11095_/B _17469_/D _17468_/D _11095_/A vssd1 vssd1 vccd1 vccd1 _10810_/Y
+ sky130_fd_sc_hd__a22oi_1
XTAP_2847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11790_ _11790_/A _16136_/A vssd1 vssd1 vccd1 vccd1 _11790_/X sky130_fd_sc_hd__or2_1
XFILLER_150_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10741_ _10742_/A _10742_/C vssd1 vssd1 vccd1 vccd1 _10747_/B sky130_fd_sc_hd__nor2_1
XFILLER_14_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_32 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13460_ _13576_/B _13460_/B vssd1 vssd1 vccd1 vccd1 _13462_/C sky130_fd_sc_hd__nand2_1
X_10672_ _10672_/A _10672_/B vssd1 vssd1 vccd1 vccd1 _10673_/B sky130_fd_sc_hd__and2_1
XFILLER_40_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12411_ _12412_/A _12412_/B vssd1 vssd1 vccd1 vccd1 _12572_/A sky130_fd_sc_hd__and2_1
XFILLER_40_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13391_ _12710_/A _13390_/X _16653_/A vssd1 vssd1 vccd1 vccd1 _13391_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_21_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15130_ _15131_/B _15129_/X _15130_/S vssd1 vssd1 vccd1 vccd1 _15130_/X sky130_fd_sc_hd__mux2_1
XFILLER_127_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12342_ _12343_/A _12343_/B _12343_/C vssd1 vssd1 vccd1 vccd1 _12344_/A sky130_fd_sc_hd__o21a_1
XFILLER_138_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15061_ _15131_/A _15061_/B vssd1 vssd1 vccd1 vccd1 _15061_/Y sky130_fd_sc_hd__nand2_1
X_12273_ _12273_/A _12273_/B vssd1 vssd1 vccd1 vccd1 _12283_/A sky130_fd_sc_hd__xnor2_1
XFILLER_4_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14012_ _14013_/A _14013_/B _14013_/C vssd1 vssd1 vccd1 vccd1 _14015_/B sky130_fd_sc_hd__a21oi_1
XFILLER_141_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11224_ _11225_/A _11225_/B vssd1 vssd1 vccd1 vccd1 _11224_/X sky130_fd_sc_hd__and2b_1
X_11155_ _11155_/A _11234_/A vssd1 vssd1 vccd1 vccd1 _11232_/B sky130_fd_sc_hd__nor2_1
XFILLER_110_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10106_ _10106_/A _10106_/B vssd1 vssd1 vccd1 vccd1 _10133_/A sky130_fd_sc_hd__xnor2_1
X_15963_ _15963_/A _15963_/B vssd1 vssd1 vccd1 vccd1 _15964_/B sky130_fd_sc_hd__xor2_1
X_11086_ _11069_/X _11070_/Y _11084_/A _11090_/A vssd1 vssd1 vccd1 vccd1 _11087_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_95_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14914_ _10014_/D _10146_/B _14914_/S vssd1 vssd1 vccd1 vccd1 _14915_/B sky130_fd_sc_hd__mux2_1
X_10037_ _10638_/B _10534_/D _10036_/D _10638_/A vssd1 vssd1 vccd1 vccd1 _10037_/Y
+ sky130_fd_sc_hd__a22oi_1
X_15894_ _15890_/X _15891_/X _15892_/Y _15893_/Y _16111_/A vssd1 vssd1 vccd1 vccd1
+ _15894_/X sky130_fd_sc_hd__a311o_1
XFILLER_48_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14845_ _15008_/A _15008_/B vssd1 vssd1 vccd1 vccd1 _14846_/B sky130_fd_sc_hd__nand2_1
XFILLER_64_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14776_ _14776_/A _16399_/A vssd1 vssd1 vccd1 vccd1 _16397_/B sky130_fd_sc_hd__or2_1
X_17564_ fanout953/X _17564_/D vssd1 vssd1 vccd1 vccd1 _17564_/Q sky130_fd_sc_hd__dfxtp_1
X_11988_ _11988_/A _11988_/B vssd1 vssd1 vccd1 vccd1 _11990_/C sky130_fd_sc_hd__xnor2_1
XFILLER_63_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16515_ _16515_/A _16515_/B vssd1 vssd1 vccd1 vccd1 _16517_/A sky130_fd_sc_hd__nand2_1
XFILLER_56_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13727_ _13727_/A _13727_/B vssd1 vssd1 vccd1 vccd1 _13936_/A sky130_fd_sc_hd__or2_1
X_10939_ _10940_/A _10940_/B vssd1 vssd1 vccd1 vccd1 _10990_/B sky130_fd_sc_hd__nand2_1
XFILLER_16_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17495_ fanout945/X _17495_/D vssd1 vssd1 vccd1 vccd1 _17495_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16446_ _16446_/A _16619_/A _16681_/C _16681_/D vssd1 vssd1 vccd1 vccd1 _16446_/X
+ sky130_fd_sc_hd__or4_1
X_13658_ _13658_/A _13852_/B _13658_/C vssd1 vssd1 vccd1 vccd1 _13659_/B sky130_fd_sc_hd__and3_1
XPHY_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12609_ _12610_/A _12610_/B vssd1 vssd1 vccd1 vccd1 _12778_/B sky130_fd_sc_hd__or2_1
X_16377_ _16378_/B _16378_/A vssd1 vssd1 vccd1 vccd1 _16470_/B sky130_fd_sc_hd__nand2b_1
XFILLER_9_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13589_ _13589_/A _13589_/B vssd1 vssd1 vccd1 vccd1 _13592_/A sky130_fd_sc_hd__xor2_1
XFILLER_76_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15328_ _14899_/X _14968_/X _16619_/A _11675_/B vssd1 vssd1 vccd1 vccd1 _15404_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_172_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15259_ _15233_/X _15234_/Y _15258_/X vssd1 vssd1 vccd1 vccd1 _15259_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_117_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout407 _14774_/A vssd1 vssd1 vccd1 vccd1 _12714_/A sky130_fd_sc_hd__buf_2
X_09820_ _09524_/A _09523_/B _09523_/A vssd1 vssd1 vccd1 vccd1 _09827_/A sky130_fd_sc_hd__o21ba_1
Xfanout418 _17529_/Q vssd1 vssd1 vccd1 vccd1 _12070_/A sky130_fd_sc_hd__buf_4
XFILLER_63_1028 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout429 _17528_/Q vssd1 vssd1 vccd1 vccd1 _10109_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_86_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09751_ _09751_/A _09880_/A vssd1 vssd1 vccd1 vccd1 _09758_/A sky130_fd_sc_hd__nor2_1
XFILLER_113_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09682_ _09674_/B _09670_/X _09631_/Y _09666_/B vssd1 vssd1 vccd1 vccd1 _09819_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_104_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09116_ _09119_/B _09119_/C vssd1 vssd1 vccd1 vccd1 _09257_/A sky130_fd_sc_hd__nand2_1
XFILLER_159_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09047_ _09047_/A _09047_/B vssd1 vssd1 vccd1 vccd1 _09049_/B sky130_fd_sc_hd__xnor2_1
XFILLER_159_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_852 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout930 _17358_/C1 vssd1 vssd1 vccd1 vccd1 _17420_/C1 sky130_fd_sc_hd__clkbuf_2
XFILLER_131_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout941 fanout957/X vssd1 vssd1 vccd1 vccd1 fanout941/X sky130_fd_sc_hd__buf_2
Xfanout952 fanout953/X vssd1 vssd1 vccd1 vccd1 fanout952/X sky130_fd_sc_hd__clkbuf_2
X_09949_ _10321_/B _10203_/B _10061_/B vssd1 vssd1 vccd1 vccd1 _09951_/C sky130_fd_sc_hd__and3_1
XFILLER_77_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12960_ _12960_/A _12960_/B vssd1 vssd1 vccd1 vccd1 _12979_/A sky130_fd_sc_hd__and2_1
XTAP_3301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11911_ _11911_/A _11911_/B _11911_/C vssd1 vssd1 vccd1 vccd1 _11911_/Y sky130_fd_sc_hd__nand3_1
XFILLER_85_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_88 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12891_ _12889_/Y _13043_/A _13302_/A _13035_/C vssd1 vssd1 vccd1 vccd1 _13043_/B
+ sky130_fd_sc_hd__and4bb_1
XFILLER_79_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14630_ _14585_/A _14582_/A _14584_/B vssd1 vssd1 vccd1 vccd1 _14631_/B sky130_fd_sc_hd__a21oi_1
XTAP_2644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11842_ _10897_/C _11841_/X _12046_/A vssd1 vssd1 vccd1 vccd1 _11842_/Y sky130_fd_sc_hd__o21ai_2
XTAP_3389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14561_ _14562_/A _14562_/B _14562_/C vssd1 vssd1 vccd1 vccd1 _14612_/A sky130_fd_sc_hd__a21o_1
XTAP_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11773_ _11773_/A _11773_/B vssd1 vssd1 vccd1 vccd1 _17105_/B sky130_fd_sc_hd__and2_1
XTAP_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13512_ _13010_/B _13511_/X _13510_/X vssd1 vssd1 vccd1 vccd1 _13514_/B sky130_fd_sc_hd__a21oi_1
XTAP_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16300_ _16300_/A _16300_/B vssd1 vssd1 vccd1 vccd1 _16301_/B sky130_fd_sc_hd__nor2_1
X_10724_ _10724_/A _10724_/B vssd1 vssd1 vccd1 vccd1 _11174_/B sky130_fd_sc_hd__nor2_1
X_17280_ _17570_/Q _17292_/B vssd1 vssd1 vccd1 vccd1 _17280_/X sky130_fd_sc_hd__and2_1
XTAP_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14492_ _14492_/A _14492_/B vssd1 vssd1 vccd1 vccd1 _14493_/C sky130_fd_sc_hd__xor2_1
XTAP_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16231_ _16232_/A _16232_/B vssd1 vssd1 vccd1 vccd1 _16231_/Y sky130_fd_sc_hd__nand2_1
XFILLER_13_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13443_ _13443_/A _13443_/B _13443_/C vssd1 vssd1 vccd1 vccd1 _13444_/A sky130_fd_sc_hd__and3_1
XFILLER_174_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10655_ _10655_/A _10655_/B vssd1 vssd1 vccd1 vccd1 _10661_/A sky130_fd_sc_hd__nor2_1
XFILLER_173_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16162_ _16068_/A _16068_/B _16069_/Y vssd1 vssd1 vccd1 vccd1 _16179_/A sky130_fd_sc_hd__a21bo_1
XFILLER_70_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13374_ _13494_/A _13373_/B _13496_/B _13373_/D vssd1 vssd1 vccd1 vccd1 _13374_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_154_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10586_ _10586_/A _10586_/B vssd1 vssd1 vccd1 vccd1 _10681_/A sky130_fd_sc_hd__xnor2_1
XFILLER_6_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15113_ _16731_/B1 _14848_/C _15110_/Y _15112_/Y _15109_/X vssd1 vssd1 vccd1 vccd1
+ _15113_/X sky130_fd_sc_hd__o311a_1
XFILLER_155_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12325_ _12325_/A _12325_/B _12325_/C vssd1 vssd1 vccd1 vccd1 _12327_/A sky130_fd_sc_hd__or3_1
XFILLER_115_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16093_ _15981_/B _15983_/B _15979_/Y vssd1 vssd1 vccd1 vccd1 _16095_/B sky130_fd_sc_hd__o21a_1
XFILLER_142_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15044_ _15041_/X _15042_/X _15043_/X vssd1 vssd1 vccd1 vccd1 _15044_/Y sky130_fd_sc_hd__a21oi_1
X_12256_ _13035_/A _12734_/B _12256_/C _12256_/D vssd1 vssd1 vccd1 vccd1 _12257_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_123_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11207_ _11175_/Y _11178_/Y _11206_/Y _10761_/A vssd1 vssd1 vccd1 vccd1 _11719_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_141_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12187_ _12188_/A _12188_/B vssd1 vssd1 vccd1 vccd1 _12189_/A sky130_fd_sc_hd__nand2_1
XFILLER_122_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11138_ _11293_/A _11138_/B vssd1 vssd1 vccd1 vccd1 _11139_/C sky130_fd_sc_hd__and2_1
X_16995_ _16996_/B _16995_/B vssd1 vssd1 vccd1 vccd1 _16997_/A sky130_fd_sc_hd__and2b_1
XFILLER_77_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15946_ _16880_/A _16054_/B vssd1 vssd1 vccd1 vccd1 _16533_/B sky130_fd_sc_hd__and2_2
X_11069_ _11069_/A _11069_/B _11069_/C vssd1 vssd1 vccd1 vccd1 _11069_/X sky130_fd_sc_hd__or3_1
XFILLER_23_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15877_ _15877_/A _15877_/B _15875_/Y vssd1 vssd1 vccd1 vccd1 _15878_/B sky130_fd_sc_hd__or3b_1
XFILLER_110_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_143 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14828_ _14492_/A _14826_/X _14827_/Y _14597_/B vssd1 vssd1 vccd1 vccd1 _14828_/Y
+ sky130_fd_sc_hd__a211oi_2
XFILLER_64_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_571 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17547_ fanout938/X _17547_/D vssd1 vssd1 vccd1 vccd1 _17547_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14759_ _14755_/A _14755_/B _14751_/A vssd1 vssd1 vccd1 vccd1 _14762_/A sky130_fd_sc_hd__o21a_1
XFILLER_44_390 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17478_ fanout949/X _17478_/D vssd1 vssd1 vccd1 vccd1 _17478_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_149_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16429_ _16747_/A _16514_/A _16938_/B _16681_/A vssd1 vssd1 vccd1 vccd1 _16431_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_20_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_763 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout204 _11849_/Y vssd1 vssd1 vccd1 vccd1 _16219_/A1 sky130_fd_sc_hd__buf_2
XFILLER_8_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout226 _14933_/Y vssd1 vssd1 vccd1 vccd1 _16799_/B1 sky130_fd_sc_hd__clkbuf_2
XFILLER_101_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09803_ _10560_/A _10072_/B _09803_/C vssd1 vssd1 vccd1 vccd1 _09939_/A sky130_fd_sc_hd__and3_1
Xfanout237 _16401_/C1 vssd1 vssd1 vccd1 vccd1 _17170_/B1 sky130_fd_sc_hd__clkbuf_4
XFILLER_115_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_170 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout248 _16007_/A vssd1 vssd1 vccd1 vccd1 _16304_/A sky130_fd_sc_hd__clkbuf_4
Xfanout259 _11783_/Y vssd1 vssd1 vccd1 vccd1 _16106_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_59_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09734_ _09894_/C _10543_/B _09607_/A _09605_/Y vssd1 vssd1 vccd1 vccd1 _09735_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_27_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09665_ _09665_/A _09665_/B vssd1 vssd1 vccd1 vccd1 _09666_/B sky130_fd_sc_hd__nand2_1
XFILLER_39_195 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09596_ _09596_/A _09596_/B vssd1 vssd1 vccd1 vccd1 _09686_/B sky130_fd_sc_hd__xnor2_1
XFILLER_70_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_922 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10440_ _10440_/A _10453_/B vssd1 vssd1 vccd1 vccd1 _10473_/A sky130_fd_sc_hd__nand2_1
XFILLER_148_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10371_ _10383_/B _10383_/C _10383_/A vssd1 vssd1 vccd1 vccd1 _10385_/A sky130_fd_sc_hd__a21o_1
XFILLER_40_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12110_ _12110_/A _12110_/B vssd1 vssd1 vccd1 vccd1 _12113_/A sky130_fd_sc_hd__xnor2_1
XFILLER_108_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13090_ _13220_/B _13090_/B vssd1 vssd1 vccd1 vccd1 _13092_/C sky130_fd_sc_hd__nand2_1
XFILLER_2_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1023 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12041_ _12463_/D _12295_/D _14942_/A vssd1 vssd1 vccd1 vccd1 _12042_/B sky130_fd_sc_hd__mux2_1
XFILLER_2_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout760 _17493_/Q vssd1 vssd1 vccd1 vccd1 _10036_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_120_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout771 fanout772/X vssd1 vssd1 vccd1 vccd1 _10532_/D sky130_fd_sc_hd__buf_4
X_15800_ _15797_/Y _15798_/Y _15799_/Y vssd1 vssd1 vccd1 vccd1 _15800_/Y sky130_fd_sc_hd__o21ai_1
Xfanout782 _10743_/C vssd1 vssd1 vccd1 vccd1 _10146_/B sky130_fd_sc_hd__clkbuf_4
X_16780_ _16781_/A _16781_/B vssd1 vssd1 vccd1 vccd1 _16846_/B sky130_fd_sc_hd__nor2_1
X_13992_ _14167_/A _14865_/B vssd1 vssd1 vccd1 vccd1 _14080_/C sky130_fd_sc_hd__and2_2
Xfanout793 fanout795/X vssd1 vssd1 vccd1 vccd1 _10743_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_59_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15731_ _15732_/A _15732_/B vssd1 vssd1 vccd1 vccd1 _15731_/X sky130_fd_sc_hd__or2_1
X_12943_ _13897_/A _13080_/C vssd1 vssd1 vccd1 vccd1 _12945_/C sky130_fd_sc_hd__nand2_1
XFILLER_74_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12874_ _12875_/B _12875_/A vssd1 vssd1 vccd1 vccd1 _13033_/A sky130_fd_sc_hd__nand2b_1
XFILLER_46_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15662_ _15750_/A _16065_/B vssd1 vssd1 vccd1 vccd1 _15663_/B sky130_fd_sc_hd__nand2_1
XTAP_3186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17401_ _17401_/A _17421_/B vssd1 vssd1 vccd1 vccd1 _17401_/X sky130_fd_sc_hd__or2_1
XTAP_2463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14613_ _14567_/A _14567_/B _14566_/A vssd1 vssd1 vccd1 vccd1 _14615_/B sky130_fd_sc_hd__a21oi_1
X_11825_ _12054_/A _15238_/A _11595_/A vssd1 vssd1 vccd1 vccd1 _11826_/B sky130_fd_sc_hd__a21bo_1
X_15593_ _15594_/A _15594_/B vssd1 vssd1 vccd1 vccd1 _15595_/A sky130_fd_sc_hd__nand2_1
XTAP_2474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_80 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17332_ _09042_/B _17356_/A2 _17331_/X _17422_/C1 vssd1 vssd1 vccd1 vccd1 _17495_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14544_ _14641_/B _14593_/D _14545_/D _14641_/A vssd1 vssd1 vccd1 vccd1 _14548_/A
+ sky130_fd_sc_hd__a22oi_1
X_11756_ _11756_/A _11756_/B vssd1 vssd1 vccd1 vccd1 _16568_/B sky130_fd_sc_hd__xor2_2
XFILLER_53_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10707_ _10708_/B _10708_/A vssd1 vssd1 vccd1 vccd1 _10715_/B sky130_fd_sc_hd__nand2b_1
XFILLER_41_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14475_ _14475_/A vssd1 vssd1 vccd1 vccd1 _14533_/C sky130_fd_sc_hd__inv_2
X_17263_ _17455_/Q _17290_/A2 _17261_/X _17262_/X _17293_/C1 vssd1 vssd1 vccd1 vccd1
+ _17455_/D sky130_fd_sc_hd__o221a_1
XFILLER_174_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11687_ _11688_/A _11688_/B vssd1 vssd1 vccd1 vccd1 _11692_/B sky130_fd_sc_hd__nand2_1
XFILLER_146_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13426_ _13421_/Y _13422_/X _13308_/A _13309_/B vssd1 vssd1 vccd1 vccd1 _13428_/B
+ sky130_fd_sc_hd__o211a_1
X_16214_ _08760_/Y _14778_/X _14813_/X vssd1 vssd1 vccd1 vccd1 _16214_/Y sky130_fd_sc_hd__a21oi_1
X_10638_ _10638_/A _10638_/B _10933_/D _10970_/B vssd1 vssd1 vccd1 vccd1 _10641_/A
+ sky130_fd_sc_hd__and4_1
X_17194_ input6/X input11/X input13/X input12/X vssd1 vssd1 vccd1 vccd1 _17195_/C
+ sky130_fd_sc_hd__or4_1
XFILLER_139_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16145_ _16146_/B _16146_/A vssd1 vssd1 vccd1 vccd1 _16145_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_154_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13357_ _13357_/A _13357_/B vssd1 vssd1 vccd1 vccd1 _13360_/A sky130_fd_sc_hd__xnor2_1
X_10569_ _10672_/A _10569_/B vssd1 vssd1 vccd1 vccd1 _10572_/B sky130_fd_sc_hd__and2_1
XFILLER_155_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12308_ _12309_/A _12309_/B _12309_/C vssd1 vssd1 vccd1 vccd1 _12310_/A sky130_fd_sc_hd__a21oi_1
XFILLER_143_958 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16076_ _16077_/A _16077_/B vssd1 vssd1 vccd1 vccd1 _16183_/B sky130_fd_sc_hd__and2_1
XFILLER_170_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13288_ _13286_/Y _13417_/A _13643_/A _13738_/B vssd1 vssd1 vccd1 vccd1 _13417_/B
+ sky130_fd_sc_hd__and4bb_1
X_15027_ _15024_/Y _15025_/Y _11518_/A vssd1 vssd1 vccd1 vccd1 _15687_/A sky130_fd_sc_hd__o21ai_4
XFILLER_142_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12239_ _12239_/A _12239_/B vssd1 vssd1 vccd1 vccd1 _12241_/B sky130_fd_sc_hd__nor2_1
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16978_ _17140_/A _17028_/B _16973_/Y _16977_/X vssd1 vssd1 vccd1 vccd1 _16978_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_37_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput4 i_wb_addr[10] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__clkbuf_1
XFILLER_110_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15929_ _15726_/A _16127_/A _16743_/C _17043_/B _15821_/X vssd1 vssd1 vccd1 vccd1
+ _15937_/A sky130_fd_sc_hd__a41o_1
XFILLER_36_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09450_ _09321_/C _09321_/D _09328_/A _09320_/Y vssd1 vssd1 vccd1 vccd1 _09451_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_65_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09381_ _09381_/A _09381_/B vssd1 vssd1 vccd1 vccd1 _09382_/C sky130_fd_sc_hd__xnor2_1
XFILLER_17_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_582 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_791 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09717_ _09717_/A _09717_/B vssd1 vssd1 vccd1 vccd1 _09719_/B sky130_fd_sc_hd__xnor2_1
XFILLER_28_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09648_ _10559_/A _09843_/C _09647_/C vssd1 vssd1 vccd1 vccd1 _09649_/B sky130_fd_sc_hd__a21oi_1
XFILLER_55_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09579_ _09579_/A _09579_/B vssd1 vssd1 vccd1 vccd1 _09581_/C sky130_fd_sc_hd__or2_1
XFILLER_31_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11610_ _11610_/A _11610_/B vssd1 vssd1 vccd1 vccd1 _11611_/B sky130_fd_sc_hd__nand2_1
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12590_ _12592_/B _12592_/C _12592_/D _12592_/A vssd1 vssd1 vccd1 vccd1 _12593_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_143_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11541_ _11541_/A _11542_/A _11541_/C vssd1 vssd1 vccd1 vccd1 _11584_/A sky130_fd_sc_hd__nor3_1
XFILLER_23_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14260_ _14257_/Y _14258_/X _14164_/X _14186_/A vssd1 vssd1 vccd1 vccd1 _14262_/C
+ sky130_fd_sc_hd__a211oi_1
XFILLER_109_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11472_ _11472_/A _11472_/B _11471_/X vssd1 vssd1 vccd1 vccd1 _11512_/A sky130_fd_sc_hd__or3b_1
XFILLER_149_590 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13211_ _13211_/A _13339_/A _13211_/C vssd1 vssd1 vccd1 vccd1 _13339_/B sky130_fd_sc_hd__nor3_1
X_10423_ _10423_/A _10423_/B vssd1 vssd1 vccd1 vccd1 _10524_/B sky130_fd_sc_hd__xnor2_1
X_14191_ _14192_/A _14192_/B _14192_/C vssd1 vssd1 vccd1 vccd1 _14270_/A sky130_fd_sc_hd__a21o_1
XFILLER_137_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13142_ _13627_/S _12047_/X _12063_/C _12858_/Y vssd1 vssd1 vccd1 vccd1 _13142_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_100_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10354_ _10330_/B _10319_/C _10319_/D _10319_/A vssd1 vssd1 vccd1 vccd1 _10354_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_151_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13073_ _13244_/A _13073_/B vssd1 vssd1 vccd1 vccd1 _13075_/C sky130_fd_sc_hd__nor2_1
XFILLER_97_308 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_500 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10285_ _10188_/A _10188_/B _10188_/C vssd1 vssd1 vccd1 vccd1 _10285_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_105_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16901_ _16900_/A _16900_/B _16900_/C vssd1 vssd1 vccd1 vccd1 _16902_/B sky130_fd_sc_hd__a21oi_1
XFILLER_78_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12024_ _14952_/A _14949_/B _14912_/B vssd1 vssd1 vccd1 vccd1 _12024_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_2_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16832_ _16832_/A _16832_/B vssd1 vssd1 vccd1 vccd1 _16897_/B sky130_fd_sc_hd__nor2_1
XFILLER_93_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout590 _17512_/Q vssd1 vssd1 vccd1 vccd1 _11518_/A sky130_fd_sc_hd__buf_4
XFILLER_93_536 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16763_ _16764_/B _16763_/B vssd1 vssd1 vccd1 vccd1 _16765_/A sky130_fd_sc_hd__and2b_1
XFILLER_47_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13975_ _13867_/A _13869_/B _13867_/B vssd1 vssd1 vccd1 vccd1 _13982_/A sky130_fd_sc_hd__o21ba_1
XFILLER_58_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15714_ _10145_/B _15804_/A2 _15713_/X vssd1 vssd1 vccd1 vccd1 _15714_/Y sky130_fd_sc_hd__a21oi_1
X_12926_ _12926_/A _12926_/B vssd1 vssd1 vccd1 vccd1 _12928_/C sky130_fd_sc_hd__xnor2_1
XFILLER_62_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16694_ _16777_/A _16694_/B vssd1 vssd1 vccd1 vccd1 _16701_/A sky130_fd_sc_hd__nand2_1
XFILLER_18_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_411 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15645_ _15734_/A _15645_/B _16514_/A vssd1 vssd1 vccd1 vccd1 _15645_/Y sky130_fd_sc_hd__nor3_1
XFILLER_62_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12857_ _12382_/X _12398_/X _16011_/B vssd1 vssd1 vccd1 vccd1 _12857_/X sky130_fd_sc_hd__mux2_1
XTAP_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_308 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11808_ _17363_/A _11808_/B vssd1 vssd1 vccd1 vccd1 _14982_/C sky130_fd_sc_hd__and2_1
X_15576_ _15393_/B _15205_/B _15617_/A vssd1 vssd1 vccd1 vccd1 _16883_/A sky130_fd_sc_hd__a21bo_1
X_12788_ _12788_/A _13080_/D vssd1 vssd1 vccd1 vccd1 _12790_/C sky130_fd_sc_hd__nand2_1
XTAP_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17315_ input67/X _17321_/B _17321_/C vssd1 vssd1 vccd1 vccd1 _17315_/X sky130_fd_sc_hd__or3_1
XFILLER_147_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11739_ _11739_/A _11739_/B _11739_/C vssd1 vssd1 vccd1 vccd1 _11753_/A sky130_fd_sc_hd__or3_1
X_14527_ _14528_/A _14528_/B vssd1 vssd1 vccd1 vccd1 _14583_/B sky130_fd_sc_hd__or2_1
XFILLER_159_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17246_ _17591_/Q _17291_/A2 _17291_/B1 vssd1 vssd1 vccd1 vccd1 _17246_/X sky130_fd_sc_hd__a21o_1
X_14458_ _14528_/A _14458_/B vssd1 vssd1 vccd1 vccd1 _14459_/C sky130_fd_sc_hd__and2_1
X_13409_ _13409_/A _13409_/B vssd1 vssd1 vccd1 vccd1 _13411_/C sky130_fd_sc_hd__xor2_1
XFILLER_143_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17177_ input30/X input32/X input31/X input34/X vssd1 vssd1 vccd1 vccd1 _17180_/B
+ sky130_fd_sc_hd__or4_1
X_14389_ _14389_/A _14389_/B vssd1 vssd1 vccd1 vccd1 _14456_/B sky130_fd_sc_hd__or2_1
XFILLER_116_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16128_ _16807_/A _16127_/X _16126_/X vssd1 vssd1 vccd1 vccd1 _16130_/A sky130_fd_sc_hd__a21o_1
XFILLER_115_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_755 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_468 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08950_ _08950_/A _09065_/A vssd1 vssd1 vccd1 vccd1 _08959_/A sky130_fd_sc_hd__nor2_1
X_16059_ _16165_/A _16533_/B vssd1 vssd1 vccd1 vccd1 _16060_/B sky130_fd_sc_hd__nand2_1
X_08881_ _08882_/A _08880_/Y _17401_/A _12340_/B vssd1 vssd1 vccd1 vccd1 _09027_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_97_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09502_ _09502_/A _09502_/B _09502_/C vssd1 vssd1 vccd1 vccd1 _09786_/A sky130_fd_sc_hd__and3_1
XFILLER_65_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_720 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09433_ _09433_/A _09433_/B vssd1 vssd1 vccd1 vccd1 _09435_/B sky130_fd_sc_hd__xnor2_1
XFILLER_64_282 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09364_ _09364_/A _09364_/B vssd1 vssd1 vccd1 vccd1 _09497_/C sky130_fd_sc_hd__nor2_1
XFILLER_21_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_20 _17575_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09295_ _09296_/A _09296_/B _09296_/C vssd1 vssd1 vccd1 vccd1 _09316_/A sky130_fd_sc_hd__a21o_2
XANTENNA_31 _17544_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_302 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_42 _14772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_53 _14765_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_64 _12338_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_75 _17510_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_86 _10638_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_97 _17480_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10070_ _10070_/A _10070_/B vssd1 vssd1 vccd1 vccd1 _10073_/A sky130_fd_sc_hd__and2_1
XFILLER_0_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13760_ _13761_/A _13761_/B vssd1 vssd1 vccd1 vccd1 _13762_/A sky130_fd_sc_hd__nor2_1
XFILLER_29_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10972_ _11115_/B _10971_/B _14806_/A vssd1 vssd1 vccd1 vccd1 _10973_/B sky130_fd_sc_hd__a21oi_1
XFILLER_44_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_496 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12711_ _11849_/A _12707_/X _12710_/X _16735_/A vssd1 vssd1 vccd1 vccd1 _12711_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_44_967 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13691_ _14167_/A _13893_/A _13691_/C _16651_/A vssd1 vssd1 vccd1 vccd1 _13793_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_102_60 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12642_ _12642_/A _12642_/B _12642_/C vssd1 vssd1 vccd1 vccd1 _12644_/A sky130_fd_sc_hd__or3_1
X_15430_ _16281_/A _16505_/A vssd1 vssd1 vccd1 vccd1 _15431_/B sky130_fd_sc_hd__nand2_1
XFILLER_31_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15361_ _15362_/B _15362_/A vssd1 vssd1 vccd1 vccd1 _15361_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_129_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12573_ _12425_/A _12427_/B _12425_/B vssd1 vssd1 vccd1 vccd1 _12583_/A sky130_fd_sc_hd__o21ba_1
XFILLER_23_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17100_ _14867_/A _17134_/C _17100_/C vssd1 vssd1 vccd1 vccd1 _17100_/X sky130_fd_sc_hd__and3b_1
X_11524_ _11514_/A _11514_/C _11558_/A vssd1 vssd1 vccd1 vccd1 _11525_/C sky130_fd_sc_hd__o21ai_1
XFILLER_129_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14312_ _14312_/A _14312_/B vssd1 vssd1 vccd1 vccd1 _14313_/B sky130_fd_sc_hd__and2_1
XFILLER_7_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15292_ _15292_/A _15292_/B vssd1 vssd1 vccd1 vccd1 _15295_/A sky130_fd_sc_hd__xnor2_1
XFILLER_168_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14243_ _14387_/A _14385_/B vssd1 vssd1 vccd1 vccd1 _14244_/B sky130_fd_sc_hd__nand2_1
X_17031_ _17023_/A _17163_/A2 _17030_/X vssd1 vssd1 vccd1 vccd1 _17033_/C sky130_fd_sc_hd__o21ba_1
X_11455_ _11451_/A _11451_/B _11495_/A vssd1 vssd1 vccd1 vccd1 _11456_/C sky130_fd_sc_hd__o21ba_1
X_10406_ _10405_/A _10406_/B vssd1 vssd1 vccd1 vccd1 _10441_/B sky130_fd_sc_hd__and2b_1
X_14174_ _14252_/A _14174_/B vssd1 vssd1 vccd1 vccd1 _14177_/A sky130_fd_sc_hd__and2_1
X_11386_ _11386_/A _11386_/B vssd1 vssd1 vccd1 vccd1 _11393_/A sky130_fd_sc_hd__xnor2_1
XFILLER_152_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13125_ _13125_/A _13125_/B _13125_/C vssd1 vssd1 vccd1 vccd1 _13125_/X sky130_fd_sc_hd__and3_1
X_10337_ _10336_/A _10336_/Y _10215_/B _10228_/Y vssd1 vssd1 vccd1 vccd1 _10337_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_97_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13056_ _13057_/A _13057_/B _13057_/C vssd1 vssd1 vccd1 vccd1 _13199_/A sky130_fd_sc_hd__o21a_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10268_ _10268_/A _10268_/B vssd1 vssd1 vccd1 vccd1 _10276_/A sky130_fd_sc_hd__xnor2_1
XFILLER_87_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12007_ _12007_/A _12007_/B vssd1 vssd1 vccd1 vccd1 _12010_/A sky130_fd_sc_hd__xor2_1
XFILLER_39_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10199_ _10321_/B _10067_/B _10067_/C vssd1 vssd1 vccd1 vccd1 _10200_/B sky130_fd_sc_hd__a21oi_1
X_16815_ _16021_/A _16589_/B _16813_/Y vssd1 vssd1 vccd1 vccd1 _16816_/C sky130_fd_sc_hd__a21o_1
X_16746_ _16746_/A _16746_/B vssd1 vssd1 vccd1 vccd1 _16750_/A sky130_fd_sc_hd__xnor2_1
X_13958_ _13958_/A _13958_/B _13958_/C vssd1 vssd1 vccd1 vccd1 _13959_/B sky130_fd_sc_hd__nor3_1
XFILLER_46_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12909_ _12910_/A _12910_/B _12910_/C vssd1 vssd1 vccd1 vccd1 _13060_/A sky130_fd_sc_hd__o21ai_1
X_16677_ _16676_/B _16677_/B vssd1 vssd1 vccd1 vccd1 _16678_/B sky130_fd_sc_hd__and2b_1
XFILLER_34_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13889_ _13990_/A _13889_/B vssd1 vssd1 vccd1 vccd1 _13891_/B sky130_fd_sc_hd__nor2_1
XFILLER_22_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15628_ _15628_/A _15628_/B vssd1 vssd1 vccd1 vccd1 _15628_/X sky130_fd_sc_hd__and2_1
XFILLER_21_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15559_ _15559_/A _15559_/B vssd1 vssd1 vccd1 vccd1 _15675_/A sky130_fd_sc_hd__nand2_1
XFILLER_147_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09080_ _09081_/A _09079_/Y _17375_/A _11900_/D vssd1 vssd1 vccd1 vccd1 _09306_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_148_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput40 i_wb_data[13] vssd1 vssd1 vccd1 vccd1 input40/X sky130_fd_sc_hd__clkbuf_1
X_17229_ _17553_/Q _17244_/B vssd1 vssd1 vccd1 vccd1 _17229_/X sky130_fd_sc_hd__and2_1
XFILLER_162_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput51 i_wb_data[23] vssd1 vssd1 vccd1 vccd1 input51/X sky130_fd_sc_hd__clkbuf_1
XFILLER_174_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput62 i_wb_data[4] vssd1 vssd1 vccd1 vccd1 input62/X sky130_fd_sc_hd__clkbuf_2
XFILLER_116_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09982_ _09982_/A _10113_/A vssd1 vssd1 vccd1 vccd1 _09989_/B sky130_fd_sc_hd__nor2_1
XFILLER_103_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08933_ _09755_/A _09325_/B _12445_/C _12445_/D vssd1 vssd1 vccd1 vccd1 _08937_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_103_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08864_ _08864_/A _08864_/B vssd1 vssd1 vccd1 vccd1 _08866_/B sky130_fd_sc_hd__xnor2_1
XFILLER_123_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_536 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08795_ _08796_/A _08796_/B vssd1 vssd1 vccd1 vccd1 _11911_/A sky130_fd_sc_hd__nand2_1
XFILLER_84_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_926 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09416_ _16983_/A _09416_/B vssd1 vssd1 vccd1 vccd1 _09546_/A sky130_fd_sc_hd__xnor2_1
X_09347_ _09654_/C _09350_/B _09161_/Y _09163_/B vssd1 vssd1 vccd1 vccd1 _09354_/B
+ sky130_fd_sc_hd__a22oi_1
XFILLER_139_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09278_ _16982_/A _09273_/A _09273_/B vssd1 vssd1 vccd1 vccd1 _09281_/A sky130_fd_sc_hd__o21ba_1
XFILLER_21_694 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1014 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11240_ _15262_/B _15472_/A _11240_/C _17466_/D vssd1 vssd1 vccd1 vccd1 _11306_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_5_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11171_ _11168_/Y _11169_/X _11021_/X _11041_/A vssd1 vssd1 vccd1 vccd1 _11171_/Y
+ sky130_fd_sc_hd__o211ai_1
XFILLER_106_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10122_ _10116_/A _10118_/B _10116_/B vssd1 vssd1 vccd1 vccd1 _10125_/A sky130_fd_sc_hd__o21ba_1
XFILLER_164_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14930_ _17476_/D _17477_/D _14836_/B vssd1 vssd1 vccd1 vccd1 _14930_/Y sky130_fd_sc_hd__nor3b_1
XFILLER_48_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10053_ _10053_/A _10053_/B _10053_/C vssd1 vssd1 vccd1 vccd1 _10054_/B sky130_fd_sc_hd__and3_1
XFILLER_57_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14861_ _16571_/A _16480_/A _16400_/B vssd1 vssd1 vccd1 vccd1 _16651_/B sky130_fd_sc_hd__and3_1
XFILLER_29_750 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16600_ _16600_/A _16600_/B vssd1 vssd1 vccd1 vccd1 _16601_/B sky130_fd_sc_hd__or2_1
X_13812_ _13812_/A _13812_/B vssd1 vssd1 vccd1 vccd1 _13814_/C sky130_fd_sc_hd__xor2_1
XFILLER_63_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17580_ fanout937/X _17580_/D vssd1 vssd1 vccd1 vccd1 _17580_/Q sky130_fd_sc_hd__dfxtp_1
X_14792_ _15126_/A _15042_/B vssd1 vssd1 vccd1 vccd1 _14796_/B sky130_fd_sc_hd__or2_1
X_16531_ _16533_/A _16533_/B vssd1 vssd1 vccd1 vccd1 _16695_/C sky130_fd_sc_hd__nand2_1
XFILLER_16_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10955_ _11010_/A vssd1 vssd1 vccd1 vccd1 _10955_/Y sky130_fd_sc_hd__inv_2
X_13743_ _13745_/B _13852_/B _13844_/C _13852_/A vssd1 vssd1 vccd1 vccd1 _13746_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_71_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16462_ _16462_/A _16462_/B _16460_/Y vssd1 vssd1 vccd1 vccd1 _16463_/B sky130_fd_sc_hd__or3b_1
XFILLER_31_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10886_ _11281_/A _11132_/C vssd1 vssd1 vccd1 vccd1 _11131_/A sky130_fd_sc_hd__nand2_1
X_13674_ _13977_/B _14050_/D _13966_/D _13977_/A vssd1 vssd1 vccd1 vccd1 _13676_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_31_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15413_ _16056_/A _16812_/A vssd1 vssd1 vccd1 vccd1 _15414_/B sky130_fd_sc_hd__nand2_1
X_12625_ _12626_/A _12626_/B _12626_/C vssd1 vssd1 vccd1 vccd1 _12820_/A sky130_fd_sc_hd__a21o_1
X_16393_ _16300_/A _16300_/B _16299_/B vssd1 vssd1 vccd1 vccd1 _16394_/B sky130_fd_sc_hd__o21ai_1
XFILLER_40_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12556_ _12871_/A _13334_/C vssd1 vssd1 vccd1 vccd1 _12560_/A sky130_fd_sc_hd__nand2_4
X_15344_ _15750_/A _16505_/A vssd1 vssd1 vccd1 vccd1 _15345_/B sky130_fd_sc_hd__nand2_1
XFILLER_129_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11507_ _11553_/A _15008_/A _11605_/B _11427_/A vssd1 vssd1 vccd1 vccd1 _11507_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_144_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12487_ _12487_/A _12787_/B _12637_/D _12487_/D vssd1 vssd1 vccd1 vccd1 _12642_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_89_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15275_ _14881_/X _14889_/X _16595_/A _15275_/C1 vssd1 vssd1 vccd1 vccd1 _15277_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_171_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17014_ _17014_/A _17014_/B _17014_/C vssd1 vssd1 vccd1 vccd1 _17016_/B sky130_fd_sc_hd__and3_1
X_11438_ _11518_/B _14895_/B _11518_/C _11518_/A vssd1 vssd1 vccd1 vccd1 _11438_/Y
+ sky130_fd_sc_hd__a22oi_1
X_14226_ _14554_/A _14301_/C vssd1 vssd1 vccd1 vccd1 _16970_/A sky130_fd_sc_hd__nand2_4
XFILLER_125_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14157_ _14158_/A _14158_/B _14158_/C vssd1 vssd1 vccd1 vccd1 _14159_/A sky130_fd_sc_hd__o21a_1
X_11369_ _11369_/A _11369_/B vssd1 vssd1 vccd1 vccd1 _11395_/A sky130_fd_sc_hd__xnor2_1
XFILLER_99_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13108_ _13109_/A _13109_/B vssd1 vssd1 vccd1 vccd1 _13241_/A sky130_fd_sc_hd__or2_1
XFILLER_98_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14088_ _14088_/A _14088_/B vssd1 vssd1 vccd1 vccd1 _14090_/A sky130_fd_sc_hd__nand2_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13039_ _13040_/A _13040_/B _13040_/C vssd1 vssd1 vccd1 vccd1 _13181_/A sky130_fd_sc_hd__o21ai_1
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16729_ _13459_/A _16729_/B vssd1 vssd1 vccd1 vccd1 _16730_/B sky130_fd_sc_hd__nand2b_1
XFILLER_50_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09201_ _09639_/C _12338_/D _09196_/B _09193_/Y vssd1 vssd1 vccd1 vccd1 _09202_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_22_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09132_ _09360_/A _09172_/A _11920_/D _09362_/D vssd1 vssd1 vccd1 vccd1 _09135_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_148_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09063_ _09063_/A _09063_/B vssd1 vssd1 vccd1 vccd1 _09293_/A sky130_fd_sc_hd__xnor2_1
XFILLER_108_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09965_ _09966_/B _09966_/A vssd1 vssd1 vccd1 vccd1 _09968_/B sky130_fd_sc_hd__and2b_1
XFILLER_104_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08916_ _08916_/A _09057_/A vssd1 vssd1 vccd1 vccd1 _08918_/B sky130_fd_sc_hd__nor2_1
XFILLER_103_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09896_ _15538_/A _14863_/B _09890_/A _09756_/Y vssd1 vssd1 vccd1 vccd1 _09898_/C
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08847_ _09078_/A _11895_/B _11902_/B _08860_/B vssd1 vssd1 vccd1 vccd1 _08996_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_100_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08778_ _17393_/A _09042_/B vssd1 vssd1 vccd1 vccd1 _08779_/B sky130_fd_sc_hd__nand2_1
XTAP_2815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10740_ _10745_/C _10647_/D _10648_/A _10646_/Y vssd1 vssd1 vccd1 vccd1 _10742_/C
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_159_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10671_ _10671_/A _10671_/B vssd1 vssd1 vccd1 vccd1 _10672_/B sky130_fd_sc_hd__nand2_1
XFILLER_159_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12410_ _12871_/A _13208_/D _12238_/A _12236_/B vssd1 vssd1 vccd1 vccd1 _12412_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_43_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_66 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_992 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13390_ _12384_/X _12400_/B _17164_/A vssd1 vssd1 vccd1 vccd1 _13390_/X sky130_fd_sc_hd__mux2_1
XFILLER_139_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_452 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12341_ _12341_/A _12341_/B vssd1 vssd1 vccd1 vccd1 _12343_/C sky130_fd_sc_hd__xnor2_1
XFILLER_127_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_327 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15060_ _15314_/A _14850_/A _15463_/A _15541_/A _14942_/A _15095_/B vssd1 vssd1 vccd1
+ vccd1 _15061_/B sky130_fd_sc_hd__mux4_1
XFILLER_154_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12272_ _12442_/A _12592_/D vssd1 vssd1 vccd1 vccd1 _12273_/B sky130_fd_sc_hd__nand2_1
XFILLER_135_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14011_ _14011_/A _14011_/B vssd1 vssd1 vccd1 vccd1 _14013_/C sky130_fd_sc_hd__xnor2_1
X_11223_ _11223_/A _11223_/B vssd1 vssd1 vccd1 vccd1 _11225_/B sky130_fd_sc_hd__xor2_1
XFILLER_5_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11154_ _11154_/A _11155_/A _11154_/C vssd1 vssd1 vccd1 vccd1 _11234_/A sky130_fd_sc_hd__nor3_1
XFILLER_1_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10105_ _10005_/A _10005_/C _10005_/B vssd1 vssd1 vccd1 vccd1 _10105_/Y sky130_fd_sc_hd__a21oi_1
X_15962_ _15963_/A _15963_/B vssd1 vssd1 vccd1 vccd1 _15962_/Y sky130_fd_sc_hd__nor2_1
X_11085_ _11084_/A _11090_/A _11069_/X _11070_/Y vssd1 vssd1 vccd1 vccd1 _11087_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_68_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14913_ _12054_/A _10016_/D _10991_/C vssd1 vssd1 vccd1 vccd1 _14913_/Y sky130_fd_sc_hd__a21oi_1
X_10036_ _10638_/A _10638_/B _10534_/D _10036_/D vssd1 vssd1 vccd1 vccd1 _10039_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_75_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15893_ _15890_/X _15891_/X _15892_/Y vssd1 vssd1 vccd1 vccd1 _15893_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_75_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14844_ _14929_/A _14938_/B vssd1 vssd1 vccd1 vccd1 _14844_/X sky130_fd_sc_hd__or2_1
XFILLER_64_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17563_ fanout952/X _17563_/D vssd1 vssd1 vccd1 vccd1 _17563_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14775_ _14775_/A _16480_/A vssd1 vssd1 vccd1 vccd1 _14775_/X sky130_fd_sc_hd__or2_1
X_11987_ _11987_/A _11987_/B vssd1 vssd1 vccd1 vccd1 _11988_/B sky130_fd_sc_hd__nor2_1
XFILLER_32_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16514_ _16514_/A _16938_/B _16514_/C vssd1 vssd1 vccd1 vccd1 _16515_/B sky130_fd_sc_hd__or3_1
XFILLER_44_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13726_ _13726_/A _13726_/B vssd1 vssd1 vccd1 vccd1 _13727_/B sky130_fd_sc_hd__and2_1
X_10938_ _10938_/A _10938_/B vssd1 vssd1 vccd1 vccd1 _10940_/B sky130_fd_sc_hd__xor2_1
X_17494_ fanout943/X _17494_/D vssd1 vssd1 vccd1 vccd1 _17494_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16445_ _16619_/A _16681_/D vssd1 vssd1 vccd1 vccd1 _16533_/C sky130_fd_sc_hd__nor2_1
XFILLER_31_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10869_ _11115_/B _11117_/D _11115_/C _11115_/A vssd1 vssd1 vccd1 vccd1 _10870_/B
+ sky130_fd_sc_hd__a22oi_1
X_13657_ _13541_/A _13657_/B vssd1 vssd1 vccd1 vccd1 _13658_/C sky130_fd_sc_hd__nand2b_1
XPHY_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12608_ _12778_/A _12608_/B vssd1 vssd1 vccd1 vccd1 _12610_/B sky130_fd_sc_hd__nand2_1
X_16376_ _16280_/B _16282_/B _16280_/A vssd1 vssd1 vccd1 vccd1 _16378_/B sky130_fd_sc_hd__o21ba_1
XPHY_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13588_ _13469_/A _13471_/B _13469_/B vssd1 vssd1 vccd1 vccd1 _13589_/B sky130_fd_sc_hd__o21ba_1
XFILLER_129_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15327_ _14882_/X _15325_/X _17377_/A vssd1 vssd1 vccd1 vccd1 _16168_/A sky130_fd_sc_hd__a21o_2
XFILLER_8_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12539_ _12540_/A _12540_/B vssd1 vssd1 vccd1 vccd1 _12539_/Y sky130_fd_sc_hd__nor2_1
XFILLER_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15258_ _16389_/A _15235_/Y _15236_/X _15257_/X vssd1 vssd1 vccd1 vccd1 _15258_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_173_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14209_ _12388_/X _12401_/B _14356_/S vssd1 vssd1 vccd1 vccd1 _14209_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15189_ _15131_/A _14921_/X _16011_/B vssd1 vssd1 vccd1 vccd1 _15189_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_99_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout408 _17530_/Q vssd1 vssd1 vccd1 vccd1 _14774_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_140_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout419 _17529_/Q vssd1 vssd1 vccd1 vccd1 _10366_/A sky130_fd_sc_hd__buf_2
XFILLER_141_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09750_ _09751_/A _09749_/Y _09894_/C _10545_/D vssd1 vssd1 vccd1 vccd1 _09880_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_39_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_940 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09681_ _09681_/A _09681_/B vssd1 vssd1 vccd1 vccd1 _09825_/A sky130_fd_sc_hd__or2_1
XFILLER_66_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_612 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09115_ _09115_/A _09115_/B _09115_/C vssd1 vssd1 vccd1 vccd1 _09119_/C sky130_fd_sc_hd__or3_1
XFILLER_164_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09046_ _09047_/B _09047_/A vssd1 vssd1 vccd1 vccd1 _09055_/B sky130_fd_sc_hd__nand2b_1
XFILLER_163_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout920 _17171_/X vssd1 vssd1 vccd1 vccd1 _17245_/A2 sky130_fd_sc_hd__clkbuf_4
Xfanout931 _17378_/C1 vssd1 vssd1 vccd1 vccd1 _17358_/C1 sky130_fd_sc_hd__clkbuf_4
Xfanout942 fanout948/X vssd1 vssd1 vccd1 vccd1 fanout942/X sky130_fd_sc_hd__buf_2
X_09948_ _09948_/A _09948_/B vssd1 vssd1 vccd1 vccd1 _10061_/B sky130_fd_sc_hd__xnor2_1
XFILLER_89_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout953 fanout954/X vssd1 vssd1 vccd1 vccd1 fanout953/X sky130_fd_sc_hd__clkbuf_2
XFILLER_57_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09879_ _09894_/C _10545_/D _09751_/A _09749_/Y vssd1 vssd1 vccd1 vccd1 _09880_/B
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_3302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11910_ _11911_/A _11911_/B _11911_/C vssd1 vssd1 vccd1 vccd1 _12148_/A sky130_fd_sc_hd__a21o_1
XFILLER_46_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12890_ _13658_/A _13414_/B _13908_/B _13802_/B vssd1 vssd1 vccd1 vccd1 _13043_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_85_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11841_ _17363_/A _11841_/B vssd1 vssd1 vccd1 vccd1 _11841_/X sky130_fd_sc_hd__and2_1
XTAP_2645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14560_ _14560_/A _14560_/B vssd1 vssd1 vccd1 vccd1 _14562_/C sky130_fd_sc_hd__xor2_1
X_11772_ _11771_/A _16972_/A _16972_/B _11770_/Y vssd1 vssd1 vccd1 vccd1 _11773_/B
+ sky130_fd_sc_hd__a31o_1
XTAP_2689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10723_ _11117_/C _10743_/D _10641_/A _10639_/Y vssd1 vssd1 vccd1 vccd1 _10724_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_13511_ _13511_/A _13511_/B vssd1 vssd1 vccd1 vccd1 _13511_/X sky130_fd_sc_hd__and2_1
XTAP_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14491_ _14599_/B _14641_/C vssd1 vssd1 vccd1 vccd1 _14492_/B sky130_fd_sc_hd__nand2_1
XTAP_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16230_ _16126_/X _16130_/B _16127_/X _16807_/A vssd1 vssd1 vccd1 vccd1 _16232_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_13_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13442_ _13442_/A _13442_/B vssd1 vssd1 vccd1 vccd1 _13443_/C sky130_fd_sc_hd__xnor2_1
XFILLER_16_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10654_ _10545_/C _10657_/B _10546_/A _10544_/Y vssd1 vssd1 vccd1 vccd1 _10655_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_139_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16161_ _16161_/A _16161_/B vssd1 vssd1 vccd1 vccd1 _16181_/A sky130_fd_sc_hd__xnor2_1
X_13373_ _13494_/A _13373_/B _13496_/B _13373_/D vssd1 vssd1 vccd1 vccd1 _13494_/B
+ sky130_fd_sc_hd__nor4_1
XFILLER_154_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10585_ _10573_/X _10574_/Y _10567_/A _10572_/A vssd1 vssd1 vccd1 vccd1 _10585_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_103_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15112_ _14791_/X _16008_/A2 _15111_/X _14944_/A vssd1 vssd1 vccd1 vccd1 _15112_/Y
+ sky130_fd_sc_hd__a211oi_1
X_12324_ _12324_/A _12492_/B vssd1 vssd1 vccd1 vccd1 _12325_/C sky130_fd_sc_hd__nor2_1
X_16092_ _16092_/A _16092_/B vssd1 vssd1 vccd1 vccd1 _16095_/A sky130_fd_sc_hd__xnor2_2
XFILLER_6_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12255_ _12734_/B _12256_/C _12256_/D _13035_/A vssd1 vssd1 vccd1 vccd1 _12257_/A
+ sky130_fd_sc_hd__a22oi_1
X_15043_ _14941_/X _15003_/X _15002_/X vssd1 vssd1 vccd1 vccd1 _15043_/X sky130_fd_sc_hd__a21bo_1
XFILLER_119_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11206_ _10760_/A _10760_/B _10760_/C vssd1 vssd1 vccd1 vccd1 _11206_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_107_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12186_ _12186_/A _12186_/B vssd1 vssd1 vccd1 vccd1 _12188_/B sky130_fd_sc_hd__xor2_1
X_11137_ _11137_/A _11137_/B _11137_/C vssd1 vssd1 vccd1 vccd1 _11138_/B sky130_fd_sc_hd__or3_1
XFILLER_123_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16994_ _16994_/A _16994_/B vssd1 vssd1 vccd1 vccd1 _16995_/B sky130_fd_sc_hd__and2_1
XFILLER_122_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11068_ _11055_/X _11056_/Y _11065_/B _11065_/Y vssd1 vssd1 vccd1 vccd1 _11069_/C
+ sky130_fd_sc_hd__o211a_1
X_15945_ _15859_/A _15859_/B _15857_/X vssd1 vssd1 vccd1 vccd1 _15969_/A sky130_fd_sc_hd__o21ai_1
XFILLER_37_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10019_ _10019_/A _10019_/B vssd1 vssd1 vccd1 vccd1 _10136_/A sky130_fd_sc_hd__xnor2_1
X_15876_ _15877_/A _15877_/B _15875_/Y vssd1 vssd1 vccd1 vccd1 _15992_/A sky130_fd_sc_hd__o21ba_1
XFILLER_64_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14827_ _17100_/C _14867_/A vssd1 vssd1 vccd1 vccd1 _14827_/Y sky130_fd_sc_hd__nor2_1
XFILLER_63_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17546_ fanout956/X _17546_/D vssd1 vssd1 vccd1 vccd1 _17546_/Q sky130_fd_sc_hd__dfxtp_4
X_14758_ _14758_/A _14758_/B vssd1 vssd1 vccd1 vccd1 _14758_/Y sky130_fd_sc_hd__nor2_1
X_13709_ _13706_/Y _13707_/X _13594_/X _13598_/A vssd1 vssd1 vccd1 vccd1 _13710_/D
+ sky130_fd_sc_hd__a211oi_1
X_17477_ fanout956/X _17477_/D vssd1 vssd1 vccd1 vccd1 _17477_/Q sky130_fd_sc_hd__dfxtp_1
X_14689_ _14717_/A _14689_/B vssd1 vssd1 vccd1 vccd1 _14691_/B sky130_fd_sc_hd__nand2_1
X_16428_ _16324_/A _16326_/B _16324_/B vssd1 vssd1 vccd1 vccd1 _16436_/A sky130_fd_sc_hd__a21bo_1
XFILLER_149_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16359_ _16443_/A _16359_/B vssd1 vssd1 vccd1 vccd1 _16361_/B sky130_fd_sc_hd__and2_1
XFILLER_146_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout205 _12046_/A vssd1 vssd1 vccd1 vccd1 _11837_/A sky130_fd_sc_hd__buf_2
Xfanout216 _16591_/B vssd1 vssd1 vccd1 vccd1 _16935_/B sky130_fd_sc_hd__buf_2
Xfanout227 _16008_/B1 vssd1 vssd1 vccd1 vccd1 _15713_/B1 sky130_fd_sc_hd__buf_2
XFILLER_8_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09802_ _09805_/B _09802_/B vssd1 vssd1 vccd1 vccd1 _09803_/C sky130_fd_sc_hd__nor2_1
XFILLER_87_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout238 _16401_/C1 vssd1 vssd1 vccd1 vccd1 _16806_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout249 _15456_/B vssd1 vssd1 vccd1 vccd1 _16007_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_87_759 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09733_ _09733_/A _09733_/B vssd1 vssd1 vccd1 vccd1 _09867_/A sky130_fd_sc_hd__xnor2_1
XFILLER_68_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09664_ _09665_/A _09665_/B vssd1 vssd1 vccd1 vccd1 _09666_/A sky130_fd_sc_hd__or2_1
XFILLER_54_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09595_ _09597_/A _09597_/B vssd1 vssd1 vccd1 vccd1 _09686_/A sky130_fd_sc_hd__nand2_1
XFILLER_82_453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_934 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10370_ _10709_/A _10370_/B _10370_/C vssd1 vssd1 vccd1 vccd1 _10383_/C sky130_fd_sc_hd__or3_1
XFILLER_156_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09029_ _17395_/A _09030_/C _11961_/B _17397_/A vssd1 vssd1 vccd1 vccd1 _09031_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_151_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12040_ _14912_/B _12040_/B vssd1 vssd1 vccd1 vccd1 _12040_/Y sky130_fd_sc_hd__nand2_1
XFILLER_46_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout750 _12942_/D vssd1 vssd1 vccd1 vccd1 _13664_/D sky130_fd_sc_hd__buf_2
XFILLER_49_98 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout761 fanout772/X vssd1 vssd1 vccd1 vccd1 _13551_/D sky130_fd_sc_hd__buf_2
XFILLER_77_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout772 _17492_/Q vssd1 vssd1 vccd1 vccd1 fanout772/X sky130_fd_sc_hd__clkbuf_8
X_13991_ _14318_/B _14485_/D _14426_/D _14318_/A vssd1 vssd1 vccd1 vccd1 _13991_/X
+ sky130_fd_sc_hd__a22o_1
Xfanout783 _17491_/Q vssd1 vssd1 vccd1 vccd1 _10743_/C sky130_fd_sc_hd__buf_4
XFILLER_46_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout794 fanout795/X vssd1 vssd1 vccd1 vccd1 _10014_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_93_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15730_ _15730_/A _15730_/B vssd1 vssd1 vccd1 vccd1 _15732_/B sky130_fd_sc_hd__xnor2_1
XFILLER_19_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12942_ _13080_/A _13450_/B _14778_/B _12942_/D vssd1 vssd1 vccd1 vccd1 _13085_/A
+ sky130_fd_sc_hd__and4_1
XTAP_3132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15661_ _15661_/A _15661_/B vssd1 vssd1 vccd1 vccd1 _15663_/A sky130_fd_sc_hd__xnor2_1
X_12873_ _12715_/A _12717_/B _12715_/B vssd1 vssd1 vccd1 vccd1 _12875_/B sky130_fd_sc_hd__o21ba_1
XTAP_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17400_ input45/X _17422_/A2 _17399_/X _17422_/C1 vssd1 vssd1 vccd1 vccd1 _17528_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14612_ _14612_/A _14612_/B vssd1 vssd1 vccd1 vccd1 _14614_/B sky130_fd_sc_hd__xnor2_1
XTAP_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_114 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11824_ _11837_/A _11824_/B vssd1 vssd1 vccd1 vccd1 _11824_/Y sky130_fd_sc_hd__nand2_1
XTAP_2464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15592_ _15750_/A _16812_/A _15498_/A _15496_/A vssd1 vssd1 vccd1 vccd1 _15594_/B
+ sky130_fd_sc_hd__a31o_1
XTAP_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17331_ input44/X _17355_/B _17355_/C vssd1 vssd1 vccd1 vccd1 _17331_/X sky130_fd_sc_hd__or3_1
XTAP_2497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14543_ _16653_/A _14543_/B vssd1 vssd1 vccd1 vccd1 _14543_/Y sky130_fd_sc_hd__nand2_1
XTAP_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11755_ _11759_/A _11755_/B vssd1 vssd1 vccd1 vccd1 _11756_/B sky130_fd_sc_hd__and2b_1
XTAP_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10706_ _11030_/A _10705_/B _10705_/A vssd1 vssd1 vccd1 vccd1 _10708_/B sky130_fd_sc_hd__o21ba_1
X_17262_ _17564_/Q _17289_/B vssd1 vssd1 vccd1 vccd1 _17262_/X sky130_fd_sc_hd__and2_1
X_14474_ _14473_/A _14473_/B _14473_/C vssd1 vssd1 vccd1 vccd1 _14475_/A sky130_fd_sc_hd__a21oi_1
X_11686_ _11686_/A _11686_/B vssd1 vssd1 vccd1 vccd1 _11688_/B sky130_fd_sc_hd__xnor2_1
XFILLER_174_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16213_ _16107_/Y _16111_/B _16210_/Y _16917_/A vssd1 vssd1 vccd1 vccd1 _16213_/X
+ sky130_fd_sc_hd__o31a_1
X_13425_ _13428_/A vssd1 vssd1 vccd1 vccd1 _13425_/Y sky130_fd_sc_hd__inv_2
X_10637_ _10637_/A _10637_/B vssd1 vssd1 vccd1 vccd1 _10653_/A sky130_fd_sc_hd__xnor2_1
X_17193_ input32/X input31/X input33/X input7/X vssd1 vssd1 vccd1 vccd1 _17195_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_10_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16144_ _16035_/A _16035_/B _16027_/Y vssd1 vssd1 vccd1 vccd1 _16146_/B sky130_fd_sc_hd__o21a_1
XFILLER_6_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13356_ _13357_/A _13357_/B vssd1 vssd1 vccd1 vccd1 _13477_/A sky130_fd_sc_hd__and2b_1
X_10568_ _10672_/A _10569_/B vssd1 vssd1 vccd1 vccd1 _10572_/A sky130_fd_sc_hd__nor2_2
XFILLER_128_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_251 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12307_ _12307_/A _12307_/B vssd1 vssd1 vccd1 vccd1 _12309_/C sky130_fd_sc_hd__xnor2_1
X_16075_ _16075_/A _16075_/B vssd1 vssd1 vccd1 vccd1 _16077_/B sky130_fd_sc_hd__xnor2_1
X_10499_ _10499_/A vssd1 vssd1 vccd1 vccd1 _10499_/Y sky130_fd_sc_hd__inv_2
X_13287_ _13852_/A _13745_/B _13735_/D _13632_/D vssd1 vssd1 vccd1 vccd1 _13417_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_108_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15026_ _15024_/Y _15025_/Y _11518_/A vssd1 vssd1 vccd1 vccd1 _15088_/B sky130_fd_sc_hd__o21a_1
X_12238_ _12238_/A _12238_/B vssd1 vssd1 vccd1 vccd1 _12241_/A sky130_fd_sc_hd__xnor2_1
XFILLER_69_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12169_ _12169_/A _12169_/B _12169_/C vssd1 vssd1 vccd1 vccd1 _12170_/B sky130_fd_sc_hd__and3_1
XFILLER_69_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16977_ _16977_/A _16977_/B _16977_/C vssd1 vssd1 vccd1 vccd1 _16977_/X sky130_fd_sc_hd__and3_1
XFILLER_96_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput5 i_wb_addr[11] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__clkbuf_1
XFILLER_65_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15928_ _15832_/A _15829_/X _15831_/B vssd1 vssd1 vccd1 vccd1 _15939_/A sky130_fd_sc_hd__o21ai_1
XFILLER_92_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15859_ _15859_/A _15859_/B vssd1 vssd1 vccd1 vccd1 _15861_/B sky130_fd_sc_hd__xor2_1
XFILLER_149_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09380_ _09381_/B _09381_/A vssd1 vssd1 vccd1 vccd1 _09383_/A sky130_fd_sc_hd__and2b_1
XFILLER_80_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17529_ fanout945/X _17529_/D vssd1 vssd1 vccd1 vccd1 _17529_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_720 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1046 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09716_ _09717_/B _09717_/A vssd1 vssd1 vccd1 vccd1 _09725_/B sky130_fd_sc_hd__nand2b_1
XFILLER_27_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_902 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09647_ _10559_/A _09843_/C _09647_/C vssd1 vssd1 vccd1 vccd1 _09969_/B sky130_fd_sc_hd__and3_1
XFILLER_76_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09578_ _09578_/A _09578_/B vssd1 vssd1 vccd1 vccd1 _09579_/B sky130_fd_sc_hd__nor2_1
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_812 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11540_ _11539_/A _11539_/B _11538_/X vssd1 vssd1 vccd1 vccd1 _11541_/C sky130_fd_sc_hd__o21ba_1
XFILLER_169_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11471_ _11506_/B _15042_/B _11468_/D _11506_/A vssd1 vssd1 vccd1 vccd1 _11471_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_167_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10422_ _10422_/A _10531_/A vssd1 vssd1 vccd1 vccd1 _10524_/A sky130_fd_sc_hd__or2_1
XFILLER_13_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13210_ _13211_/A _13339_/A _13211_/C vssd1 vssd1 vccd1 vccd1 _13212_/A sky130_fd_sc_hd__o21a_1
XFILLER_167_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_904 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14190_ _14190_/A _14190_/B vssd1 vssd1 vccd1 vccd1 _14192_/C sky130_fd_sc_hd__xnor2_1
XFILLER_152_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13141_ _16922_/A _13139_/X _13140_/Y _13013_/Y _13016_/X vssd1 vssd1 vccd1 vccd1
+ _17584_/D sky130_fd_sc_hd__a32o_1
X_10353_ _10336_/A _10336_/C _10336_/B vssd1 vssd1 vccd1 vccd1 _10353_/X sky130_fd_sc_hd__o21a_1
X_13072_ _13072_/A _13072_/B _13072_/C vssd1 vssd1 vccd1 vccd1 _13073_/B sky130_fd_sc_hd__nor3_1
XFILLER_3_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10284_ _10263_/X _10283_/X _10157_/Y _10230_/X vssd1 vssd1 vccd1 vccd1 _10319_/A
+ sky130_fd_sc_hd__o211ai_4
X_16900_ _16900_/A _16900_/B _16900_/C vssd1 vssd1 vccd1 vccd1 _16902_/A sky130_fd_sc_hd__and3_1
XFILLER_78_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12023_ _12025_/A _14864_/A vssd1 vssd1 vccd1 vccd1 _14949_/B sky130_fd_sc_hd__and2_1
XFILLER_78_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16831_ _16832_/A _16832_/B vssd1 vssd1 vccd1 vccd1 _16833_/A sky130_fd_sc_hd__and2_1
XFILLER_66_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout580 _10180_/A vssd1 vssd1 vccd1 vccd1 _12845_/S sky130_fd_sc_hd__clkbuf_4
Xfanout591 _12700_/B vssd1 vssd1 vccd1 vccd1 _09654_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_76_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16762_ _16762_/A _16762_/B vssd1 vssd1 vccd1 vccd1 _16763_/B sky130_fd_sc_hd__xor2_1
XFILLER_76_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13974_ _13974_/A _13974_/B vssd1 vssd1 vccd1 vccd1 _14016_/A sky130_fd_sc_hd__xnor2_1
XFILLER_58_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15713_ _15707_/B _16008_/A2 _15713_/B1 _15709_/A _14944_/A vssd1 vssd1 vccd1 vccd1
+ _15713_/X sky130_fd_sc_hd__a221o_1
X_12925_ _13069_/A _13194_/D vssd1 vssd1 vccd1 vccd1 _12926_/B sky130_fd_sc_hd__nand2_1
X_16693_ _16692_/B _16693_/B vssd1 vssd1 vccd1 vccd1 _16694_/B sky130_fd_sc_hd__nand2b_1
XFILLER_20_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15644_ _16129_/A _16604_/B _16758_/B _15918_/A vssd1 vssd1 vccd1 vccd1 _15644_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_61_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12856_ _12856_/A _12856_/B vssd1 vssd1 vccd1 vccd1 _17582_/D sky130_fd_sc_hd__nand2_1
XTAP_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11807_ _11837_/A _11807_/B vssd1 vssd1 vccd1 vccd1 _11807_/Y sky130_fd_sc_hd__nand2_1
XTAP_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15575_ _15393_/B _15205_/B _15617_/A vssd1 vssd1 vccd1 vccd1 _15575_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_33_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12787_ _13080_/A _12787_/B _12942_/D _12787_/D vssd1 vssd1 vccd1 vccd1 _12947_/A
+ sky130_fd_sc_hd__and4_1
XTAP_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17314_ _12338_/D _17322_/A2 _17313_/X _17388_/C1 vssd1 vssd1 vccd1 vccd1 _17486_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_42_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14526_ _14583_/A _14526_/B vssd1 vssd1 vccd1 vccd1 _14528_/B sky130_fd_sc_hd__nand2_1
X_11738_ _11736_/A _11736_/B _11735_/Y vssd1 vssd1 vccd1 vccd1 _11739_/C sky130_fd_sc_hd__o21ba_1
X_17245_ _17449_/Q _17245_/A2 _17243_/X _17244_/X _17284_/C1 vssd1 vssd1 vccd1 vccd1
+ _17449_/D sky130_fd_sc_hd__o221a_1
X_14457_ _14456_/A _14456_/B _14456_/C vssd1 vssd1 vccd1 vccd1 _14458_/B sky130_fd_sc_hd__a21o_1
X_11669_ _15524_/C _11670_/C vssd1 vssd1 vccd1 vccd1 _11690_/B sky130_fd_sc_hd__and2b_1
X_13408_ _13408_/A _13408_/B vssd1 vssd1 vccd1 vccd1 _13409_/B sky130_fd_sc_hd__xnor2_1
X_17176_ input33/X input5/X input4/X input7/X vssd1 vssd1 vccd1 vccd1 _17180_/A sky130_fd_sc_hd__or4_1
XFILLER_128_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14388_ _14388_/A _14388_/B vssd1 vssd1 vccd1 vccd1 _14456_/A sky130_fd_sc_hd__xnor2_1
XFILLER_155_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16127_ _16127_/A _16226_/C _17119_/C vssd1 vssd1 vccd1 vccd1 _16127_/X sky130_fd_sc_hd__and3_1
XFILLER_116_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13339_ _13339_/A _13339_/B _13339_/C vssd1 vssd1 vccd1 vccd1 _13341_/A sky130_fd_sc_hd__or3_1
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16058_ _16058_/A _16058_/B vssd1 vssd1 vccd1 vccd1 _16060_/A sky130_fd_sc_hd__nor2_1
XFILLER_88_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15009_ _15248_/C _14846_/B _15008_/X _16008_/B1 _15008_/A vssd1 vssd1 vccd1 vccd1
+ _15009_/X sky130_fd_sc_hd__a32o_1
XFILLER_69_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08880_ _17399_/A _09272_/D _12338_/C _12068_/A vssd1 vssd1 vccd1 vccd1 _08880_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_97_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09501_ _09502_/A _17478_/Q vssd1 vssd1 vccd1 vccd1 _10074_/A sky130_fd_sc_hd__nand2_1
XFILLER_53_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09432_ _09433_/B _09433_/A vssd1 vssd1 vccd1 vccd1 _09441_/B sky130_fd_sc_hd__nand2b_1
XFILLER_80_732 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09363_ _09502_/A _10067_/B _09357_/A _09174_/Y vssd1 vssd1 vccd1 vccd1 _09364_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_52_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09294_ _09294_/A _09294_/B vssd1 vssd1 vccd1 vccd1 _09296_/C sky130_fd_sc_hd__or2_1
XANTENNA_10 _17428_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_21 _17502_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_32 _17545_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_43 _09412_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_54 fanout699/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_65 _09265_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_76 _13142_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_358 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_87 _14863_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_98 _16935_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10971_ _11115_/B _10971_/B _14806_/A vssd1 vssd1 vccd1 vccd1 _10973_/A sky130_fd_sc_hd__and3_1
XFILLER_28_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_423 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12710_ _12710_/A _12710_/B vssd1 vssd1 vccd1 vccd1 _12710_/X sky130_fd_sc_hd__or2_1
X_13690_ _13893_/A _13691_/C _16651_/A _14167_/A vssd1 vssd1 vccd1 vccd1 _13693_/B
+ sky130_fd_sc_hd__a22oi_1
XFILLER_44_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12641_ _12641_/A _12792_/B vssd1 vssd1 vccd1 vccd1 _12642_/C sky130_fd_sc_hd__nor2_1
XFILLER_70_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15360_ _15292_/A _15292_/B _15286_/Y vssd1 vssd1 vccd1 vccd1 _15362_/B sky130_fd_sc_hd__a21oi_1
XFILLER_168_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12572_ _12572_/A _12572_/B _12572_/C vssd1 vssd1 vccd1 vccd1 _12585_/B sky130_fd_sc_hd__or3_1
XFILLER_157_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14311_ _14312_/A _14312_/B vssd1 vssd1 vccd1 vccd1 _14381_/A sky130_fd_sc_hd__nor2_1
X_11523_ _11523_/A _11523_/B vssd1 vssd1 vccd1 vccd1 _11525_/B sky130_fd_sc_hd__xnor2_1
XFILLER_8_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15291_ _15291_/A _15291_/B vssd1 vssd1 vccd1 vccd1 _15292_/B sky130_fd_sc_hd__xnor2_1
XFILLER_7_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17030_ _17023_/B _17162_/A2 _16974_/B _17028_/A _17162_/C1 vssd1 vssd1 vccd1 vccd1
+ _17030_/X sky130_fd_sc_hd__a221o_1
XFILLER_7_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14242_ _14242_/A _14242_/B vssd1 vssd1 vccd1 vccd1 _14244_/A sky130_fd_sc_hd__nor2_1
X_11454_ _11460_/A _11454_/B vssd1 vssd1 vccd1 vccd1 _11456_/B sky130_fd_sc_hd__nand2_1
XFILLER_137_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10405_ _10405_/A _10405_/B _10405_/C _10405_/D vssd1 vssd1 vccd1 vccd1 _10406_/B
+ sky130_fd_sc_hd__or4_1
X_11385_ _11395_/B _11435_/A _11395_/A vssd1 vssd1 vccd1 vccd1 _11396_/A sky130_fd_sc_hd__a21o_1
X_14173_ _14173_/A _14173_/B _14173_/C vssd1 vssd1 vccd1 vccd1 _14174_/B sky130_fd_sc_hd__or3_1
XFILLER_109_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13124_ _13125_/A _13125_/B _13125_/C vssd1 vssd1 vccd1 vccd1 _13258_/A sky130_fd_sc_hd__a21oi_2
XFILLER_11_91 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10336_ _10336_/A _10336_/B _10336_/C vssd1 vssd1 vccd1 vccd1 _10336_/Y sky130_fd_sc_hd__nor3_2
XFILLER_3_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13055_ _13055_/A _13055_/B vssd1 vssd1 vccd1 vccd1 _13057_/C sky130_fd_sc_hd__xor2_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10267_ _10267_/A _10267_/B _10267_/C vssd1 vssd1 vccd1 vccd1 _10267_/Y sky130_fd_sc_hd__nand3_1
XFILLER_112_439 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12006_ _12007_/A _12007_/B vssd1 vssd1 vccd1 vccd1 _12006_/X sky130_fd_sc_hd__and2_1
XFILLER_39_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10198_ _10198_/A _10322_/A _10198_/C vssd1 vssd1 vccd1 vccd1 _10202_/A sky130_fd_sc_hd__or3_1
XFILLER_66_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_995 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16814_ _16814_/A _16814_/B _16938_/D _16883_/C vssd1 vssd1 vccd1 vccd1 _16888_/A
+ sky130_fd_sc_hd__or4b_1
XFILLER_93_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16745_ _16745_/A _16935_/B vssd1 vssd1 vccd1 vccd1 _16746_/B sky130_fd_sc_hd__nand2_1
X_13957_ _13958_/A _13958_/B _13958_/C vssd1 vssd1 vccd1 vccd1 _14044_/B sky130_fd_sc_hd__o21a_1
XFILLER_19_475 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_272 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12908_ _12908_/A _12908_/B vssd1 vssd1 vccd1 vccd1 _12910_/C sky130_fd_sc_hd__xnor2_1
X_16676_ _16677_/B _16676_/B vssd1 vssd1 vccd1 vccd1 _16770_/A sky130_fd_sc_hd__and2b_1
X_13888_ _13888_/A _13888_/B vssd1 vssd1 vccd1 vccd1 _13889_/B sky130_fd_sc_hd__and2_1
XFILLER_50_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15627_ _16011_/A _15627_/B vssd1 vssd1 vccd1 vccd1 _15628_/B sky130_fd_sc_hd__or2_1
X_12839_ _12689_/A _12691_/A _13001_/B _12837_/Y vssd1 vssd1 vccd1 vccd1 _12840_/B
+ sky130_fd_sc_hd__o211ai_1
XTAP_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15558_ _15559_/A _15559_/B vssd1 vssd1 vccd1 vccd1 _15558_/Y sky130_fd_sc_hd__nor2_1
XTAP_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14509_ _14509_/A _14509_/B _14509_/C vssd1 vssd1 vccd1 vccd1 _14512_/A sky130_fd_sc_hd__nor3_1
XFILLER_174_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15489_ _15489_/A _15489_/B vssd1 vssd1 vccd1 vccd1 _15499_/A sky130_fd_sc_hd__xor2_1
X_17228_ _17585_/Q _17273_/A2 _17273_/B1 vssd1 vssd1 vccd1 vccd1 _17228_/X sky130_fd_sc_hd__a21o_1
Xinput30 i_wb_addr[5] vssd1 vssd1 vccd1 vccd1 input30/X sky130_fd_sc_hd__clkbuf_1
Xinput41 i_wb_data[14] vssd1 vssd1 vccd1 vccd1 input41/X sky130_fd_sc_hd__clkbuf_1
Xinput52 i_wb_data[24] vssd1 vssd1 vccd1 vccd1 input52/X sky130_fd_sc_hd__clkbuf_1
XFILLER_116_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput63 i_wb_data[5] vssd1 vssd1 vccd1 vccd1 input63/X sky130_fd_sc_hd__clkbuf_1
XFILLER_128_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17159_ _11778_/Y _17157_/Y _17158_/Y vssd1 vssd1 vccd1 vccd1 _17166_/A sky130_fd_sc_hd__o21ai_1
XFILLER_155_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09981_ _09982_/A _09980_/Y _10111_/C _09981_/D vssd1 vssd1 vccd1 vccd1 _10113_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_131_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08932_ _08872_/X _08874_/X _08930_/A _08929_/Y vssd1 vssd1 vccd1 vccd1 _09016_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_112_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08863_ _08864_/B _08864_/A vssd1 vssd1 vccd1 vccd1 _08863_/X sky130_fd_sc_hd__and2b_1
XFILLER_69_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08794_ _11878_/B _08794_/B vssd1 vssd1 vccd1 vccd1 _08796_/B sky130_fd_sc_hd__nor2_1
XFILLER_26_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09415_ _09415_/A _09415_/B vssd1 vssd1 vccd1 vccd1 _09416_/B sky130_fd_sc_hd__nor2_1
XFILLER_13_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09346_ _09346_/A _09346_/B vssd1 vssd1 vccd1 vccd1 _09370_/A sky130_fd_sc_hd__or2_1
XFILLER_139_826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09277_ _09290_/B _09290_/C _09290_/A vssd1 vssd1 vccd1 vccd1 _09292_/A sky130_fd_sc_hd__a21o_1
XFILLER_166_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11170_ _11021_/X _11041_/A _11168_/Y _11169_/X vssd1 vssd1 vccd1 vccd1 _11202_/A
+ sky130_fd_sc_hd__a211o_1
X_10121_ _10133_/B _10133_/C _10133_/A vssd1 vssd1 vccd1 vccd1 _10134_/A sky130_fd_sc_hd__a21o_1
XFILLER_79_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10052_ _10074_/B _10052_/B vssd1 vssd1 vccd1 vccd1 _10053_/C sky130_fd_sc_hd__and2_1
XFILLER_0_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14860_ _16399_/A _16399_/B vssd1 vssd1 vccd1 vccd1 _16400_/B sky130_fd_sc_hd__and2_1
XFILLER_29_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13811_ _13812_/A _13812_/B vssd1 vssd1 vccd1 vccd1 _13921_/B sky130_fd_sc_hd__or2_1
XFILLER_75_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14791_ _15715_/A _15110_/A vssd1 vssd1 vccd1 vccd1 _14791_/X sky130_fd_sc_hd__or2_1
XFILLER_28_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16530_ _16437_/A _16437_/B _16435_/X vssd1 vssd1 vccd1 vccd1 _16543_/A sky130_fd_sc_hd__a21o_1
XFILLER_44_732 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13742_ _13742_/A _13742_/B vssd1 vssd1 vccd1 vccd1 _13748_/A sky130_fd_sc_hd__nor2_1
XFILLER_113_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10954_ _10954_/A _11006_/B _17468_/D _10954_/D vssd1 vssd1 vccd1 vccd1 _11010_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_16_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16461_ _16462_/A _16462_/B _16460_/Y vssd1 vssd1 vccd1 vccd1 _16557_/A sky130_fd_sc_hd__o21ba_1
XFILLER_73_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13673_ _13670_/Y _13770_/B _13558_/A _13559_/Y vssd1 vssd1 vccd1 vccd1 _13710_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_71_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10885_ _11629_/A _11132_/B _10932_/B _14893_/B vssd1 vssd1 vccd1 vccd1 _10891_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_31_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15412_ _15493_/A _15932_/A vssd1 vssd1 vccd1 vccd1 _15414_/A sky130_fd_sc_hd__nor2_1
X_12624_ _12780_/A _12624_/B vssd1 vssd1 vccd1 vccd1 _12626_/C sky130_fd_sc_hd__nand2_1
X_16392_ _14776_/A _16391_/Y _16390_/Y vssd1 vssd1 vccd1 vccd1 _16396_/A sky130_fd_sc_hd__a21o_1
XFILLER_129_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_611 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15343_ _15342_/A _15661_/A _15340_/X vssd1 vssd1 vccd1 vccd1 _15345_/A sky130_fd_sc_hd__a21oi_1
X_12555_ _12542_/Y _12555_/B vssd1 vssd1 vccd1 vccd1 _17580_/D sky130_fd_sc_hd__nand2b_1
XFILLER_12_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11506_ _11506_/A _11506_/B _11629_/D _11605_/B vssd1 vssd1 vccd1 vccd1 _11506_/X
+ sky130_fd_sc_hd__and4_1
X_15274_ _15274_/A _15493_/A _15402_/B vssd1 vssd1 vccd1 vccd1 _15277_/A sky130_fd_sc_hd__or3b_1
XFILLER_7_143 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12486_ _12787_/B _12637_/D _12487_/D _12487_/A vssd1 vssd1 vccd1 vccd1 _12490_/A
+ sky130_fd_sc_hd__a22oi_1
X_17013_ _17013_/A vssd1 vssd1 vccd1 vccd1 _17014_/C sky130_fd_sc_hd__inv_2
X_14225_ _14225_/A _14225_/B vssd1 vssd1 vccd1 vccd1 _14227_/A sky130_fd_sc_hd__nor2_1
XFILLER_171_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11437_ _11518_/A _11518_/B _14895_/B _11437_/D vssd1 vssd1 vccd1 vccd1 _11440_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_171_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14156_ _14156_/A _14156_/B vssd1 vssd1 vccd1 vccd1 _14158_/C sky130_fd_sc_hd__xnor2_1
X_11368_ _11367_/A _11367_/C _11448_/A vssd1 vssd1 vccd1 vccd1 _11368_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_98_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13107_ _13107_/A _13107_/B vssd1 vssd1 vccd1 vccd1 _13109_/B sky130_fd_sc_hd__nor2_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10319_ _10319_/A _10330_/B _10319_/C _10319_/D vssd1 vssd1 vccd1 vccd1 _10319_/Y
+ sky130_fd_sc_hd__nand4_4
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14087_ _14086_/B _14087_/B vssd1 vssd1 vccd1 vccd1 _14088_/B sky130_fd_sc_hd__nand2b_1
XFILLER_113_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11299_ _11299_/A _11299_/B _11299_/C vssd1 vssd1 vccd1 vccd1 _11415_/A sky130_fd_sc_hd__or3_1
XFILLER_3_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13038_ _13038_/A _13038_/B vssd1 vssd1 vccd1 vccd1 _13040_/C sky130_fd_sc_hd__xnor2_1
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_526 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14989_ _14986_/Y _14988_/Y _15384_/S vssd1 vssd1 vccd1 vccd1 _14989_/X sky130_fd_sc_hd__mux2_1
XFILLER_93_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16728_ _16727_/B _16728_/B vssd1 vssd1 vccd1 vccd1 _16728_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_35_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16659_ _08743_/A _16639_/Y _16658_/X vssd1 vssd1 vccd1 vccd1 _16659_/X sky130_fd_sc_hd__o21a_1
XFILLER_90_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09200_ _09227_/B _09200_/B vssd1 vssd1 vccd1 vccd1 _09211_/A sky130_fd_sc_hd__and2_1
XFILLER_22_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09131_ _09167_/A _09137_/B vssd1 vssd1 vccd1 vccd1 _09131_/X sky130_fd_sc_hd__and2_1
XFILLER_147_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_667 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09062_ _09063_/B _09063_/A vssd1 vssd1 vccd1 vccd1 _09062_/X sky130_fd_sc_hd__and2b_1
XFILLER_163_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_188 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09964_ _09964_/A _10091_/A vssd1 vssd1 vccd1 vccd1 _09966_/B sky130_fd_sc_hd__nor2_1
XFILLER_89_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08915_ _08916_/A _08914_/Y _17381_/A _12088_/D vssd1 vssd1 vccd1 vccd1 _09057_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_58_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09895_ _09895_/A _10021_/A vssd1 vssd1 vccd1 vccd1 _09902_/A sky130_fd_sc_hd__nor2_1
XFILLER_112_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_59 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08846_ _08947_/B _11902_/B _08860_/B _09078_/A vssd1 vssd1 vccd1 vccd1 _08846_/Y
+ sky130_fd_sc_hd__a22oi_1
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_827 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08777_ _08777_/A _08777_/B vssd1 vssd1 vccd1 vccd1 _08779_/A sky130_fd_sc_hd__nor2_1
XFILLER_45_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10670_ _10670_/A _10670_/B vssd1 vssd1 vccd1 vccd1 _10673_/A sky130_fd_sc_hd__nand2_1
XFILLER_167_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09329_ _09332_/B _09329_/B vssd1 vssd1 vccd1 vccd1 _09462_/C sky130_fd_sc_hd__and2_1
XFILLER_139_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12340_ _17415_/A _12340_/B vssd1 vssd1 vccd1 vccd1 _12341_/B sky130_fd_sc_hd__nand2_1
XFILLER_166_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12271_ _12271_/A _12271_/B vssd1 vssd1 vccd1 vccd1 _12273_/A sky130_fd_sc_hd__nor2_1
XFILLER_153_136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14010_ _14115_/B _14010_/B vssd1 vssd1 vccd1 vccd1 _14011_/B sky130_fd_sc_hd__and2_1
XFILLER_153_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11222_ _11222_/A _11222_/B vssd1 vssd1 vccd1 vccd1 _11223_/B sky130_fd_sc_hd__or2_1
XFILLER_135_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1014 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11153_ _11153_/A _11153_/B _11153_/C vssd1 vssd1 vccd1 vccd1 _11154_/C sky130_fd_sc_hd__nor3_1
XFILLER_96_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10104_ _10027_/B _10027_/C _10025_/Y _10028_/A vssd1 vssd1 vccd1 vccd1 _10104_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_150_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11084_ _11084_/A _11084_/B _11084_/C vssd1 vssd1 vccd1 vccd1 _11090_/A sky130_fd_sc_hd__nor3_1
X_15961_ _15855_/A _15855_/B _15852_/Y vssd1 vssd1 vccd1 vccd1 _15963_/B sky130_fd_sc_hd__o21a_1
XFILLER_150_898 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14912_ _12442_/A _14912_/B vssd1 vssd1 vccd1 vccd1 _14912_/Y sky130_fd_sc_hd__nand2b_1
X_10035_ _10035_/A _10035_/B vssd1 vssd1 vccd1 vccd1 _10050_/A sky130_fd_sc_hd__nand2_1
XFILLER_103_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15892_ _15797_/Y _15798_/Y _15797_/A vssd1 vssd1 vccd1 vccd1 _15892_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_48_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14843_ _14929_/A _14938_/B vssd1 vssd1 vccd1 vccd1 _15248_/C sky130_fd_sc_hd__nor2_2
XFILLER_84_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17562_ fanout952/X _17562_/D vssd1 vssd1 vccd1 vccd1 _17562_/Q sky130_fd_sc_hd__dfxtp_1
X_14774_ _14774_/A _16571_/A vssd1 vssd1 vccd1 vccd1 _16576_/B sky130_fd_sc_hd__or2_1
XFILLER_95_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11986_ _11985_/B _11986_/B vssd1 vssd1 vccd1 vccd1 _11987_/B sky130_fd_sc_hd__and2b_1
XFILLER_16_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16513_ _16514_/A _16938_/B _16514_/C vssd1 vssd1 vccd1 vccd1 _16515_/A sky130_fd_sc_hd__o21ai_1
XFILLER_16_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13725_ _13726_/A _13726_/B vssd1 vssd1 vccd1 vccd1 _13727_/A sky130_fd_sc_hd__nor2_1
X_10937_ _10938_/A _10938_/B vssd1 vssd1 vccd1 vccd1 _10990_/A sky130_fd_sc_hd__nand2_1
X_17493_ fanout943/X _17493_/D vssd1 vssd1 vccd1 vccd1 _17493_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_44_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16444_ _16444_/A _16444_/B vssd1 vssd1 vccd1 vccd1 _16455_/A sky130_fd_sc_hd__or2_1
XFILLER_149_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13656_ _13654_/X _13656_/B vssd1 vssd1 vccd1 vccd1 _13659_/A sky130_fd_sc_hd__nand2b_1
XFILLER_31_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10868_ _11117_/C _10963_/C vssd1 vssd1 vccd1 vccd1 _11100_/A sky130_fd_sc_hd__nand2_2
XFILLER_31_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12607_ _12607_/A _12607_/B _12607_/C vssd1 vssd1 vccd1 vccd1 _12608_/B sky130_fd_sc_hd__or3_1
X_16375_ _16375_/A _16375_/B vssd1 vssd1 vccd1 vccd1 _16378_/A sky130_fd_sc_hd__xnor2_2
XPHY_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13587_ _13587_/A _13587_/B vssd1 vssd1 vccd1 vccd1 _13589_/A sky130_fd_sc_hd__nor2_1
XPHY_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10799_ _14787_/A _10799_/B vssd1 vssd1 vccd1 vccd1 _10799_/Y sky130_fd_sc_hd__nand2_1
XFILLER_9_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15326_ _14882_/X _15325_/X _17377_/A vssd1 vssd1 vccd1 vccd1 _16695_/A sky130_fd_sc_hd__a21oi_4
XFILLER_12_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_818 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12538_ _12540_/A _12540_/B vssd1 vssd1 vccd1 vccd1 _12538_/Y sky130_fd_sc_hd__nand2_1
XFILLER_117_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15257_ _15257_/A _15257_/B _15257_/C _15256_/X vssd1 vssd1 vccd1 vccd1 _15257_/X
+ sky130_fd_sc_hd__or4b_1
XFILLER_172_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12469_ _12271_/A _12273_/B _12271_/B vssd1 vssd1 vccd1 vccd1 _12473_/A sky130_fd_sc_hd__o21ba_1
X_14208_ _14763_/S _14206_/Y _14207_/X _14129_/Y vssd1 vssd1 vccd1 vccd1 _17594_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_132_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15188_ _15188_/A _15188_/B vssd1 vssd1 vccd1 vccd1 _15188_/Y sky130_fd_sc_hd__nor2_1
XFILLER_113_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14139_ _14221_/A _14139_/B vssd1 vssd1 vccd1 vccd1 _14148_/A sky130_fd_sc_hd__or2_1
Xfanout409 _12068_/A vssd1 vssd1 vccd1 vccd1 _17403_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_3_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09680_ _09678_/B _09675_/C _09675_/B vssd1 vssd1 vccd1 vccd1 _09681_/B sky130_fd_sc_hd__o21a_1
XFILLER_67_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_624 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09114_ _09115_/A _09115_/B _09115_/C vssd1 vssd1 vccd1 vccd1 _09114_/Y sky130_fd_sc_hd__nor3_1
XFILLER_136_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09045_ _17387_/A _09042_/B _09044_/B _09041_/Y vssd1 vssd1 vccd1 vccd1 _09047_/B
+ sky130_fd_sc_hd__a31oi_1
XFILLER_163_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout910 _10905_/D vssd1 vssd1 vccd1 vccd1 _11095_/D sky130_fd_sc_hd__buf_2
Xfanout921 _17284_/C1 vssd1 vssd1 vccd1 vccd1 _17293_/C1 sky130_fd_sc_hd__buf_2
XFILLER_131_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout932 _17428_/B vssd1 vssd1 vccd1 vccd1 _17378_/C1 sky130_fd_sc_hd__clkbuf_4
XFILLER_89_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09947_ _10321_/B _10203_/B vssd1 vssd1 vccd1 vccd1 _10061_/A sky130_fd_sc_hd__nand2_1
XFILLER_104_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout943 fanout944/X vssd1 vssd1 vccd1 vccd1 fanout943/X sky130_fd_sc_hd__clkbuf_2
Xfanout954 fanout957/X vssd1 vssd1 vccd1 vccd1 fanout954/X sky130_fd_sc_hd__clkbuf_4
XFILLER_58_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09878_ _09878_/A _09878_/B vssd1 vssd1 vccd1 vccd1 _10007_/A sky130_fd_sc_hd__xnor2_1
XFILLER_100_740 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08829_ _08828_/B _08829_/B vssd1 vssd1 vccd1 vccd1 _08869_/B sky130_fd_sc_hd__nand2b_1
XFILLER_45_304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11840_ _12046_/A _11840_/B vssd1 vssd1 vccd1 vccd1 _11840_/Y sky130_fd_sc_hd__nand2_1
XTAP_2635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11771_ _11771_/A _11771_/B vssd1 vssd1 vccd1 vccd1 _11771_/Y sky130_fd_sc_hd__nand2_1
XFILLER_54_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13510_ _13267_/X _13511_/B _13509_/Y _13385_/B vssd1 vssd1 vccd1 vccd1 _13510_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10722_ _10722_/A _10722_/B vssd1 vssd1 vccd1 vccd1 _11174_/A sky130_fd_sc_hd__xnor2_1
XFILLER_14_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14490_ _14557_/B _14490_/B vssd1 vssd1 vccd1 vccd1 _14519_/A sky130_fd_sc_hd__nor2_1
XFILLER_13_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13441_ _13441_/A vssd1 vssd1 vccd1 vccd1 _13600_/A sky130_fd_sc_hd__inv_2
X_10653_ _10653_/A _10653_/B _10653_/C vssd1 vssd1 vccd1 vccd1 _10662_/B sky130_fd_sc_hd__nand3_1
XFILLER_110_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16160_ _16161_/A _16161_/B vssd1 vssd1 vccd1 vccd1 _16160_/X sky130_fd_sc_hd__or2_1
XFILLER_139_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13372_ _13496_/A _13370_/Y _13240_/Y _13244_/B vssd1 vssd1 vccd1 vccd1 _13373_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_154_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10584_ _10579_/A _10577_/X _10325_/A _10329_/B vssd1 vssd1 vccd1 vccd1 _10584_/X
+ sky130_fd_sc_hd__o211a_1
X_15111_ _11469_/X _15804_/A2 _15713_/B1 _15110_/A vssd1 vssd1 vccd1 vccd1 _15111_/X
+ sky130_fd_sc_hd__a22o_1
X_12323_ _12323_/A _12492_/A _12323_/C vssd1 vssd1 vccd1 vccd1 _12492_/B sky130_fd_sc_hd__nor3_1
X_16091_ _16092_/A _16092_/B vssd1 vssd1 vccd1 vccd1 _16200_/A sky130_fd_sc_hd__nand2b_1
XFILLER_154_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15042_ _15130_/S _15042_/B _15450_/B vssd1 vssd1 vccd1 vccd1 _15042_/X sky130_fd_sc_hd__or3_1
XFILLER_114_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12254_ _12078_/A _12080_/B _12078_/B vssd1 vssd1 vccd1 vccd1 _12261_/A sky130_fd_sc_hd__o21ba_1
XFILLER_141_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_692 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11205_ _11739_/A _11205_/B vssd1 vssd1 vccd1 vccd1 _11221_/A sky130_fd_sc_hd__nand2_1
XFILLER_79_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12185_ _11988_/A _11988_/B _11987_/A vssd1 vssd1 vccd1 vccd1 _12186_/B sky130_fd_sc_hd__a21oi_1
XFILLER_123_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11136_ _11137_/B _11137_/C _11137_/A vssd1 vssd1 vccd1 vccd1 _11293_/A sky130_fd_sc_hd__o21ai_1
X_16993_ _17046_/B _16993_/B vssd1 vssd1 vccd1 vccd1 _16996_/B sky130_fd_sc_hd__and2b_1
XFILLER_62_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11067_ _11069_/B vssd1 vssd1 vccd1 vccd1 _11067_/Y sky130_fd_sc_hd__inv_2
X_15944_ _15944_/A _15944_/B vssd1 vssd1 vccd1 vccd1 _15972_/A sky130_fd_sc_hd__xnor2_1
XFILLER_110_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_62 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10018_ _10018_/A _10018_/B _10019_/B vssd1 vssd1 vccd1 vccd1 _10023_/B sky130_fd_sc_hd__or3_1
XFILLER_92_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15875_ _15875_/A _15875_/B vssd1 vssd1 vccd1 vccd1 _15875_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17614_ fanout954/X _17614_/D vssd1 vssd1 vccd1 vccd1 _17614_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_64_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14826_ _17023_/A _14825_/Y _14764_/Y _14434_/Y vssd1 vssd1 vccd1 vccd1 _14826_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_45_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14757_ _13832_/B _13834_/A _14757_/S vssd1 vssd1 vccd1 vccd1 _14758_/B sky130_fd_sc_hd__mux2_1
X_17545_ fanout954/X _17545_/D vssd1 vssd1 vccd1 vccd1 _17545_/Q sky130_fd_sc_hd__dfxtp_4
X_11969_ _11970_/A _11970_/B vssd1 vssd1 vccd1 vccd1 _11971_/A sky130_fd_sc_hd__or2_1
X_13708_ _13594_/X _13598_/A _13706_/Y _13707_/X vssd1 vssd1 vccd1 vccd1 _13817_/A
+ sky130_fd_sc_hd__o211a_1
X_17476_ fanout956/X _17476_/D vssd1 vssd1 vccd1 vccd1 _17476_/Q sky130_fd_sc_hd__dfxtp_1
X_14688_ _14688_/A _14688_/B vssd1 vssd1 vccd1 vccd1 _14689_/B sky130_fd_sc_hd__nand2_1
X_16427_ _16333_/X _16337_/B _16335_/B vssd1 vssd1 vccd1 vccd1 _16437_/A sky130_fd_sc_hd__o21ai_1
X_13639_ _13638_/A _13638_/B _13638_/C vssd1 vssd1 vccd1 vccd1 _13645_/B sky130_fd_sc_hd__a21o_1
XFILLER_32_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16358_ _16358_/A _16358_/B _16358_/C vssd1 vssd1 vccd1 vccd1 _16359_/B sky130_fd_sc_hd__or3_1
XFILLER_158_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_615 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15309_ _15309_/A _16111_/A _15307_/X vssd1 vssd1 vccd1 vccd1 _15321_/A sky130_fd_sc_hd__or3b_1
XFILLER_172_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16289_ _16290_/A _16290_/B _16290_/C vssd1 vssd1 vccd1 vccd1 _16382_/B sky130_fd_sc_hd__o21a_1
XFILLER_145_467 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_82 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout206 _14912_/B vssd1 vssd1 vccd1 vccd1 _14911_/B sky130_fd_sc_hd__buf_2
Xfanout217 _15638_/Y vssd1 vssd1 vccd1 vccd1 _16591_/B sky130_fd_sc_hd__buf_2
X_09801_ _09801_/A _09801_/B _09941_/A vssd1 vssd1 vccd1 vccd1 _09802_/B sky130_fd_sc_hd__nor3_1
XFILLER_87_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout228 _14933_/Y vssd1 vssd1 vccd1 vccd1 _16008_/B1 sky130_fd_sc_hd__clkbuf_2
XFILLER_101_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout239 _16401_/C1 vssd1 vssd1 vccd1 vccd1 _17162_/C1 sky130_fd_sc_hd__clkbuf_4
XFILLER_101_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09732_ _09733_/B _09733_/A vssd1 vssd1 vccd1 vccd1 _09732_/X sky130_fd_sc_hd__and2b_1
XFILLER_55_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09663_ _09499_/Y _09500_/X _09789_/A _09774_/B _09774_/A vssd1 vssd1 vccd1 vccd1
+ _09665_/B sky130_fd_sc_hd__a32o_1
XFILLER_82_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09594_ _09588_/X _09723_/A _09580_/X _09581_/Y vssd1 vssd1 vccd1 vccd1 _09597_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_82_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_721 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_795 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09028_ _13028_/A _12787_/D vssd1 vssd1 vccd1 vccd1 _17081_/A sky130_fd_sc_hd__nand2_8
XFILLER_164_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout740 _10171_/D vssd1 vssd1 vccd1 vccd1 _11841_/B sky130_fd_sc_hd__buf_4
XFILLER_104_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout751 _12334_/B vssd1 vssd1 vccd1 vccd1 _12942_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_131_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout762 fanout772/X vssd1 vssd1 vccd1 vccd1 _12787_/D sky130_fd_sc_hd__buf_2
Xfanout773 _17491_/Q vssd1 vssd1 vccd1 vccd1 _13434_/D sky130_fd_sc_hd__buf_2
X_13990_ _13990_/A _13990_/B vssd1 vssd1 vccd1 vccd1 _14011_/A sky130_fd_sc_hd__xor2_1
Xfanout784 fanout795/X vssd1 vssd1 vccd1 vccd1 _13321_/D sky130_fd_sc_hd__buf_2
Xfanout795 _17490_/Q vssd1 vssd1 vccd1 vccd1 fanout795/X sky130_fd_sc_hd__buf_6
XTAP_3100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12941_ _13450_/B _13080_/D _12942_/D _13080_/A vssd1 vssd1 vccd1 vccd1 _12945_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_46_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15660_ _16056_/A _15661_/A _16259_/B vssd1 vssd1 vccd1 vccd1 _15660_/X sky130_fd_sc_hd__and3_1
XTAP_3155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12872_ _12872_/A _12872_/B vssd1 vssd1 vccd1 vccd1 _12875_/A sky130_fd_sc_hd__xnor2_1
XANTENNA_100 _09412_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14611_ _14612_/A _14612_/B vssd1 vssd1 vccd1 vccd1 _14693_/A sky130_fd_sc_hd__and2b_1
XTAP_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11823_ _17304_/A1 _17302_/A1 _12050_/S vssd1 vssd1 vccd1 vccd1 _11824_/B sky130_fd_sc_hd__mux2_1
XTAP_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15591_ _15591_/A _15591_/B vssd1 vssd1 vccd1 vccd1 _15601_/A sky130_fd_sc_hd__or2_1
XFILLER_14_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17330_ _10297_/D _17360_/A2 _17329_/X _17408_/C1 vssd1 vssd1 vccd1 vccd1 _17494_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14542_ _12710_/A _13015_/B _14210_/B _13012_/X vssd1 vssd1 vccd1 vccd1 _14543_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11754_ _11753_/A _11753_/B _11753_/C vssd1 vssd1 vccd1 vccd1 _11755_/B sky130_fd_sc_hd__a21o_1
XFILLER_60_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10705_ _10705_/A _10705_/B vssd1 vssd1 vccd1 vccd1 _11030_/B sky130_fd_sc_hd__nor2_1
XFILLER_42_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17261_ _17596_/Q _17282_/A2 _17282_/B1 vssd1 vssd1 vccd1 vccd1 _17261_/X sky130_fd_sc_hd__a21o_1
XTAP_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14473_ _14473_/A _14473_/B _14473_/C vssd1 vssd1 vccd1 vccd1 _14533_/B sky130_fd_sc_hd__nand3_1
X_11685_ _15235_/A _15235_/B vssd1 vssd1 vccd1 vccd1 _11688_/A sky130_fd_sc_hd__nor2_1
XFILLER_128_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16212_ _16107_/Y _16111_/B _16210_/Y vssd1 vssd1 vccd1 vccd1 _16212_/Y sky130_fd_sc_hd__o21ai_1
X_13424_ _13308_/A _13309_/B _13421_/Y _13422_/X vssd1 vssd1 vccd1 vccd1 _13428_/A
+ sky130_fd_sc_hd__a211oi_2
XFILLER_174_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10636_ _10550_/X _10634_/Y _10632_/B _10614_/X vssd1 vssd1 vccd1 vccd1 _10636_/Y
+ sky130_fd_sc_hd__o211ai_1
X_17192_ input18/X input17/X input19/X input23/X vssd1 vssd1 vccd1 vccd1 _17195_/A
+ sky130_fd_sc_hd__or4b_1
XFILLER_167_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16143_ _16241_/B _16143_/B vssd1 vssd1 vccd1 vccd1 _16146_/A sky130_fd_sc_hd__nor2_1
X_13355_ _13355_/A _13355_/B vssd1 vssd1 vccd1 vccd1 _13357_/B sky130_fd_sc_hd__xnor2_1
XFILLER_127_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10567_ _10567_/A _10567_/B vssd1 vssd1 vccd1 vccd1 _10569_/B sky130_fd_sc_hd__or2_1
XFILLER_155_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12306_ _12306_/A _12306_/B vssd1 vssd1 vccd1 vccd1 _12307_/B sky130_fd_sc_hd__nor2_1
X_16074_ _16075_/A _16075_/B vssd1 vssd1 vccd1 vccd1 _16188_/B sky130_fd_sc_hd__and2b_1
X_13286_ _13745_/B _13735_/D _13632_/D _13852_/A vssd1 vssd1 vccd1 vccd1 _13286_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_5_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10498_ _10589_/A _10589_/B vssd1 vssd1 vccd1 vccd1 _10499_/A sky130_fd_sc_hd__or2_2
XFILLER_142_437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15025_ _15305_/C _15025_/B vssd1 vssd1 vccd1 vccd1 _15025_/Y sky130_fd_sc_hd__nor2_1
X_12237_ _12871_/A _13208_/D vssd1 vssd1 vccd1 vccd1 _12238_/B sky130_fd_sc_hd__nand2_1
XFILLER_69_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_90 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12168_ _12169_/A _12169_/B _12169_/C vssd1 vssd1 vccd1 vccd1 _12170_/A sky130_fd_sc_hd__a21oi_1
XFILLER_111_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11119_ _11124_/C _10971_/B _10878_/A _10876_/Y vssd1 vssd1 vccd1 vccd1 _11121_/C
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_1_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12099_ _11891_/A _11891_/Y _12097_/X _12268_/B vssd1 vssd1 vccd1 vccd1 _12122_/A
+ sky130_fd_sc_hd__o211ai_4
X_16976_ _16735_/A _14590_/B _17164_/C _15628_/B vssd1 vssd1 vccd1 vccd1 _16977_/C
+ sky130_fd_sc_hd__o22a_1
X_15927_ _15925_/Y _15927_/B vssd1 vssd1 vccd1 vccd1 _15941_/A sky130_fd_sc_hd__and2b_1
Xinput6 i_wb_addr[12] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__clkbuf_1
XFILLER_49_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15858_ _15858_/A _15858_/B vssd1 vssd1 vccd1 vccd1 _15859_/B sky130_fd_sc_hd__xnor2_1
XFILLER_18_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_774 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14809_ _15707_/B _15707_/C _10145_/B vssd1 vssd1 vccd1 vccd1 _15802_/A sky130_fd_sc_hd__a21o_1
XFILLER_17_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15789_ _15610_/A _15698_/A _15698_/B vssd1 vssd1 vccd1 vccd1 _15789_/X sky130_fd_sc_hd__o21ba_1
XFILLER_33_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17528_ fanout945/X _17528_/D vssd1 vssd1 vccd1 vccd1 _17528_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_60_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17459_ fanout933/X _17459_/D vssd1 vssd1 vccd1 vccd1 _17459_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_118_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_580 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_49 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_194 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09715_ _09711_/X _09713_/X _16982_/B _09710_/Y vssd1 vssd1 vccd1 vccd1 _09717_/B
+ sky130_fd_sc_hd__o2bb2a_2
XFILLER_28_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_410 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09646_ _09969_/A _09646_/B vssd1 vssd1 vccd1 vccd1 _09647_/C sky130_fd_sc_hd__nor2_1
XFILLER_71_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_115 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09577_ _09577_/A _09577_/B _09596_/B vssd1 vssd1 vccd1 vccd1 _09624_/B sky130_fd_sc_hd__and3_1
XFILLER_35_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_958 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_824 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_34 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11470_ _11470_/A _11561_/D vssd1 vssd1 vccd1 vccd1 _11472_/B sky130_fd_sc_hd__nand2_1
XFILLER_137_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10421_ _10422_/A _10420_/Y _15805_/A _10421_/D vssd1 vssd1 vccd1 vccd1 _10531_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_13_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_916 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13140_ _13268_/B _13140_/B vssd1 vssd1 vccd1 vccd1 _13140_/Y sky130_fd_sc_hd__nand2_1
X_10352_ _10352_/A _10352_/B vssd1 vssd1 vccd1 vccd1 _10465_/A sky130_fd_sc_hd__xor2_1
XFILLER_164_595 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_908 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13071_ _13072_/A _13072_/B _13072_/C vssd1 vssd1 vccd1 vccd1 _13244_/A sky130_fd_sc_hd__o21a_1
X_10283_ _10283_/A _10283_/B _10283_/C _10283_/D vssd1 vssd1 vccd1 vccd1 _10283_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_105_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12022_ _10180_/C _14952_/B wire209/X vssd1 vssd1 vccd1 vccd1 _12022_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_105_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16830_ _16830_/A _16830_/B vssd1 vssd1 vccd1 vccd1 _16832_/B sky130_fd_sc_hd__xnor2_1
XFILLER_93_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout570 _17513_/Q vssd1 vssd1 vccd1 vccd1 _15538_/A sky130_fd_sc_hd__buf_2
Xfanout581 _16011_/B vssd1 vssd1 vccd1 vccd1 _15254_/S sky130_fd_sc_hd__buf_2
Xfanout592 _14982_/A vssd1 vssd1 vccd1 vccd1 _12700_/B sky130_fd_sc_hd__clkbuf_4
X_16761_ _16761_/A _16761_/B vssd1 vssd1 vccd1 vccd1 _16762_/B sky130_fd_sc_hd__xnor2_1
XFILLER_19_624 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13973_ _13864_/B _13870_/B _13862_/X vssd1 vssd1 vccd1 vccd1 _13974_/B sky130_fd_sc_hd__a21oi_1
XFILLER_46_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12924_ _12924_/A _12924_/B vssd1 vssd1 vccd1 vccd1 _12926_/A sky130_fd_sc_hd__nor2_1
X_15712_ _15715_/A _15103_/X _15711_/Y _16582_/A vssd1 vssd1 vccd1 vccd1 _15712_/X
+ sky130_fd_sc_hd__a211o_1
X_16692_ _16693_/B _16692_/B vssd1 vssd1 vccd1 vccd1 _16777_/A sky130_fd_sc_hd__nand2b_1
XFILLER_74_763 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_605 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15643_ _15732_/A _15643_/B vssd1 vssd1 vccd1 vccd1 _15742_/A sky130_fd_sc_hd__nand2_1
X_12855_ _14421_/S _12852_/X _14482_/B1 _12850_/X vssd1 vssd1 vccd1 vccd1 _12856_/B
+ sky130_fd_sc_hd__o31a_1
XTAP_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11806_ _12025_/A _14863_/A _09926_/C vssd1 vssd1 vccd1 vccd1 _11807_/B sky130_fd_sc_hd__a21o_1
X_15574_ _16760_/A _08731_/A _16315_/D vssd1 vssd1 vccd1 vccd1 _15658_/B sky130_fd_sc_hd__a21oi_1
XFILLER_33_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12786_ _12787_/B _12942_/D _12787_/D _13080_/A vssd1 vssd1 vccd1 vccd1 _12790_/A
+ sky130_fd_sc_hd__a22oi_1
XTAP_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17313_ input66/X _17321_/B _17321_/C vssd1 vssd1 vccd1 vccd1 _17313_/X sky130_fd_sc_hd__or3_1
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14525_ _14524_/A _14524_/B _14524_/C vssd1 vssd1 vccd1 vccd1 _14526_/B sky130_fd_sc_hd__o21ai_1
X_11737_ _11739_/B vssd1 vssd1 vccd1 vccd1 _11737_/Y sky130_fd_sc_hd__inv_2
XTAP_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14456_ _14456_/A _14456_/B _14456_/C vssd1 vssd1 vccd1 vccd1 _14528_/A sky130_fd_sc_hd__nand3_1
X_17244_ _17558_/Q _17244_/B vssd1 vssd1 vccd1 vccd1 _17244_/X sky130_fd_sc_hd__and2_1
X_11668_ _11646_/A _11646_/B _11646_/C vssd1 vssd1 vccd1 vccd1 _11670_/C sky130_fd_sc_hd__a21o_1
XFILLER_174_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13407_ _13643_/A _13846_/B vssd1 vssd1 vccd1 vccd1 _13408_/B sky130_fd_sc_hd__nand2_1
X_10619_ _10719_/C _10736_/D vssd1 vssd1 vccd1 vccd1 _10716_/A sky130_fd_sc_hd__nand2_4
X_17175_ input15/X input18/X input17/X input20/X vssd1 vssd1 vccd1 vccd1 _17181_/C
+ sky130_fd_sc_hd__or4_1
X_14387_ _14387_/A _14450_/B vssd1 vssd1 vccd1 vccd1 _14388_/B sky130_fd_sc_hd__nand2_1
X_11599_ _11555_/A _11555_/B _11637_/A vssd1 vssd1 vccd1 vccd1 _11600_/B sky130_fd_sc_hd__o21bai_1
X_16126_ _16315_/B _16681_/D _16938_/D _16025_/A vssd1 vssd1 vccd1 vccd1 _16126_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_115_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13338_ _13338_/A _13455_/B vssd1 vssd1 vccd1 vccd1 _13339_/C sky130_fd_sc_hd__nor2_1
XFILLER_116_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16057_ _16055_/A _15658_/Y _16827_/D _15081_/A vssd1 vssd1 vccd1 vccd1 _16058_/B
+ sky130_fd_sc_hd__o22a_1
X_13269_ _13010_/B _13511_/A _13267_/X vssd1 vssd1 vccd1 vccd1 _13271_/B sky130_fd_sc_hd__a21oi_1
XFILLER_143_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15008_ _15008_/A _15008_/B vssd1 vssd1 vccd1 vccd1 _15008_/X sky130_fd_sc_hd__or2_1
XFILLER_170_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16959_ _17008_/A _17012_/A vssd1 vssd1 vccd1 vccd1 _16960_/B sky130_fd_sc_hd__nand2_1
XFILLER_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09500_ _09620_/A _09500_/B vssd1 vssd1 vccd1 vccd1 _09500_/X sky130_fd_sc_hd__or2_1
XFILLER_110_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_988 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09431_ _10255_/A _10899_/D _09430_/B _09427_/Y vssd1 vssd1 vccd1 vccd1 _09433_/B
+ sky130_fd_sc_hd__a31oi_4
XFILLER_37_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09362_ _09497_/A _09361_/Y _09502_/A _09362_/D vssd1 vssd1 vccd1 vccd1 _09504_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_80_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_1046 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09293_ _09293_/A _09293_/B vssd1 vssd1 vccd1 vccd1 _09294_/B sky130_fd_sc_hd__nor2_1
XFILLER_123_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_11 _12869_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_22 _17529_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_33 _17546_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_44 _17389_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_55 fanout699/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_66 _09843_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_77 _14939_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_88 fanout699/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_99 _16935_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10970_ _10970_/A _10970_/B vssd1 vssd1 vccd1 vccd1 _10974_/A sky130_fd_sc_hd__nand2_1
XFILLER_44_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09629_ _09629_/A _09629_/B vssd1 vssd1 vccd1 vccd1 _09632_/A sky130_fd_sc_hd__nand2_1
XFILLER_83_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12640_ _12640_/A _12792_/A _12640_/C vssd1 vssd1 vccd1 vccd1 _12792_/B sky130_fd_sc_hd__nor3_1
XFILLER_62_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12571_ _12572_/A _12572_/B _12572_/C vssd1 vssd1 vccd1 vccd1 _12585_/A sky130_fd_sc_hd__o21ai_1
X_14310_ _14230_/B _14232_/B _14230_/A vssd1 vssd1 vccd1 vccd1 _14312_/B sky130_fd_sc_hd__o21ba_1
X_11522_ _11522_/A _11522_/B _11523_/B vssd1 vssd1 vccd1 vccd1 _11576_/A sky130_fd_sc_hd__or3_1
XFILLER_129_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15290_ _16086_/A _16317_/B _15291_/A vssd1 vssd1 vccd1 vccd1 _15363_/A sky130_fd_sc_hd__and3_1
XFILLER_156_326 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14241_ _14318_/A _14318_/B _14433_/B _14366_/B vssd1 vssd1 vccd1 vccd1 _14242_/B
+ sky130_fd_sc_hd__and4_1
X_11453_ _11453_/A _11453_/B vssd1 vssd1 vccd1 vccd1 _11454_/B sky130_fd_sc_hd__nand2_1
XFILLER_137_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10404_ _10262_/X _10357_/Y _10385_/A _10385_/Y vssd1 vssd1 vccd1 vccd1 _10405_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_139_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14172_ _14173_/A _14173_/B _14173_/C vssd1 vssd1 vccd1 vccd1 _14252_/A sky130_fd_sc_hd__o21ai_1
X_11384_ _11395_/B _11435_/A _11395_/A vssd1 vssd1 vccd1 vccd1 _11384_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_164_381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13123_ _13123_/A _13123_/B vssd1 vssd1 vccd1 vccd1 _13125_/C sky130_fd_sc_hd__or2_1
X_10335_ _10193_/B _10229_/X _10319_/A _10319_/Y vssd1 vssd1 vccd1 vccd1 _10336_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_113_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13054_ _13055_/A _13055_/B vssd1 vssd1 vccd1 vccd1 _13186_/A sky130_fd_sc_hd__or2_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10266_ _10267_/A _10267_/B _10267_/C vssd1 vssd1 vccd1 vccd1 _10266_/X sky130_fd_sc_hd__a21o_2
XFILLER_3_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12005_ _12005_/A _12005_/B vssd1 vssd1 vccd1 vccd1 _12007_/B sky130_fd_sc_hd__nand2_1
XFILLER_78_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10197_ _10198_/A _10198_/C vssd1 vssd1 vccd1 vccd1 _10322_/B sky130_fd_sc_hd__nor2_1
X_16813_ _16883_/A _16813_/B vssd1 vssd1 vccd1 vccd1 _16813_/Y sky130_fd_sc_hd__nor2_1
XFILLER_78_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16744_ _16744_/A _16744_/B vssd1 vssd1 vccd1 vccd1 _16746_/A sky130_fd_sc_hd__nor2_1
X_13956_ _13958_/A _13958_/B vssd1 vssd1 vccd1 vccd1 _14130_/A sky130_fd_sc_hd__nor2_1
XFILLER_47_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12907_ _12907_/A _13948_/C vssd1 vssd1 vccd1 vccd1 _12908_/B sky130_fd_sc_hd__nand2_1
XFILLER_62_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16675_ _16503_/Y _16670_/B _16597_/B _16597_/A vssd1 vssd1 vccd1 vccd1 _16676_/B
+ sky130_fd_sc_hd__a2bb2o_1
X_13887_ _13888_/A _13888_/B vssd1 vssd1 vccd1 vccd1 _13990_/A sky130_fd_sc_hd__nor2_1
XFILLER_46_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12838_ _13001_/B _12837_/Y _12689_/A _12691_/A vssd1 vssd1 vccd1 vccd1 _12838_/Y
+ sky130_fd_sc_hd__a211oi_1
XTAP_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15626_ _15622_/B _16008_/A2 _15625_/X _14944_/A vssd1 vssd1 vccd1 vccd1 _15626_/Y
+ sky130_fd_sc_hd__a211oi_1
XTAP_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15557_ _15557_/A _15557_/B vssd1 vssd1 vccd1 vccd1 _15559_/B sky130_fd_sc_hd__xnor2_1
X_12769_ _12770_/B _12923_/D _12770_/D _12770_/A vssd1 vssd1 vccd1 vccd1 _12771_/A
+ sky130_fd_sc_hd__a22oi_1
XTAP_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14508_ _14508_/A _14508_/B vssd1 vssd1 vccd1 vccd1 _14514_/A sky130_fd_sc_hd__xnor2_1
XFILLER_174_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15488_ _15489_/A _15489_/B vssd1 vssd1 vccd1 vccd1 _15488_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_159_186 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput20 i_wb_addr[25] vssd1 vssd1 vccd1 vccd1 input20/X sky130_fd_sc_hd__clkbuf_1
X_17227_ _17443_/Q _17275_/A2 _17225_/X _17226_/X _17275_/C1 vssd1 vssd1 vccd1 vccd1
+ _17443_/D sky130_fd_sc_hd__o221a_1
Xinput31 i_wb_addr[6] vssd1 vssd1 vccd1 vccd1 input31/X sky130_fd_sc_hd__clkbuf_1
X_14439_ _14440_/A _14440_/B _14440_/C vssd1 vssd1 vccd1 vccd1 _14441_/A sky130_fd_sc_hd__o21a_1
Xinput42 i_wb_data[15] vssd1 vssd1 vccd1 vccd1 input42/X sky130_fd_sc_hd__clkbuf_1
Xinput53 i_wb_data[25] vssd1 vssd1 vccd1 vccd1 input53/X sky130_fd_sc_hd__clkbuf_1
XFILLER_116_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput64 i_wb_data[6] vssd1 vssd1 vccd1 vccd1 input64/X sky130_fd_sc_hd__clkbuf_1
X_17158_ _11778_/Y _17157_/Y _17070_/B vssd1 vssd1 vccd1 vccd1 _17158_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_171_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16109_ _16001_/A _16003_/X _16107_/Y _16108_/X vssd1 vssd1 vccd1 vccd1 _16111_/B
+ sky130_fd_sc_hd__a211oi_2
X_17089_ _17089_/A _17089_/B vssd1 vssd1 vccd1 vccd1 _17118_/A sky130_fd_sc_hd__nor2_1
X_09980_ _10109_/B _09979_/C _10111_/D _09979_/A vssd1 vssd1 vccd1 vccd1 _09980_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_131_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08931_ _08930_/A _08929_/Y _08872_/X _08874_/X vssd1 vssd1 vccd1 vccd1 _09016_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_130_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08862_ _08862_/A _08862_/B vssd1 vssd1 vccd1 vccd1 _08864_/B sky130_fd_sc_hd__nor2_1
XFILLER_57_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08793_ _17387_/A _09319_/C _08790_/Y _11878_/A vssd1 vssd1 vccd1 vccd1 _08794_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_96_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09414_ _09414_/A _17395_/A _09557_/B _12340_/B vssd1 vssd1 vccd1 vccd1 _09415_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_53_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09345_ _09358_/A _09345_/B vssd1 vssd1 vccd1 vccd1 _09346_/B sky130_fd_sc_hd__nor2_1
XFILLER_139_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09276_ _09404_/A _09404_/B vssd1 vssd1 vccd1 vccd1 _09290_/C sky130_fd_sc_hd__nand2_1
XFILLER_138_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_36 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10120_ _10232_/A _10232_/B vssd1 vssd1 vccd1 vccd1 _10133_/C sky130_fd_sc_hd__nand2_1
XFILLER_161_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10051_ _09930_/A _09930_/B _09930_/C vssd1 vssd1 vccd1 vccd1 _10052_/B sky130_fd_sc_hd__o21ai_1
XFILLER_75_302 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13810_ _13923_/A _13810_/B vssd1 vssd1 vccd1 vccd1 _13812_/B sky130_fd_sc_hd__or2_1
XFILLER_75_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14790_ _14889_/C _15175_/B vssd1 vssd1 vccd1 vccd1 _14790_/Y sky130_fd_sc_hd__nor2_1
XFILLER_29_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13741_ _13741_/A _13741_/B _13741_/C vssd1 vssd1 vccd1 vccd1 _13742_/B sky130_fd_sc_hd__nor3_1
X_10953_ _10953_/A _10953_/B vssd1 vssd1 vccd1 vccd1 _11069_/A sky130_fd_sc_hd__xnor2_1
XFILLER_73_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16460_ _16550_/B _16460_/B vssd1 vssd1 vccd1 vccd1 _16460_/Y sky130_fd_sc_hd__nand2_1
X_13672_ _13558_/A _13559_/Y _13670_/Y _13770_/B vssd1 vssd1 vccd1 vccd1 _13814_/A
+ sky130_fd_sc_hd__a211oi_2
XFILLER_32_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10884_ _10884_/A _10884_/B vssd1 vssd1 vccd1 vccd1 _10891_/A sky130_fd_sc_hd__xnor2_1
X_15411_ _15140_/Y _15206_/B _14895_/B vssd1 vssd1 vccd1 vccd1 _16334_/A sky130_fd_sc_hd__o21ai_2
X_12623_ _12623_/A _12623_/B vssd1 vssd1 vccd1 vccd1 _12624_/B sky130_fd_sc_hd__or2_1
X_16391_ _16399_/A _16571_/B vssd1 vssd1 vccd1 vccd1 _16391_/Y sky130_fd_sc_hd__nor2_1
XFILLER_31_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15342_ _15342_/A _15661_/A vssd1 vssd1 vccd1 vccd1 _15342_/Y sky130_fd_sc_hd__nand2_1
X_12554_ _11849_/A _12550_/X _12553_/X _16735_/A vssd1 vssd1 vccd1 vccd1 _12555_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_156_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11505_ _11487_/A _11487_/B _11485_/X vssd1 vssd1 vccd1 vccd1 _11527_/B sky130_fd_sc_hd__o21ba_1
XFILLER_8_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_808 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15273_ _15493_/A _16416_/A vssd1 vssd1 vccd1 vccd1 _15578_/B sky130_fd_sc_hd__nor2_1
X_12485_ _12311_/A _12311_/B _12310_/A vssd1 vssd1 vccd1 vccd1 _12519_/A sky130_fd_sc_hd__a21oi_1
XFILLER_138_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17012_ _17012_/A _17012_/B vssd1 vssd1 vccd1 vccd1 _17013_/A sky130_fd_sc_hd__nor2_1
XFILLER_7_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14224_ _14680_/A _14599_/B _14485_/D _14426_/D vssd1 vssd1 vccd1 vccd1 _14225_/B
+ sky130_fd_sc_hd__and4_1
X_11436_ _11436_/A _11436_/B vssd1 vssd1 vccd1 vccd1 _11442_/A sky130_fd_sc_hd__xnor2_1
XFILLER_7_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14155_ _14155_/A _14485_/D vssd1 vssd1 vccd1 vccd1 _14156_/B sky130_fd_sc_hd__nand2_1
X_11367_ _11367_/A _11448_/A _11367_/C vssd1 vssd1 vccd1 vccd1 _11403_/A sky130_fd_sc_hd__or3_1
XFILLER_153_874 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13106_ _13106_/A _13106_/B vssd1 vssd1 vccd1 vccd1 _13109_/A sky130_fd_sc_hd__xor2_1
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10318_ _10157_/Y _10230_/X _10263_/X _10283_/X vssd1 vssd1 vccd1 vccd1 _10319_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_3_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14086_ _14087_/B _14086_/B vssd1 vssd1 vccd1 vccd1 _14088_/A sky130_fd_sc_hd__nand2b_1
X_11298_ _11153_/C _11235_/X _11290_/Y _11296_/Y vssd1 vssd1 vccd1 vccd1 _11299_/C
+ sky130_fd_sc_hd__o211a_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13037_ _13302_/A _13037_/B vssd1 vssd1 vccd1 vccd1 _13038_/B sky130_fd_sc_hd__nand2_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10249_ _10262_/A vssd1 vssd1 vccd1 vccd1 _10249_/Y sky130_fd_sc_hd__inv_2
XFILLER_140_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_696 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14988_ _15100_/A _14988_/B vssd1 vssd1 vccd1 vccd1 _14988_/Y sky130_fd_sc_hd__nand2_1
XFILLER_75_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16727_ _16728_/B _16727_/B vssd1 vssd1 vccd1 vccd1 _16794_/B sky130_fd_sc_hd__nand2b_1
X_13939_ wire116/X vssd1 vssd1 vccd1 vccd1 _13939_/Y sky130_fd_sc_hd__inv_2
XFILLER_19_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16658_ _17070_/B _16641_/Y _16648_/X _16657_/X vssd1 vssd1 vccd1 vccd1 _16658_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_34_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15609_ _15609_/A _15609_/B _15609_/C vssd1 vssd1 vccd1 vccd1 _15610_/B sky130_fd_sc_hd__nor3_1
X_16589_ _16812_/A _16589_/B _16743_/C _17043_/B vssd1 vssd1 vccd1 vccd1 _16686_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_50_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09130_ _09139_/B _09130_/B vssd1 vssd1 vccd1 vccd1 _09137_/B sky130_fd_sc_hd__nor2_1
XFILLER_31_972 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09061_ _09061_/A _09298_/A vssd1 vssd1 vccd1 vccd1 _09063_/B sky130_fd_sc_hd__nor2_1
XFILLER_8_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_524 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09963_ _09923_/A _09957_/A _09964_/A _09962_/X vssd1 vssd1 vccd1 vccd1 _10091_/A
+ sky130_fd_sc_hd__a211oi_1
XFILLER_89_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08914_ _17383_/A _12079_/B _09058_/C _17385_/A vssd1 vssd1 vccd1 vccd1 _08914_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_134_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09894_ _09895_/A _09893_/Y _09894_/C _10299_/D vssd1 vssd1 vccd1 vccd1 _10021_/A
+ sky130_fd_sc_hd__and4bb_1
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08845_ _08845_/A _08845_/B vssd1 vssd1 vccd1 vccd1 _08907_/A sky130_fd_sc_hd__xnor2_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08776_ _17397_/A _11861_/B _08776_/C vssd1 vssd1 vccd1 vccd1 _08777_/B sky130_fd_sc_hd__and3_1
XFILLER_150_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_891 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09328_ _09328_/A _09451_/A _09328_/C vssd1 vssd1 vccd1 vccd1 _09329_/B sky130_fd_sc_hd__or3_1
XFILLER_167_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_624 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09259_ _09259_/A _09259_/B vssd1 vssd1 vccd1 vccd1 _09338_/A sky130_fd_sc_hd__or2_1
XFILLER_126_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12270_ _12592_/A _12592_/B _12439_/D _12447_/B vssd1 vssd1 vccd1 vccd1 _12271_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_5_637 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11221_ _11221_/A _11221_/B vssd1 vssd1 vccd1 vccd1 _11223_/A sky130_fd_sc_hd__xor2_1
XFILLER_4_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_502 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11152_ _11153_/B _11153_/C _11153_/A vssd1 vssd1 vccd1 vccd1 _11155_/A sky130_fd_sc_hd__o21a_1
XFILLER_136_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10103_ _10057_/A _10057_/C _10057_/B vssd1 vssd1 vccd1 vccd1 _10194_/B sky130_fd_sc_hd__a21oi_1
XFILLER_150_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15960_ _15960_/A _15960_/B vssd1 vssd1 vccd1 vccd1 _15963_/A sky130_fd_sc_hd__xnor2_1
X_11083_ _11064_/X _11071_/Y _11080_/B _11145_/A vssd1 vssd1 vccd1 vccd1 _11084_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_68_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14911_ _12442_/A _14911_/B vssd1 vssd1 vccd1 vccd1 _14911_/X sky130_fd_sc_hd__and2b_1
X_10034_ _10034_/A _10042_/A _10034_/C vssd1 vssd1 vccd1 vccd1 _10035_/B sky130_fd_sc_hd__or3_1
XFILLER_75_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15891_ _15898_/A _16571_/B _16809_/A vssd1 vssd1 vccd1 vccd1 _15891_/X sky130_fd_sc_hd__or3b_1
XFILLER_49_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14842_ _14842_/A1 _14839_/Y _14840_/Y _14841_/Y _11848_/Y vssd1 vssd1 vccd1 vccd1
+ _14842_/X sky130_fd_sc_hd__o32a_1
XFILLER_36_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17561_ fanout952/X _17561_/D vssd1 vssd1 vccd1 vccd1 _17561_/Q sky130_fd_sc_hd__dfxtp_1
X_11985_ _11986_/B _11985_/B vssd1 vssd1 vccd1 vccd1 _11987_/A sky130_fd_sc_hd__and2b_1
X_14773_ _16644_/C _16651_/A vssd1 vssd1 vccd1 vccd1 _16649_/B sky130_fd_sc_hd__or2_1
XFILLER_91_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16512_ _16604_/B _16809_/C vssd1 vssd1 vccd1 vccd1 _16514_/C sky130_fd_sc_hd__nand2_1
XFILLER_56_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10936_ _10936_/A _10936_/B vssd1 vssd1 vccd1 vccd1 _10938_/B sky130_fd_sc_hd__xnor2_1
X_13724_ _13614_/A _13614_/B _13612_/A vssd1 vssd1 vccd1 vccd1 _13726_/B sky130_fd_sc_hd__a21oi_1
X_17492_ fanout943/X _17492_/D vssd1 vssd1 vccd1 vccd1 _17492_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16443_ _16443_/A _16443_/B vssd1 vssd1 vccd1 vccd1 _16457_/A sky130_fd_sc_hd__nand2_1
XFILLER_71_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10867_ _11117_/C _10963_/C vssd1 vssd1 vccd1 vccd1 _14801_/A sky130_fd_sc_hd__and2_1
X_13655_ _13654_/B _13655_/B vssd1 vssd1 vccd1 vccd1 _13656_/B sky130_fd_sc_hd__nand2b_1
XFILLER_90_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12606_ _12607_/A _12607_/B _12607_/C vssd1 vssd1 vccd1 vccd1 _12778_/A sky130_fd_sc_hd__o21ai_1
X_16374_ _16375_/B _16375_/A vssd1 vssd1 vccd1 vccd1 _16470_/A sky130_fd_sc_hd__nand2b_1
XPHY_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13586_ _13586_/A _13586_/B _13586_/C vssd1 vssd1 vccd1 vccd1 _13587_/B sky130_fd_sc_hd__nor3_1
XFILLER_31_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10798_ _14787_/A _15381_/A vssd1 vssd1 vccd1 vccd1 _10800_/C sky130_fd_sc_hd__and2_1
XPHY_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15325_ _16021_/A _15147_/A _15147_/D _15270_/B vssd1 vssd1 vccd1 vccd1 _15325_/X
+ sky130_fd_sc_hd__a211o_1
X_12537_ _12366_/A _12366_/B _12368_/B _12370_/A _12370_/B vssd1 vssd1 vccd1 vccd1
+ _12540_/B sky130_fd_sc_hd__o32ai_4
XFILLER_118_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12468_ _12662_/B _12468_/B vssd1 vssd1 vccd1 vccd1 _12474_/A sky130_fd_sc_hd__nor2_1
XFILLER_8_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15256_ _16012_/S _17143_/A1 _12553_/B _14962_/B _15255_/X vssd1 vssd1 vccd1 vccd1
+ _15256_/X sky130_fd_sc_hd__o32a_1
XFILLER_144_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11419_ _11419_/A _11419_/B vssd1 vssd1 vccd1 vccd1 _11703_/A sky130_fd_sc_hd__xnor2_2
X_14207_ _14278_/B _14207_/B vssd1 vssd1 vccd1 vccd1 _14207_/X sky130_fd_sc_hd__or2_1
X_15187_ _11321_/X _15804_/A2 _15184_/X _15186_/X _16869_/C1 vssd1 vssd1 vccd1 vccd1
+ _15188_/B sky130_fd_sc_hd__a2111o_1
X_12399_ _13837_/C _12398_/X _12865_/S vssd1 vssd1 vccd1 vccd1 _12400_/B sky130_fd_sc_hd__mux2_1
XFILLER_141_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14138_ _14138_/A _14138_/B vssd1 vssd1 vccd1 vccd1 _14139_/B sky130_fd_sc_hd__and2_1
XFILLER_140_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14069_ _13978_/A _13980_/B _13978_/B vssd1 vssd1 vccd1 vccd1 _14071_/B sky130_fd_sc_hd__o21ba_1
XFILLER_113_579 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_708 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09113_ _09115_/A _09115_/B _09115_/C vssd1 vssd1 vccd1 vccd1 _09119_/B sky130_fd_sc_hd__o21ai_1
XFILLER_129_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_616 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09044_ _09041_/Y _09044_/B vssd1 vssd1 vccd1 vccd1 _09279_/B sky130_fd_sc_hd__and2b_1
XFILLER_135_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_833 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_310 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout900 fanout904/X vssd1 vssd1 vccd1 vccd1 _17467_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_143_192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout911 _10905_/D vssd1 vssd1 vccd1 vccd1 _11027_/D sky130_fd_sc_hd__buf_4
Xfanout922 _17275_/C1 vssd1 vssd1 vccd1 vccd1 _17284_/C1 sky130_fd_sc_hd__buf_2
X_09946_ _09948_/B _09948_/A vssd1 vssd1 vccd1 vccd1 _09951_/B sky130_fd_sc_hd__and2b_1
XFILLER_104_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout933 fanout935/X vssd1 vssd1 vccd1 vccd1 fanout933/X sky130_fd_sc_hd__buf_2
Xfanout944 fanout948/X vssd1 vssd1 vccd1 vccd1 fanout944/X sky130_fd_sc_hd__buf_2
Xfanout955 fanout956/X vssd1 vssd1 vccd1 vccd1 fanout955/X sky130_fd_sc_hd__buf_2
XFILLER_57_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09877_ _09878_/B _09878_/A vssd1 vssd1 vccd1 vccd1 _09877_/X sky130_fd_sc_hd__and2b_1
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08828_ _08829_/B _08828_/B vssd1 vssd1 vccd1 vccd1 _08830_/A sky130_fd_sc_hd__nand2b_1
XFILLER_100_774 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08759_ _12077_/B _12500_/B vssd1 vssd1 vccd1 vccd1 _08776_/C sky130_fd_sc_hd__and2_4
XTAP_2625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_12 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11770_ _10583_/A _11771_/B _11771_/A vssd1 vssd1 vccd1 vccd1 _11770_/Y sky130_fd_sc_hd__a21boi_1
XTAP_2669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10721_ _10722_/B _10722_/A vssd1 vssd1 vccd1 vccd1 _10721_/X sky130_fd_sc_hd__and2b_1
XTAP_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13440_ _13442_/A _13442_/B vssd1 vssd1 vccd1 vccd1 _13441_/A sky130_fd_sc_hd__and2b_1
X_10652_ _10653_/B _10653_/C _10653_/A vssd1 vssd1 vccd1 vccd1 _10662_/A sky130_fd_sc_hd__a21o_1
XFILLER_70_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13371_ _13240_/Y _13244_/B _13496_/A _13370_/Y vssd1 vssd1 vccd1 vccd1 _13496_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_166_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10583_ _10583_/A _10583_/B vssd1 vssd1 vccd1 vccd1 _16972_/A sky130_fd_sc_hd__and2_1
XFILLER_167_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15110_ _15110_/A _15110_/B vssd1 vssd1 vccd1 vccd1 _15110_/Y sky130_fd_sc_hd__nor2_1
XFILLER_10_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12322_ _12323_/A _12492_/A _12323_/C vssd1 vssd1 vccd1 vccd1 _12324_/A sky130_fd_sc_hd__o21a_1
XFILLER_70_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16090_ _15984_/A _15984_/B _15975_/Y vssd1 vssd1 vccd1 vccd1 _16092_/B sky130_fd_sc_hd__a21bo_1
XFILLER_103_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15041_ _11518_/A _15373_/B _15274_/A vssd1 vssd1 vccd1 vccd1 _15041_/X sky130_fd_sc_hd__a21o_1
XFILLER_170_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12253_ _12089_/A _12091_/B _12089_/B vssd1 vssd1 vccd1 vccd1 _12263_/A sky130_fd_sc_hd__o21ba_1
XFILLER_119_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11204_ _11204_/A _11204_/B vssd1 vssd1 vccd1 vccd1 _11205_/B sky130_fd_sc_hd__nand2_1
XFILLER_123_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12184_ _12351_/A _12351_/B vssd1 vssd1 vccd1 vccd1 _12186_/A sky130_fd_sc_hd__xnor2_1
XFILLER_69_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11135_ _11281_/A _14893_/B _11135_/C vssd1 vssd1 vccd1 vccd1 _11137_/C sky130_fd_sc_hd__and3_1
XFILLER_122_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16992_ _17083_/A _16991_/C _16991_/D _16991_/B vssd1 vssd1 vccd1 vccd1 _16993_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_1_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11066_ _11065_/B _11065_/Y _11055_/X _11056_/Y vssd1 vssd1 vccd1 vccd1 _11069_/B
+ sky130_fd_sc_hd__a211oi_2
X_15943_ _15944_/A _15944_/B vssd1 vssd1 vccd1 vccd1 _16080_/A sky130_fd_sc_hd__nor2_1
XFILLER_48_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10017_ _10017_/A _10140_/A vssd1 vssd1 vccd1 vccd1 _10019_/B sky130_fd_sc_hd__nor2_1
XFILLER_37_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15874_ _15989_/B _15874_/B vssd1 vssd1 vccd1 vccd1 _15875_/B sky130_fd_sc_hd__nor2_1
XFILLER_36_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17613_ fanout954/X _17613_/D vssd1 vssd1 vccd1 vccd1 _17613_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14825_ _17023_/B _17024_/A vssd1 vssd1 vccd1 vccd1 _14825_/Y sky130_fd_sc_hd__nand2_1
XFILLER_17_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17544_ fanout956/X _17544_/D vssd1 vssd1 vccd1 vccd1 _17544_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_45_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14756_ _14756_/A1 _14754_/Y _14755_/X _14734_/Y _14735_/X vssd1 vssd1 vccd1 vccd1
+ _17605_/D sky130_fd_sc_hd__a32o_1
XFILLER_91_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11968_ _17405_/A _12166_/B vssd1 vssd1 vccd1 vccd1 _11970_/B sky130_fd_sc_hd__nand2_1
XFILLER_91_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13707_ _13707_/A _13707_/B vssd1 vssd1 vccd1 vccd1 _13707_/X sky130_fd_sc_hd__or2_1
X_17475_ fanout955/X _17608_/Q vssd1 vssd1 vccd1 vccd1 _17475_/Q sky130_fd_sc_hd__dfxtp_1
X_10919_ _14788_/A _10971_/B vssd1 vssd1 vccd1 vccd1 _10924_/A sky130_fd_sc_hd__nand2_1
X_11899_ _17383_/A _12258_/B _11900_/D _17385_/A vssd1 vssd1 vccd1 vccd1 _11901_/A
+ sky130_fd_sc_hd__a22oi_1
X_14687_ _14688_/A _14688_/B vssd1 vssd1 vccd1 vccd1 _14717_/A sky130_fd_sc_hd__or2_1
XFILLER_149_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16426_ _16527_/A _16426_/B vssd1 vssd1 vccd1 vccd1 _16439_/A sky130_fd_sc_hd__nand2b_1
X_13638_ _13638_/A _13638_/B _13638_/C vssd1 vssd1 vccd1 vccd1 _13749_/A sky130_fd_sc_hd__nand3_1
X_16357_ _16358_/A _16358_/B _16358_/C vssd1 vssd1 vccd1 vccd1 _16443_/A sky130_fd_sc_hd__o21ai_1
XFILLER_146_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13569_ _13569_/A _13569_/B _13569_/C vssd1 vssd1 vccd1 vccd1 _13571_/A sky130_fd_sc_hd__or3_1
XFILLER_74_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15308_ _15307_/A _15307_/B _15307_/C vssd1 vssd1 vccd1 vccd1 _15309_/A sky130_fd_sc_hd__o21a_1
X_16288_ _16288_/A _16288_/B vssd1 vssd1 vccd1 vccd1 _16290_/C sky130_fd_sc_hd__xnor2_1
XFILLER_145_479 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15239_ _15175_/X _15176_/Y _15174_/Y vssd1 vssd1 vccd1 vccd1 _15241_/C sky130_fd_sc_hd__a21bo_1
XFILLER_126_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_94 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09800_ _09801_/B _09941_/A _09801_/A vssd1 vssd1 vccd1 vccd1 _09805_/B sky130_fd_sc_hd__o21a_1
Xfanout207 _12046_/A vssd1 vssd1 vccd1 vccd1 _14912_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_119_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout218 _16021_/B vssd1 vssd1 vccd1 vccd1 _16054_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_86_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout229 _14931_/X vssd1 vssd1 vccd1 vccd1 _17163_/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_101_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09731_ _09731_/A _09872_/A vssd1 vssd1 vccd1 vccd1 _09733_/B sky130_fd_sc_hd__nor2_1
XFILLER_39_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09662_ _09662_/A _09662_/B vssd1 vssd1 vccd1 vccd1 _09774_/B sky130_fd_sc_hd__nor2_1
XFILLER_83_912 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09593_ _09580_/X _09581_/Y _09588_/X _09723_/A vssd1 vssd1 vccd1 vccd1 _09597_/A
+ sky130_fd_sc_hd__a211o_1
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1047 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09027_ _09027_/A _09027_/B _09033_/B vssd1 vssd1 vccd1 vccd1 _09048_/B sky130_fd_sc_hd__or3_1
XFILLER_151_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout730 _17496_/Q vssd1 vssd1 vccd1 vccd1 _12077_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_133_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout741 _17495_/Q vssd1 vssd1 vccd1 vccd1 _10171_/D sky130_fd_sc_hd__buf_4
XFILLER_77_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout752 _12334_/B vssd1 vssd1 vccd1 vccd1 _11861_/B sky130_fd_sc_hd__buf_4
X_09929_ _09929_/A _10184_/A vssd1 vssd1 vccd1 vccd1 _09930_/C sky130_fd_sc_hd__nor2_1
XFILLER_120_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout763 _12328_/B vssd1 vssd1 vccd1 vccd1 _11859_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_59_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout774 _17491_/Q vssd1 vssd1 vccd1 vccd1 _12637_/D sky130_fd_sc_hd__clkbuf_2
Xfanout785 fanout795/X vssd1 vssd1 vccd1 vccd1 _12487_/D sky130_fd_sc_hd__buf_2
XFILLER_59_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout796 fanout805/X vssd1 vssd1 vccd1 vccd1 _13194_/D sky130_fd_sc_hd__buf_2
XFILLER_92_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12940_ _12780_/A _12779_/B _12779_/A vssd1 vssd1 vccd1 vccd1 _12981_/A sky130_fd_sc_hd__o21ba_1
XFILLER_58_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12871_ _12871_/A _12871_/B vssd1 vssd1 vccd1 vccd1 _12872_/B sky130_fd_sc_hd__nand2_1
XTAP_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14610_ _14683_/A _14610_/B vssd1 vssd1 vccd1 vccd1 _14612_/B sky130_fd_sc_hd__nor2_1
XTAP_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11822_ _11820_/Y _11821_/X _13516_/S vssd1 vssd1 vccd1 vccd1 _11822_/X sky130_fd_sc_hd__mux2_1
XTAP_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15590_ _15590_/A _15590_/B _15590_/C vssd1 vssd1 vccd1 vccd1 _15591_/B sky130_fd_sc_hd__and3_1
XTAP_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11753_ _11753_/A _11753_/B _11753_/C vssd1 vssd1 vccd1 vccd1 _11759_/A sky130_fd_sc_hd__and3_2
XFILLER_14_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14541_ _14421_/S _14735_/A1 _11820_/A _14636_/A vssd1 vssd1 vccd1 vccd1 _14541_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_81_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10704_ _10904_/A _11005_/B _10805_/D _10954_/A vssd1 vssd1 vccd1 vccd1 _10705_/B
+ sky130_fd_sc_hd__a22oi_1
XTAP_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17260_ _17454_/Q _17290_/A2 _17258_/X _17259_/X _17293_/C1 vssd1 vssd1 vccd1 vccd1
+ _17454_/D sky130_fd_sc_hd__o221a_1
XFILLER_159_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11684_ _15235_/A _15235_/C vssd1 vssd1 vccd1 vccd1 _15302_/A sky130_fd_sc_hd__nor2_1
X_14472_ _14531_/B _14472_/B vssd1 vssd1 vccd1 vccd1 _14473_/C sky130_fd_sc_hd__or2_1
XTAP_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16211_ _16107_/Y _16111_/B _16210_/B vssd1 vssd1 vccd1 vccd1 _16300_/B sky130_fd_sc_hd__o21ba_1
XFILLER_139_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10635_ _10614_/X _10632_/B _10634_/Y _10550_/X vssd1 vssd1 vccd1 vccd1 _10670_/A
+ sky130_fd_sc_hd__a211o_1
X_13423_ _13545_/A _13423_/B _13423_/C vssd1 vssd1 vccd1 vccd1 _13545_/B sky130_fd_sc_hd__nand3_1
X_17191_ _17191_/A _17191_/B _17191_/C _17191_/D vssd1 vssd1 vccd1 vccd1 _17196_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_128_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16142_ _16142_/A _16142_/B vssd1 vssd1 vccd1 vccd1 _16143_/B sky130_fd_sc_hd__and2_1
XFILLER_127_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13354_ _14155_/A _13866_/D vssd1 vssd1 vccd1 vccd1 _13355_/B sky130_fd_sc_hd__nand2_1
XFILLER_6_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10566_ _10566_/A _10566_/B _10566_/C vssd1 vssd1 vccd1 vccd1 _10567_/B sky130_fd_sc_hd__and3_1
XFILLER_143_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12305_ _12305_/A _12305_/B _12305_/C vssd1 vssd1 vccd1 vccd1 _12306_/B sky130_fd_sc_hd__and3_1
X_16073_ _16188_/A _16073_/B vssd1 vssd1 vccd1 vccd1 _16075_/B sky130_fd_sc_hd__nor2_1
X_13285_ _13285_/A _13285_/B vssd1 vssd1 vccd1 vccd1 _13292_/A sky130_fd_sc_hd__xnor2_1
X_10497_ _10497_/A _10497_/B vssd1 vssd1 vccd1 vccd1 _10589_/B sky130_fd_sc_hd__xnor2_1
XFILLER_108_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12236_ _12236_/A _12236_/B vssd1 vssd1 vccd1 vccd1 _12238_/A sky130_fd_sc_hd__nor2_1
X_15024_ _14874_/X _14878_/X _15147_/D vssd1 vssd1 vccd1 vccd1 _15024_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_142_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12167_ _12167_/A _12167_/B vssd1 vssd1 vccd1 vccd1 _12169_/C sky130_fd_sc_hd__xor2_1
XFILLER_110_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11118_ _11118_/A _11246_/A vssd1 vssd1 vccd1 vccd1 _11126_/A sky130_fd_sc_hd__nor2_1
XFILLER_122_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12098_ _12268_/A _12098_/B _12098_/C vssd1 vssd1 vccd1 vccd1 _12268_/B sky130_fd_sc_hd__nand3_2
X_16975_ _14767_/Y _14929_/X _17163_/A2 _16970_/A _16974_/Y vssd1 vssd1 vccd1 vccd1
+ _16977_/B sky130_fd_sc_hd__o221a_1
X_11049_ _11049_/A _11049_/B _11049_/C vssd1 vssd1 vccd1 vccd1 _11051_/C sky130_fd_sc_hd__or3_1
X_15926_ _15926_/A _15926_/B vssd1 vssd1 vccd1 vccd1 _15927_/B sky130_fd_sc_hd__nand2_1
XFILLER_37_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput7 i_wb_addr[13] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__clkbuf_1
XFILLER_65_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_271 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15857_ _15858_/A _15858_/B vssd1 vssd1 vccd1 vccd1 _15857_/X sky130_fd_sc_hd__or2_1
XFILLER_36_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_786 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14808_ _15622_/B _15623_/A _10269_/X vssd1 vssd1 vccd1 vccd1 _15707_/C sky130_fd_sc_hd__a21o_1
XFILLER_52_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15788_ _15788_/A _15788_/B vssd1 vssd1 vccd1 vccd1 _15788_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_17_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17527_ fanout944/X _17527_/D vssd1 vssd1 vccd1 vccd1 _17527_/Q sky130_fd_sc_hd__dfxtp_4
X_14739_ _17167_/A _14739_/B vssd1 vssd1 vccd1 vccd1 _14739_/Y sky130_fd_sc_hd__nand2_1
XFILLER_44_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17458_ fanout934/X _17458_/D vssd1 vssd1 vccd1 vccd1 _17458_/Q sky130_fd_sc_hd__dfxtp_2
X_16409_ _16410_/A _16595_/B vssd1 vssd1 vccd1 vccd1 _16503_/A sky130_fd_sc_hd__nor2_1
X_17389_ _17389_/A _17389_/B vssd1 vssd1 vccd1 vccd1 _17389_/X sky130_fd_sc_hd__or2_1
XFILLER_146_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_592 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09714_ _16982_/B _09710_/Y _09713_/X vssd1 vssd1 vccd1 vccd1 _09852_/B sky130_fd_sc_hd__o21a_1
XFILLER_56_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09645_ _09645_/A _09645_/B _09793_/A vssd1 vssd1 vccd1 vccd1 _09646_/B sky130_fd_sc_hd__nor3_1
XFILLER_16_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09576_ _09576_/A _09721_/A vssd1 vssd1 vccd1 vccd1 _09596_/B sky130_fd_sc_hd__nand2_1
XFILLER_71_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_639 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10420_ _10419_/B _10534_/D _10647_/D _14789_/A vssd1 vssd1 vccd1 vccd1 _10420_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_167_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_552 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10351_ _10345_/A _10343_/Y _10070_/A _10072_/Y vssd1 vssd1 vccd1 vccd1 _10581_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_124_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13070_ _13070_/A _13070_/B vssd1 vssd1 vccd1 vccd1 _13072_/C sky130_fd_sc_hd__xnor2_1
X_10282_ _10134_/Y _10231_/X _10249_/Y _10262_/X vssd1 vssd1 vccd1 vccd1 _10283_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_133_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12021_ _17363_/A _14863_/B vssd1 vssd1 vccd1 vccd1 _14952_/B sky130_fd_sc_hd__and2_1
XFILLER_2_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_780 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_493 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout560 _17514_/Q vssd1 vssd1 vccd1 vccd1 _09899_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_116_94 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout571 _11470_/A vssd1 vssd1 vccd1 vccd1 _15715_/A sky130_fd_sc_hd__buf_4
X_16760_ _16760_/A _16760_/B vssd1 vssd1 vccd1 vccd1 _16761_/B sky130_fd_sc_hd__nand2_1
Xfanout582 _10180_/A vssd1 vssd1 vccd1 vccd1 _16011_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_120_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13972_ _14058_/B _13972_/B vssd1 vssd1 vccd1 vccd1 _13974_/A sky130_fd_sc_hd__nand2_1
XFILLER_59_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout593 _14954_/A vssd1 vssd1 vccd1 vccd1 _15095_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_58_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15711_ _15805_/A _15711_/B vssd1 vssd1 vccd1 vccd1 _15711_/Y sky130_fd_sc_hd__nor2_1
X_12923_ _14213_/A _14050_/B _13067_/D _12923_/D vssd1 vssd1 vccd1 vccd1 _12924_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_20_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16691_ _16601_/A _16614_/B _16601_/B vssd1 vssd1 vccd1 vccd1 _16693_/B sky130_fd_sc_hd__a21boi_1
XFILLER_132_60 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_775 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15642_ _16226_/C _16812_/A _16591_/B _15726_/A vssd1 vssd1 vccd1 vccd1 _15643_/B
+ sky130_fd_sc_hd__a22o_1
XTAP_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12854_ _14636_/A _13626_/B vssd1 vssd1 vccd1 vccd1 _14758_/A sky130_fd_sc_hd__nand2_1
XFILLER_74_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11805_ _11802_/Y _11804_/Y _17365_/A vssd1 vssd1 vccd1 vccd1 _11805_/X sky130_fd_sc_hd__mux2_1
XTAP_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15573_ _15573_/A _15573_/B vssd1 vssd1 vccd1 vccd1 _15584_/A sky130_fd_sc_hd__xnor2_1
XTAP_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12785_ _12655_/A _12655_/B _12671_/B _12670_/B _12670_/A vssd1 vssd1 vccd1 vccd1
+ _12822_/B sky130_fd_sc_hd__a32o_1
XTAP_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17312_ _12618_/D _17322_/A2 _17311_/X _17378_/C1 vssd1 vssd1 vccd1 vccd1 _17485_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14524_ _14524_/A _14524_/B _14524_/C vssd1 vssd1 vccd1 vccd1 _14583_/A sky130_fd_sc_hd__or3_1
XFILLER_70_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11736_ _11736_/A _11736_/B _11735_/Y vssd1 vssd1 vccd1 vccd1 _11739_/B sky130_fd_sc_hd__nor3b_1
XFILLER_15_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17243_ _17590_/Q _17273_/A2 _17273_/B1 vssd1 vssd1 vccd1 vccd1 _17243_/X sky130_fd_sc_hd__a21o_1
XFILLER_30_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14455_ _14509_/C _14455_/B vssd1 vssd1 vccd1 vccd1 _14456_/C sky130_fd_sc_hd__and2_1
X_11667_ _11686_/B _11686_/A vssd1 vssd1 vccd1 vccd1 _11690_/A sky130_fd_sc_hd__and2b_1
X_13406_ _13406_/A _13406_/B vssd1 vssd1 vccd1 vccd1 _13408_/A sky130_fd_sc_hd__nor2_1
XFILLER_174_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10618_ _10963_/A _10963_/B _10875_/C _10962_/B vssd1 vssd1 vccd1 vccd1 _10621_/A
+ sky130_fd_sc_hd__and4_1
X_17174_ input19/X input22/X input21/X input23/X vssd1 vssd1 vccd1 vccd1 _17181_/B
+ sky130_fd_sc_hd__or4b_1
XFILLER_167_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11598_ _11598_/A _11598_/B vssd1 vssd1 vccd1 vccd1 _11639_/A sky130_fd_sc_hd__xor2_1
XFILLER_128_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14386_ _14386_/A _14386_/B vssd1 vssd1 vccd1 vccd1 _14388_/A sky130_fd_sc_hd__nor2_1
XFILLER_155_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16125_ _16125_/A vssd1 vssd1 vccd1 vccd1 _17558_/D sky130_fd_sc_hd__clkinv_2
X_13337_ _13337_/A _13455_/A _13337_/C vssd1 vssd1 vccd1 vccd1 _13455_/B sky130_fd_sc_hd__nor3_1
X_10549_ _10671_/A _10549_/B vssd1 vssd1 vccd1 vccd1 _10550_/C sky130_fd_sc_hd__and2_1
XFILLER_170_511 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16056_ _16056_/A _16259_/B _16454_/A vssd1 vssd1 vccd1 vccd1 _16058_/A sky130_fd_sc_hd__and3_1
XFILLER_115_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13268_ _13268_/A _13268_/B vssd1 vssd1 vccd1 vccd1 _13511_/A sky130_fd_sc_hd__nor2_1
XFILLER_124_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15007_ _11675_/C _11655_/A _14793_/Y _15108_/A _15006_/Y vssd1 vssd1 vccd1 vccd1
+ _15007_/X sky130_fd_sc_hd__o311a_1
XFILLER_29_1043 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12219_ _12213_/X _12218_/Y _13833_/S vssd1 vssd1 vccd1 vccd1 _12219_/X sky130_fd_sc_hd__mux2_1
XFILLER_69_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13199_ _13199_/A _13199_/B _13199_/C vssd1 vssd1 vccd1 vccd1 _13200_/B sky130_fd_sc_hd__nor3_1
XFILLER_116_1002 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16958_ _16958_/A _16958_/B vssd1 vssd1 vccd1 vccd1 _17012_/B sky130_fd_sc_hd__xor2_1
XFILLER_37_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_580 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15909_ _15884_/Y _15885_/Y _15884_/A vssd1 vssd1 vccd1 vccd1 _15994_/A sky130_fd_sc_hd__o21ai_2
X_16889_ _16888_/A _16888_/B _16888_/C vssd1 vssd1 vccd1 vccd1 _16952_/A sky130_fd_sc_hd__a21o_1
XFILLER_80_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09430_ _09427_/Y _09430_/B vssd1 vssd1 vccd1 vccd1 _09563_/B sky130_fd_sc_hd__and2b_1
XFILLER_25_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09361_ _09360_/A _09502_/B _09502_/C vssd1 vssd1 vccd1 vccd1 _09361_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_52_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09292_ _09292_/A _09437_/A vssd1 vssd1 vccd1 vccd1 _09310_/B sky130_fd_sc_hd__nand2_1
XFILLER_36_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_12 _17023_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_23 _17529_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_34 _17546_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_45 _13302_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_56 _10308_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_67 _12770_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_78 _15715_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_89 fanout699/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09628_ _09628_/A _09628_/B _09628_/C vssd1 vssd1 vccd1 vccd1 _09668_/A sky130_fd_sc_hd__or3_2
XFILLER_71_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_756 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09559_ _09559_/A _09559_/B vssd1 vssd1 vccd1 vccd1 _09689_/B sky130_fd_sc_hd__xnor2_1
XFILLER_169_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12570_ _12570_/A _12570_/B vssd1 vssd1 vccd1 vccd1 _12572_/C sky130_fd_sc_hd__xor2_1
XFILLER_52_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_806 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11521_ _11521_/A _11565_/A vssd1 vssd1 vccd1 vccd1 _11523_/B sky130_fd_sc_hd__nor2_1
XFILLER_157_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11452_ _11453_/A _11453_/B vssd1 vssd1 vccd1 vccd1 _11460_/A sky130_fd_sc_hd__or2_1
X_14240_ _13893_/A _14433_/B _14366_/B _14318_/A vssd1 vssd1 vccd1 vccd1 _14242_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10403_ _10402_/A _10402_/B _10402_/C vssd1 vssd1 vccd1 vccd1 _10405_/C sky130_fd_sc_hd__a21oi_1
X_14171_ _14171_/A _14245_/B vssd1 vssd1 vccd1 vccd1 _14173_/C sky130_fd_sc_hd__nor2_1
X_11383_ _11395_/B _11383_/B _11383_/C vssd1 vssd1 vccd1 vccd1 _11435_/A sky130_fd_sc_hd__nand3_2
XFILLER_164_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13122_ _13121_/A _13121_/B _13121_/C vssd1 vssd1 vccd1 vccd1 _13123_/B sky130_fd_sc_hd__o21a_1
X_10334_ _10451_/A _10334_/B vssd1 vssd1 vccd1 vccd1 _10336_/B sky130_fd_sc_hd__xnor2_1
XFILLER_124_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13053_ _12907_/A _13948_/C _12908_/A _12905_/X vssd1 vssd1 vccd1 vccd1 _13055_/B
+ sky130_fd_sc_hd__a31oi_1
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10265_ _10265_/A _10265_/B vssd1 vssd1 vccd1 vccd1 _10267_/C sky130_fd_sc_hd__xnor2_1
XFILLER_79_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12004_ _12200_/B _12004_/B vssd1 vssd1 vccd1 vccd1 _12007_/A sky130_fd_sc_hd__nor2_1
XFILLER_121_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10196_ _10321_/A _09172_/B _10062_/B _09514_/B vssd1 vssd1 vccd1 vccd1 _10198_/C
+ sky130_fd_sc_hd__a22oi_1
XFILLER_120_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16812_ _16812_/A _16883_/A _16938_/D _16883_/C vssd1 vssd1 vccd1 vccd1 _16816_/A
+ sky130_fd_sc_hd__or4b_1
XFILLER_78_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout390 _14772_/A vssd1 vssd1 vccd1 vccd1 _16723_/A sky130_fd_sc_hd__buf_4
XFILLER_93_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16743_ _16814_/B _16743_/B _16743_/C _17043_/B vssd1 vssd1 vccd1 vccd1 _16744_/B
+ sky130_fd_sc_hd__and4_1
X_13955_ _14134_/A _13955_/B vssd1 vssd1 vccd1 vccd1 _13958_/C sky130_fd_sc_hd__and2_1
XFILLER_35_904 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12906_ _12749_/Y _13182_/C _12905_/X vssd1 vssd1 vccd1 vccd1 _12908_/A sky130_fd_sc_hd__a21oi_1
X_16674_ _16751_/B _16674_/B vssd1 vssd1 vccd1 vccd1 _16677_/B sky130_fd_sc_hd__nand2_1
XFILLER_47_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13886_ _13779_/B _13781_/B _13779_/A vssd1 vssd1 vccd1 vccd1 _13888_/B sky130_fd_sc_hd__o21ba_1
XFILLER_62_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15625_ _10269_/X _15804_/A2 _15713_/B1 _15624_/A vssd1 vssd1 vccd1 vccd1 _15625_/X
+ sky130_fd_sc_hd__a22o_1
X_12837_ _12833_/Y _12835_/X _12651_/A _12655_/A vssd1 vssd1 vccd1 vccd1 _12837_/Y
+ sky130_fd_sc_hd__o211ai_1
XFILLER_61_244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15556_ _16226_/B _16152_/A vssd1 vssd1 vccd1 vccd1 _15557_/B sky130_fd_sc_hd__nand2_1
XTAP_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12768_ _12765_/Y _12920_/B _12612_/A _12612_/Y vssd1 vssd1 vccd1 vccd1 _12782_/B
+ sky130_fd_sc_hd__a211o_1
XTAP_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14507_ _14508_/A _14508_/B vssd1 vssd1 vccd1 vccd1 _14569_/A sky130_fd_sc_hd__nand2b_1
XFILLER_147_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11719_ _11719_/A _11719_/B vssd1 vssd1 vccd1 vccd1 _11726_/B sky130_fd_sc_hd__and2_1
X_15487_ _15406_/A _15406_/B _15403_/X vssd1 vssd1 vccd1 vccd1 _15489_/B sky130_fd_sc_hd__a21o_1
X_12699_ _13003_/A _12698_/B _15998_/A vssd1 vssd1 vccd1 vccd1 _12699_/X sky130_fd_sc_hd__a21o_1
XFILLER_174_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17226_ _17552_/Q _17274_/B vssd1 vssd1 vccd1 vccd1 _17226_/X sky130_fd_sc_hd__and2_1
Xinput10 i_wb_addr[16] vssd1 vssd1 vccd1 vccd1 input10/X sky130_fd_sc_hd__clkbuf_1
X_14438_ _14438_/A _14438_/B vssd1 vssd1 vccd1 vccd1 _14440_/C sky130_fd_sc_hd__nor2_1
Xinput21 i_wb_addr[26] vssd1 vssd1 vccd1 vccd1 input21/X sky130_fd_sc_hd__clkbuf_1
XFILLER_122_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput32 i_wb_addr[7] vssd1 vssd1 vccd1 vccd1 input32/X sky130_fd_sc_hd__clkbuf_1
XFILLER_128_552 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput43 i_wb_data[16] vssd1 vssd1 vccd1 vccd1 input43/X sky130_fd_sc_hd__clkbuf_1
Xinput54 i_wb_data[26] vssd1 vssd1 vccd1 vccd1 input54/X sky130_fd_sc_hd__clkbuf_1
XFILLER_128_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17157_ _17138_/A _17138_/B _10098_/A vssd1 vssd1 vccd1 vccd1 _17157_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_155_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput65 i_wb_data[7] vssd1 vssd1 vccd1 vccd1 input65/X sky130_fd_sc_hd__clkbuf_2
X_14369_ _14554_/A _14433_/B _14368_/C vssd1 vssd1 vccd1 vccd1 _14370_/B sky130_fd_sc_hd__a21oi_1
XFILLER_155_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16108_ _16114_/A _16644_/B _16108_/C vssd1 vssd1 vccd1 vccd1 _16108_/X sky130_fd_sc_hd__and3b_1
X_17088_ _17088_/A _17088_/B _17088_/C vssd1 vssd1 vccd1 vccd1 _17089_/B sky130_fd_sc_hd__nor3_1
XFILLER_171_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16039_ _16416_/A _16681_/A vssd1 vssd1 vccd1 vccd1 _16040_/B sky130_fd_sc_hd__nor2_1
X_08930_ _08930_/A _08930_/B _08930_/C vssd1 vssd1 vccd1 vccd1 _08930_/X sky130_fd_sc_hd__or3_1
XFILLER_88_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08861_ _08861_/A _08861_/B vssd1 vssd1 vccd1 vccd1 _08864_/A sky130_fd_sc_hd__xnor2_1
XFILLER_111_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08792_ _11878_/A _09319_/C _17387_/A _08792_/D vssd1 vssd1 vccd1 vccd1 _11878_/B
+ sky130_fd_sc_hd__and4b_1
XFILLER_84_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09413_ _10242_/A1 _09557_/B _09555_/C _09414_/A vssd1 vssd1 vccd1 vccd1 _09415_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_34_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09344_ _09344_/A _09344_/B _09344_/C vssd1 vssd1 vccd1 vccd1 _09344_/Y sky130_fd_sc_hd__nor3_2
XFILLER_80_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09275_ _09275_/A _09275_/B vssd1 vssd1 vccd1 vccd1 _09404_/B sky130_fd_sc_hd__xnor2_1
XFILLER_138_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_931 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10050_ _10050_/A _10050_/B _10163_/A vssd1 vssd1 vccd1 vccd1 _10053_/B sky130_fd_sc_hd__nand3_1
XFILLER_88_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13740_ _13741_/A _13741_/B _13741_/C vssd1 vssd1 vccd1 vccd1 _13742_/A sky130_fd_sc_hd__o21a_1
XFILLER_44_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10952_ _10953_/A _10953_/B vssd1 vssd1 vccd1 vccd1 _11195_/A sky130_fd_sc_hd__or2_1
XFILLER_17_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13671_ _13671_/A _13671_/B _13671_/C vssd1 vssd1 vccd1 vccd1 _13770_/B sky130_fd_sc_hd__and3_1
X_10883_ _10883_/A _10883_/B _10883_/C vssd1 vssd1 vccd1 vccd1 _10893_/B sky130_fd_sc_hd__nand3_1
X_15410_ _15140_/Y _15206_/B _14895_/B vssd1 vssd1 vccd1 vccd1 _15854_/B sky130_fd_sc_hd__o21a_1
X_12622_ _12623_/A _12623_/B vssd1 vssd1 vccd1 vccd1 _12780_/A sky130_fd_sc_hd__nand2_1
XFILLER_169_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16390_ _14776_/A _16644_/B _16399_/A vssd1 vssd1 vccd1 vccd1 _16390_/Y sky130_fd_sc_hd__a21boi_1
X_15341_ _15493_/A _15755_/B vssd1 vssd1 vccd1 vccd1 _15661_/A sky130_fd_sc_hd__nor2_1
X_12553_ _15457_/B _12553_/B vssd1 vssd1 vccd1 vccd1 _12553_/X sky130_fd_sc_hd__or2_1
XFILLER_169_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11504_ _11499_/A _11499_/C _11499_/B vssd1 vssd1 vccd1 vccd1 _11539_/B sky130_fd_sc_hd__o21a_1
XFILLER_11_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15272_ _15207_/X _15270_/X _11437_/D vssd1 vssd1 vccd1 vccd1 _16595_/A sky130_fd_sc_hd__a21bo_2
X_12484_ _12354_/A _12353_/B _12353_/A vssd1 vssd1 vccd1 vccd1 _12521_/A sky130_fd_sc_hd__a21bo_1
XFILLER_172_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1029 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17011_ _17014_/A _17014_/B vssd1 vssd1 vccd1 vccd1 _17060_/A sky130_fd_sc_hd__nor2_1
XFILLER_8_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14223_ _14599_/B _14485_/D _14426_/D _14680_/A vssd1 vssd1 vccd1 vccd1 _14225_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_171_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11435_ _11435_/A _11435_/B _11435_/C vssd1 vssd1 vccd1 vccd1 _11444_/A sky130_fd_sc_hd__nand3_1
XFILLER_138_883 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11366_ _11341_/A _11341_/B _11341_/C vssd1 vssd1 vccd1 vccd1 _11367_/C sky130_fd_sc_hd__a21oi_1
XFILLER_153_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14154_ _14154_/A _14154_/B vssd1 vssd1 vccd1 vccd1 _14156_/A sky130_fd_sc_hd__nor2_1
XFILLER_153_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13105_ _13106_/B _13106_/A vssd1 vssd1 vccd1 vccd1 _13236_/B sky130_fd_sc_hd__and2b_1
X_10317_ _10330_/A _10287_/Y _10303_/Y _10315_/X vssd1 vssd1 vccd1 vccd1 _10319_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_153_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11297_ _11290_/Y _11296_/Y _11153_/C _11235_/X vssd1 vssd1 vccd1 vccd1 _11299_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_125_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14085_ _16864_/A _16918_/A _13998_/B vssd1 vssd1 vccd1 vccd1 _14086_/B sky130_fd_sc_hd__o21ba_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13036_ _13036_/A _13036_/B vssd1 vssd1 vccd1 vccd1 _13038_/A sky130_fd_sc_hd__nor2_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10248_ _10261_/B _10261_/C _10261_/A vssd1 vssd1 vccd1 vccd1 _10262_/A sky130_fd_sc_hd__a21o_1
XFILLER_79_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10179_ _10430_/A _10431_/B vssd1 vssd1 vccd1 vccd1 _10180_/C sky130_fd_sc_hd__and2_2
XFILLER_94_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14987_ _11841_/B _12054_/B _10657_/B _10308_/B _09925_/A _10182_/C vssd1 vssd1 vccd1
+ vccd1 _14988_/B sky130_fd_sc_hd__mux4_1
XFILLER_47_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16726_ _16568_/A _16568_/B _16641_/A _11762_/X vssd1 vssd1 vccd1 vccd1 _16728_/B
+ sky130_fd_sc_hd__a31oi_1
XFILLER_19_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13938_ _13010_/B _13511_/X _13934_/Y _13935_/Y _13937_/X vssd1 vssd1 vccd1 vccd1
+ wire116/A sky130_fd_sc_hd__a311oi_2
XFILLER_93_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_222 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16657_ _16304_/A _16649_/X _16650_/Y _16652_/X _16656_/X vssd1 vssd1 vccd1 vccd1
+ _16657_/X sky130_fd_sc_hd__o311a_1
X_13869_ _13869_/A _13869_/B vssd1 vssd1 vccd1 vccd1 _13870_/B sky130_fd_sc_hd__xnor2_1
XFILLER_23_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15608_ _15609_/A _15609_/B _15609_/C vssd1 vssd1 vccd1 vccd1 _15610_/A sky130_fd_sc_hd__o21a_1
XFILLER_50_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16588_ _16747_/A _16497_/C _16497_/D _16814_/A vssd1 vssd1 vccd1 vccd1 _16590_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_31_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15539_ _15901_/S _14989_/X _15538_/X _17371_/A vssd1 vssd1 vccd1 vccd1 _15539_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_33_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09060_ _09061_/A _09059_/Y _17381_/A _12079_/B vssd1 vssd1 vccd1 vccd1 _09298_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_163_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17209_ _17437_/Q _17275_/A2 _17207_/X _17208_/X _17364_/C1 vssd1 vssd1 vccd1 vccd1
+ _17437_/D sky130_fd_sc_hd__o221a_1
XFILLER_129_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09962_ _09813_/X _09829_/Y _09960_/A _09960_/Y vssd1 vssd1 vccd1 vccd1 _09962_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_131_536 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08913_ _08913_/A _17383_/A _12079_/B _09058_/C vssd1 vssd1 vccd1 vccd1 _08916_/A
+ sky130_fd_sc_hd__and4_1
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09893_ _09892_/B _10421_/D _10534_/D _09892_/A vssd1 vssd1 vccd1 vccd1 _09893_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_112_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08844_ _08845_/B _08845_/A vssd1 vssd1 vccd1 vccd1 _08844_/X sky130_fd_sc_hd__and2b_1
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08775_ _17397_/A _11861_/B _08776_/C vssd1 vssd1 vccd1 vccd1 _08777_/A sky130_fd_sc_hd__a21oi_1
XTAP_2807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09327_ _09462_/A _09326_/Y _09327_/C _11808_/B vssd1 vssd1 vccd1 vccd1 _09468_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_167_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09258_ _09071_/A _09071_/C _09071_/B vssd1 vssd1 vccd1 vccd1 _09259_/B sky130_fd_sc_hd__o21a_1
XFILLER_167_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09189_ _09189_/A _09221_/A _09189_/C vssd1 vssd1 vccd1 vccd1 _09221_/B sky130_fd_sc_hd__nor3_1
XFILLER_153_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11220_ _11220_/A _11220_/B vssd1 vssd1 vccd1 vccd1 _11221_/B sky130_fd_sc_hd__xnor2_1
XFILLER_5_649 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_330 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_1035 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11151_ _11153_/B _11151_/B _11151_/C vssd1 vssd1 vccd1 vccd1 _11153_/C sky130_fd_sc_hd__nor3_2
XFILLER_135_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10102_ _10086_/A _10086_/C _10086_/B vssd1 vssd1 vccd1 vccd1 _10216_/B sky130_fd_sc_hd__o21ai_1
XFILLER_161_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11082_ _11082_/A _11082_/B vssd1 vssd1 vccd1 vccd1 _11084_/B sky130_fd_sc_hd__xnor2_1
XFILLER_49_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10033_ _10033_/A _10033_/B vssd1 vssd1 vccd1 vccd1 _10055_/A sky130_fd_sc_hd__nor2_1
X_14910_ _17131_/A _15846_/A _15726_/A vssd1 vssd1 vccd1 vccd1 _14910_/X sky130_fd_sc_hd__and3_1
XFILLER_48_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15890_ _16809_/A _16644_/B _15898_/A vssd1 vssd1 vccd1 vccd1 _15890_/X sky130_fd_sc_hd__a21bo_1
XFILLER_76_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14841_ _15457_/B _14841_/B vssd1 vssd1 vccd1 vccd1 _14841_/Y sky130_fd_sc_hd__nor2_1
XFILLER_36_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17560_ fanout951/X _17560_/D vssd1 vssd1 vccd1 vccd1 _17560_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_583 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14772_ _14772_/A _16722_/A vssd1 vssd1 vccd1 vccd1 _16729_/B sky130_fd_sc_hd__or2_1
XFILLER_17_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11984_ _11984_/A _11984_/B vssd1 vssd1 vccd1 vccd1 _11985_/B sky130_fd_sc_hd__xnor2_1
X_16511_ _16511_/A _16511_/B vssd1 vssd1 vccd1 vccd1 _16522_/A sky130_fd_sc_hd__or2_1
XFILLER_44_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13723_ _13723_/A _13723_/B vssd1 vssd1 vccd1 vccd1 _13726_/A sky130_fd_sc_hd__xnor2_1
XFILLER_90_158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10935_ _10935_/A _10935_/B vssd1 vssd1 vccd1 vccd1 _10936_/B sky130_fd_sc_hd__nor2_1
X_17491_ fanout943/X _17491_/D vssd1 vssd1 vccd1 vccd1 _17491_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_56_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16442_ _16442_/A _16442_/B vssd1 vssd1 vccd1 vccd1 _16459_/A sky130_fd_sc_hd__xor2_1
XFILLER_71_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13654_ _13655_/B _13654_/B vssd1 vssd1 vccd1 vccd1 _13654_/X sky130_fd_sc_hd__and2b_1
X_10866_ _11115_/A _11115_/B _11117_/D _11115_/C vssd1 vssd1 vccd1 vccd1 _10870_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_143_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12605_ _12605_/A _12605_/B vssd1 vssd1 vccd1 vccd1 _12607_/C sky130_fd_sc_hd__xnor2_1
X_16373_ _16283_/A _16283_/B _16277_/A vssd1 vssd1 vccd1 vccd1 _16375_/B sky130_fd_sc_hd__o21a_1
XPHY_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13585_ _13586_/A _13586_/B _13586_/C vssd1 vssd1 vccd1 vccd1 _13587_/A sky130_fd_sc_hd__o21a_1
XFILLER_12_450 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10797_ _11117_/C _10875_/C vssd1 vssd1 vccd1 vccd1 _10803_/A sky130_fd_sc_hd__nand2_1
XFILLER_129_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15324_ _16226_/C _16317_/B vssd1 vssd1 vccd1 vccd1 _15350_/A sky130_fd_sc_hd__nand2_1
X_12536_ _12536_/A _12536_/B vssd1 vssd1 vccd1 vccd1 _12540_/A sky130_fd_sc_hd__xnor2_2
XFILLER_173_915 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15255_ _15245_/X _15252_/X _15254_/X _15253_/X _13627_/S _17371_/A vssd1 vssd1 vccd1
+ vccd1 _15255_/X sky130_fd_sc_hd__mux4_1
X_12467_ _12467_/A _12467_/B vssd1 vssd1 vccd1 vccd1 _12468_/B sky130_fd_sc_hd__and2_1
X_14206_ _14278_/B _14207_/B vssd1 vssd1 vccd1 vccd1 _14206_/Y sky130_fd_sc_hd__nand2_1
X_11418_ _11418_/A _11418_/B vssd1 vssd1 vccd1 vccd1 _11708_/B sky130_fd_sc_hd__xnor2_1
X_15186_ _15175_/B _14848_/C _15185_/Y vssd1 vssd1 vccd1 vccd1 _15186_/X sky130_fd_sc_hd__o21a_1
X_12398_ _12040_/Y _12061_/Y _15095_/B vssd1 vssd1 vccd1 vccd1 _12398_/X sky130_fd_sc_hd__mux2_1
XFILLER_140_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14137_ _14138_/A _14138_/B vssd1 vssd1 vccd1 vccd1 _14221_/A sky130_fd_sc_hd__nor2_1
XFILLER_113_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11349_ _11349_/A _11349_/B _11349_/C vssd1 vssd1 vccd1 vccd1 _11402_/A sky130_fd_sc_hd__and3_1
XFILLER_153_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14068_ _14068_/A _14068_/B vssd1 vssd1 vccd1 vccd1 _14071_/A sky130_fd_sc_hd__xnor2_1
XFILLER_113_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13019_ _13019_/A _13019_/B vssd1 vssd1 vccd1 vccd1 _13021_/A sky130_fd_sc_hd__nor2_1
XFILLER_100_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16709_ _16709_/A _16709_/B vssd1 vssd1 vccd1 vccd1 _16711_/C sky130_fd_sc_hd__xnor2_1
XFILLER_62_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09112_ _09092_/A _09314_/B _09093_/A vssd1 vssd1 vccd1 vccd1 _09115_/C sky130_fd_sc_hd__o21a_1
XFILLER_148_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09043_ _09043_/A _17081_/B vssd1 vssd1 vccd1 vccd1 _09044_/B sky130_fd_sc_hd__nand2_1
XFILLER_164_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout901 fanout904/X vssd1 vssd1 vccd1 vccd1 _11240_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_131_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_878 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout912 _17478_/Q vssd1 vssd1 vccd1 vccd1 _10905_/D sky130_fd_sc_hd__clkbuf_4
X_09945_ _09945_/A _10064_/A vssd1 vssd1 vccd1 vccd1 _09948_/B sky130_fd_sc_hd__nor2_1
Xfanout923 _17364_/C1 vssd1 vssd1 vccd1 vccd1 _17275_/C1 sky130_fd_sc_hd__clkbuf_2
Xfanout934 fanout935/X vssd1 vssd1 vccd1 vccd1 fanout934/X sky130_fd_sc_hd__clkbuf_2
Xfanout945 fanout947/X vssd1 vssd1 vccd1 vccd1 fanout945/X sky130_fd_sc_hd__clkbuf_2
Xfanout956 fanout957/X vssd1 vssd1 vccd1 vccd1 fanout956/X sky130_fd_sc_hd__clkbuf_4
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09876_ _09876_/A _10018_/A vssd1 vssd1 vccd1 vccd1 _09878_/B sky130_fd_sc_hd__nor2_1
XFILLER_161_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08827_ _08893_/A _08826_/B _08826_/A vssd1 vssd1 vccd1 vccd1 _08828_/B sky130_fd_sc_hd__o21ba_1
XFILLER_58_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08758_ _12077_/B _13208_/D _13080_/D _12077_/A vssd1 vssd1 vccd1 vccd1 _08758_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_72_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_840 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10720_ _10720_/A _11013_/A vssd1 vssd1 vccd1 vccd1 _10722_/B sky130_fd_sc_hd__nor2_1
XTAP_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10651_ _10653_/B _10653_/C _10653_/A vssd1 vssd1 vccd1 vccd1 _10651_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_110_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13370_ _13369_/B _13369_/C _13369_/A vssd1 vssd1 vccd1 vccd1 _13370_/Y sky130_fd_sc_hd__a21oi_1
X_10582_ _10582_/A _10582_/B vssd1 vssd1 vccd1 vccd1 _10583_/B sky130_fd_sc_hd__nand2_1
XFILLER_70_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12321_ _17409_/A _12637_/D vssd1 vssd1 vccd1 vccd1 _12323_/C sky130_fd_sc_hd__nand2_1
XFILLER_70_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15040_ _16011_/C _15034_/Y _15037_/X _15039_/X _15312_/S _15901_/S vssd1 vssd1 vccd1
+ vccd1 _15040_/X sky130_fd_sc_hd__mux4_1
X_12252_ _12252_/A _12252_/B _12252_/C vssd1 vssd1 vccd1 vccd1 _12265_/B sky130_fd_sc_hd__or3_1
XFILLER_5_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11203_ _11204_/A _11204_/B vssd1 vssd1 vccd1 vccd1 _11739_/A sky130_fd_sc_hd__or2_1
XFILLER_79_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12183_ _12183_/A _12183_/B vssd1 vssd1 vccd1 vccd1 _12351_/B sky130_fd_sc_hd__nor2_1
X_11134_ _11137_/B _11134_/B vssd1 vssd1 vccd1 vccd1 _11135_/C sky130_fd_sc_hd__nor2_1
X_16991_ _17083_/A _16991_/B _16991_/C _16991_/D vssd1 vssd1 vccd1 vccd1 _17046_/B
+ sky130_fd_sc_hd__and4_1
X_11065_ _11065_/A _11065_/B _11065_/C _11065_/D vssd1 vssd1 vccd1 vccd1 _11065_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_135_82 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15942_ _15837_/A _15837_/B _15826_/Y vssd1 vssd1 vccd1 vccd1 _15944_/B sky130_fd_sc_hd__a21oi_1
XFILLER_89_792 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10016_ _10017_/A _10015_/Y _10271_/A _10016_/D vssd1 vssd1 vccd1 vccd1 _10140_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_64_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15873_ _16281_/A _16259_/B _15872_/C vssd1 vssd1 vccd1 vccd1 _15874_/B sky130_fd_sc_hd__a21oi_1
XFILLER_36_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14824_ _14767_/Y _16971_/A _16970_/A vssd1 vssd1 vccd1 vccd1 _17024_/A sky130_fd_sc_hd__o21ai_1
X_17612_ fanout954/X _17612_/D vssd1 vssd1 vccd1 vccd1 _17612_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17543_ fanout954/X _17543_/D vssd1 vssd1 vccd1 vccd1 _17543_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_63_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14755_ _14755_/A _14755_/B vssd1 vssd1 vccd1 vccd1 _14755_/X sky130_fd_sc_hd__or2_1
X_11967_ _11967_/A _11967_/B vssd1 vssd1 vccd1 vccd1 _11970_/A sky130_fd_sc_hd__nand2_1
XFILLER_32_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13706_ _13707_/A _13707_/B vssd1 vssd1 vccd1 vccd1 _13706_/Y sky130_fd_sc_hd__nand2_1
X_17474_ fanout955/X _17607_/Q vssd1 vssd1 vccd1 vccd1 _17474_/Q sky130_fd_sc_hd__dfxtp_1
X_10918_ _10918_/A _10918_/B vssd1 vssd1 vccd1 vccd1 _10926_/A sky130_fd_sc_hd__xnor2_1
XFILLER_44_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14686_ _14719_/A _14686_/B vssd1 vssd1 vccd1 vccd1 _14688_/B sky130_fd_sc_hd__xnor2_1
X_11898_ _12138_/B _11898_/B vssd1 vssd1 vccd1 vccd1 _11908_/A sky130_fd_sc_hd__nor2_1
XFILLER_32_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16425_ _16425_/A _16425_/B _16423_/Y vssd1 vssd1 vccd1 vccd1 _16426_/B sky130_fd_sc_hd__or3b_1
X_13637_ _13637_/A _13637_/B vssd1 vssd1 vccd1 vccd1 _13638_/C sky130_fd_sc_hd__nand2_1
X_10849_ _10850_/A _10850_/C vssd1 vssd1 vccd1 vccd1 _10855_/B sky130_fd_sc_hd__nor2_1
XFILLER_32_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16356_ _16356_/A _16356_/B vssd1 vssd1 vccd1 vccd1 _16358_/C sky130_fd_sc_hd__xnor2_1
XFILLER_158_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13568_ _13568_/A _13568_/B vssd1 vssd1 vccd1 vccd1 _13569_/C sky130_fd_sc_hd__xnor2_1
XFILLER_12_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15307_ _15307_/A _15307_/B _15307_/C vssd1 vssd1 vccd1 vccd1 _15307_/X sky130_fd_sc_hd__or3_1
XFILLER_9_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12519_ _12519_/A _12519_/B vssd1 vssd1 vccd1 vccd1 _12521_/B sky130_fd_sc_hd__xnor2_1
X_16287_ _16288_/B _16288_/A vssd1 vssd1 vccd1 vccd1 _16287_/Y sky130_fd_sc_hd__nand2b_1
X_13499_ _13500_/A _13500_/B _13500_/C vssd1 vssd1 vccd1 vccd1 _13501_/A sky130_fd_sc_hd__o21a_1
XFILLER_8_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15238_ _15238_/A _15450_/B _14924_/A vssd1 vssd1 vccd1 vccd1 _15241_/B sky130_fd_sc_hd__or3b_1
XFILLER_126_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15169_ _15169_/A _15169_/B vssd1 vssd1 vccd1 vccd1 _15171_/A sky130_fd_sc_hd__xnor2_1
Xfanout208 wire209/X vssd1 vssd1 vccd1 vccd1 _12046_/A sky130_fd_sc_hd__buf_4
Xfanout219 _17083_/A vssd1 vssd1 vccd1 vccd1 _16021_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_113_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09730_ _09731_/A _09729_/Y _09730_/C _10534_/D vssd1 vssd1 vccd1 vccd1 _09872_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_39_133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09661_ _09658_/A _09789_/A _09499_/Y _09500_/X vssd1 vssd1 vccd1 vccd1 _09662_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_39_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_924 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_795 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09592_ _09722_/A _09722_/B vssd1 vssd1 vccd1 vccd1 _09723_/A sky130_fd_sc_hd__and2_1
XFILLER_82_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09026_ _09026_/A _09269_/A vssd1 vssd1 vccd1 vccd1 _09033_/B sky130_fd_sc_hd__nor2_1
XFILLER_2_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_675 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout720 _17497_/Q vssd1 vssd1 vccd1 vccd1 _16480_/A sky130_fd_sc_hd__buf_4
XFILLER_104_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout731 _12054_/B vssd1 vssd1 vccd1 vccd1 _10299_/D sky130_fd_sc_hd__buf_2
Xfanout742 _14778_/B vssd1 vssd1 vccd1 vccd1 _13080_/D sky130_fd_sc_hd__buf_4
XFILLER_49_79 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09928_ _09929_/A _09927_/Y _10182_/C _14863_/A vssd1 vssd1 vccd1 vccd1 _10184_/A
+ sky130_fd_sc_hd__and4bb_1
Xfanout753 _17493_/Q vssd1 vssd1 vccd1 vccd1 _12334_/B sky130_fd_sc_hd__buf_4
Xfanout764 fanout772/X vssd1 vssd1 vccd1 vccd1 _12328_/B sky130_fd_sc_hd__buf_4
Xfanout775 _12166_/B vssd1 vssd1 vccd1 vccd1 _09030_/C sky130_fd_sc_hd__clkbuf_4
Xfanout786 _09229_/B vssd1 vssd1 vccd1 vccd1 _11961_/B sky130_fd_sc_hd__buf_4
XFILLER_74_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09859_ _15393_/A _16938_/A vssd1 vssd1 vccd1 vccd1 _15801_/A sky130_fd_sc_hd__nand2_4
Xfanout797 fanout805/X vssd1 vssd1 vccd1 vccd1 _12320_/D sky130_fd_sc_hd__buf_2
XTAP_3102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12870_ _12870_/A _12870_/B vssd1 vssd1 vccd1 vccd1 _12872_/A sky130_fd_sc_hd__nor2_1
XFILLER_73_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11821_ _11802_/Y _11804_/Y _11807_/Y _11809_/Y _17365_/A _12848_/S vssd1 vssd1 vccd1
+ vccd1 _11821_/X sky130_fd_sc_hd__mux4_1
XTAP_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_1003 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14540_ _14763_/S _14538_/X _14585_/B _14483_/Y vssd1 vssd1 vccd1 vccd1 _17599_/D
+ sky130_fd_sc_hd__a31o_1
XTAP_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11752_ _11223_/A _11223_/B _11224_/X vssd1 vssd1 vccd1 vccd1 _11753_/C sky130_fd_sc_hd__a21o_1
XTAP_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_854 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10703_ _11005_/A _10703_/B vssd1 vssd1 vccd1 vccd1 _11030_/A sky130_fd_sc_hd__nand2_1
XFILLER_41_353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14471_ _14471_/A _14471_/B vssd1 vssd1 vccd1 vccd1 _14472_/B sky130_fd_sc_hd__and2_1
XTAP_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11683_ _15106_/A _11683_/B vssd1 vssd1 vccd1 vccd1 _15235_/C sky130_fd_sc_hd__or2_1
XFILLER_14_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16210_ _16300_/A _16210_/B vssd1 vssd1 vccd1 vccd1 _16210_/Y sky130_fd_sc_hd__nor2_1
X_13422_ _13545_/A _13423_/B _13423_/C vssd1 vssd1 vccd1 vccd1 _13422_/X sky130_fd_sc_hd__and3_1
X_10634_ _10550_/A _10550_/B _10550_/C vssd1 vssd1 vccd1 vccd1 _10634_/Y sky130_fd_sc_hd__a21oi_1
X_17190_ input9/X input8/X input10/X input16/X vssd1 vssd1 vccd1 vccd1 _17191_/D sky130_fd_sc_hd__or4_1
XFILLER_167_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16141_ _16142_/A _16142_/B vssd1 vssd1 vccd1 vccd1 _16241_/B sky130_fd_sc_hd__nor2_1
X_13353_ _13353_/A _13353_/B vssd1 vssd1 vccd1 vccd1 _13355_/A sky130_fd_sc_hd__nor2_1
X_10565_ _10566_/A _10566_/B _10566_/C vssd1 vssd1 vccd1 vccd1 _10567_/A sky130_fd_sc_hd__a21oi_2
XFILLER_127_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12304_ _12305_/A _12305_/B _12305_/C vssd1 vssd1 vccd1 vccd1 _12306_/A sky130_fd_sc_hd__a21oi_1
X_16072_ _16072_/A _16072_/B _16072_/C vssd1 vssd1 vccd1 vccd1 _16073_/B sky130_fd_sc_hd__nor3_1
X_13284_ _13285_/B _13285_/A vssd1 vssd1 vccd1 vccd1 _13411_/A sky130_fd_sc_hd__nand2b_1
X_10496_ _10496_/A _10496_/B vssd1 vssd1 vccd1 vccd1 _10589_/A sky130_fd_sc_hd__xor2_1
XFILLER_136_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15023_ _15081_/A _16025_/A _15415_/A _15734_/A vssd1 vssd1 vccd1 vccd1 _15089_/S
+ sky130_fd_sc_hd__or4_2
X_12235_ _12714_/A _13080_/D _12235_/C vssd1 vssd1 vccd1 vccd1 _12236_/B sky130_fd_sc_hd__and3_1
XFILLER_146_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12166_ _17407_/A _12166_/B vssd1 vssd1 vccd1 vccd1 _12167_/B sky130_fd_sc_hd__nand2_1
XFILLER_69_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11117_ _11118_/A _11116_/Y _11117_/C _11117_/D vssd1 vssd1 vccd1 vccd1 _11246_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_7_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12097_ _12268_/A _12098_/B _12098_/C vssd1 vssd1 vccd1 vccd1 _12097_/X sky130_fd_sc_hd__a21o_1
X_16974_ _16974_/A _16974_/B vssd1 vssd1 vccd1 vccd1 _16974_/Y sky130_fd_sc_hd__nand2_1
X_11048_ _11048_/A _11048_/B vssd1 vssd1 vccd1 vccd1 _11051_/B sky130_fd_sc_hd__xor2_1
X_15925_ _15926_/A _15926_/B vssd1 vssd1 vccd1 vccd1 _15925_/Y sky130_fd_sc_hd__nor2_1
XFILLER_65_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput8 i_wb_addr[14] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__clkbuf_1
XFILLER_37_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15856_ _15666_/B _15853_/A _15756_/A _15756_/B vssd1 vssd1 vccd1 vccd1 _15858_/B
+ sky130_fd_sc_hd__a22oi_2
XFILLER_76_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14807_ _14785_/X _14806_/X _10716_/A vssd1 vssd1 vccd1 vccd1 _15623_/A sky130_fd_sc_hd__a21bo_1
XFILLER_24_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15787_ _15883_/B _15787_/B _15788_/B vssd1 vssd1 vccd1 vccd1 _15787_/X sky130_fd_sc_hd__or3b_1
X_12999_ _12999_/A _12999_/B vssd1 vssd1 vccd1 vccd1 _13001_/C sky130_fd_sc_hd__nand2_1
XFILLER_45_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17526_ fanout944/X _17526_/D vssd1 vssd1 vccd1 vccd1 _17526_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14738_ _14738_/A _14738_/B vssd1 vssd1 vccd1 vccd1 _17151_/A sky130_fd_sc_hd__nand2_2
XTAP_2990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17457_ fanout951/X _17457_/D vssd1 vssd1 vccd1 vccd1 _17457_/Q sky130_fd_sc_hd__dfxtp_2
X_14669_ _14638_/A _14669_/B vssd1 vssd1 vccd1 vccd1 _14669_/X sky130_fd_sc_hd__and2b_1
X_16408_ _16021_/A _16317_/B _15397_/A _16129_/B vssd1 vssd1 vccd1 vccd1 _16411_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_32_397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17388_ input39/X _17426_/A2 _17387_/X _17388_/C1 vssd1 vssd1 vccd1 vccd1 _17522_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_146_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16339_ _16339_/A _16339_/B _16339_/C vssd1 vssd1 vccd1 vccd1 _16340_/B sky130_fd_sc_hd__and3_1
XFILLER_145_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09713_ _10126_/B _10014_/D _10142_/B _10254_/A vssd1 vssd1 vccd1 vccd1 _09713_/X
+ sky130_fd_sc_hd__a22o_1
X_09644_ _09645_/B _09793_/A _09645_/A vssd1 vssd1 vccd1 vccd1 _09969_/A sky130_fd_sc_hd__o21a_1
XFILLER_56_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09575_ _09576_/A _09575_/B _09575_/C vssd1 vssd1 vccd1 vccd1 _09721_/A sky130_fd_sc_hd__nand3_1
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_990 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10350_ _17105_/A _10350_/B vssd1 vssd1 vccd1 vccd1 _11773_/A sky130_fd_sc_hd__nor2_1
XFILLER_136_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09009_ _09009_/A _09009_/B vssd1 vssd1 vccd1 vccd1 _09010_/B sky130_fd_sc_hd__nand2_1
XFILLER_151_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10281_ _10275_/X _10388_/A _10266_/X _10267_/Y vssd1 vssd1 vccd1 vccd1 _10283_/C
+ sky130_fd_sc_hd__o211ai_4
XFILLER_3_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12020_ _14911_/B _12020_/B vssd1 vssd1 vccd1 vccd1 _12020_/Y sky130_fd_sc_hd__nand2_1
XFILLER_104_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout550 _11930_/B vssd1 vssd1 vccd1 vccd1 _09325_/B sky130_fd_sc_hd__buf_2
Xfanout561 _17112_/A1 vssd1 vssd1 vccd1 vccd1 _14735_/A1 sky130_fd_sc_hd__buf_2
Xfanout572 _11470_/A vssd1 vssd1 vccd1 vccd1 _11553_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_59_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13971_ _13971_/A _13971_/B vssd1 vssd1 vccd1 vccd1 _13972_/B sky130_fd_sc_hd__or2_1
Xfanout583 _17164_/B vssd1 vssd1 vccd1 vccd1 _10180_/A sky130_fd_sc_hd__buf_2
XFILLER_65_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout594 _14954_/A vssd1 vssd1 vccd1 vccd1 _10182_/C sky130_fd_sc_hd__buf_2
X_15710_ _16015_/A _15811_/B _15710_/C vssd1 vssd1 vccd1 vccd1 _15710_/X sky130_fd_sc_hd__or3_1
X_12922_ _14050_/B _13067_/D _12923_/D _13434_/A vssd1 vssd1 vccd1 vccd1 _12924_/A
+ sky130_fd_sc_hd__a22oi_1
X_16690_ _16690_/A _16690_/B vssd1 vssd1 vccd1 vccd1 _16692_/B sky130_fd_sc_hd__xnor2_1
XFILLER_74_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15641_ _15913_/A _16419_/A vssd1 vssd1 vccd1 vccd1 _15732_/A sky130_fd_sc_hd__or2_1
X_12853_ _14636_/A _13626_/B vssd1 vssd1 vccd1 vccd1 _12853_/X sky130_fd_sc_hd__and2_1
XFILLER_74_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11804_ _11837_/A _11804_/B vssd1 vssd1 vccd1 vccd1 _11804_/Y sky130_fd_sc_hd__nand2_1
XTAP_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15572_ _15573_/B _15573_/A vssd1 vssd1 vccd1 vccd1 _15572_/Y sky130_fd_sc_hd__nand2b_1
XTAP_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12784_ _12781_/X _12938_/B _12631_/A _12631_/Y vssd1 vssd1 vccd1 vccd1 _12825_/B
+ sky130_fd_sc_hd__a211oi_1
XTAP_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17311_ input65/X _17321_/B _17321_/C vssd1 vssd1 vccd1 vccd1 _17311_/X sky130_fd_sc_hd__or3_1
XTAP_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14523_ _14577_/A _14523_/B vssd1 vssd1 vccd1 vccd1 _14524_/C sky130_fd_sc_hd__nand2_1
X_11735_ _11221_/A _11221_/B _11219_/Y vssd1 vssd1 vccd1 vccd1 _11735_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_30_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17242_ _17448_/Q _17293_/A2 _17240_/X _17241_/X _17284_/C1 vssd1 vssd1 vccd1 vccd1
+ _17448_/D sky130_fd_sc_hd__o221a_1
X_14454_ _14454_/A _14454_/B vssd1 vssd1 vccd1 vccd1 _14455_/B sky130_fd_sc_hd__or2_1
X_11666_ _11666_/A _11674_/A vssd1 vssd1 vccd1 vccd1 _11686_/B sky130_fd_sc_hd__nor2_1
XFILLER_174_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13405_ _13852_/A _13745_/B _13738_/B _13735_/D vssd1 vssd1 vccd1 vccd1 _13406_/B
+ sky130_fd_sc_hd__and4_1
X_10617_ _10617_/A _10617_/B vssd1 vssd1 vccd1 vccd1 _10624_/A sky130_fd_sc_hd__nor2_1
X_17173_ input27/X input26/X input24/X vssd1 vssd1 vccd1 vccd1 _17191_/A sky130_fd_sc_hd__or3b_1
XFILLER_127_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14385_ _16913_/C _14385_/B _14509_/A vssd1 vssd1 vccd1 vccd1 _14386_/B sky130_fd_sc_hd__and3_1
X_11597_ _11598_/A _11598_/B vssd1 vssd1 vccd1 vccd1 _11641_/A sky130_fd_sc_hd__and2_1
XFILLER_10_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16124_ _16103_/Y _16106_/Y _16123_/X _16494_/B1 _16114_/A vssd1 vssd1 vccd1 vccd1
+ _16125_/A sky130_fd_sc_hd__a32o_1
X_13336_ _13337_/A _13455_/A _13337_/C vssd1 vssd1 vccd1 vccd1 _13338_/A sky130_fd_sc_hd__o21a_1
XFILLER_41_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10548_ _10547_/A _10547_/B _10547_/C vssd1 vssd1 vccd1 vccd1 _10549_/B sky130_fd_sc_hd__o21ai_1
XFILLER_143_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16055_ _16055_/A _16827_/D vssd1 vssd1 vccd1 vccd1 _16454_/A sky130_fd_sc_hd__nor2_2
X_13267_ _13002_/A _13134_/Y _13137_/B vssd1 vssd1 vccd1 vccd1 _13267_/X sky130_fd_sc_hd__o21a_1
XFILLER_170_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10479_ _11027_/B _10479_/B vssd1 vssd1 vccd1 vccd1 _10480_/B sky130_fd_sc_hd__nand2_1
X_15006_ _11655_/A _14793_/Y _11675_/C vssd1 vssd1 vccd1 vccd1 _15006_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_130_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12218_ _12218_/A vssd1 vssd1 vccd1 vccd1 _12218_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_170_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13198_ _13199_/A _13199_/B _13199_/C vssd1 vssd1 vccd1 vccd1 _13369_/A sky130_fd_sc_hd__o21a_1
XFILLER_29_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1014 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12149_ _12149_/A _12149_/B vssd1 vssd1 vccd1 vccd1 _12150_/B sky130_fd_sc_hd__nor2_1
XFILLER_69_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16957_ _16958_/A _16958_/B vssd1 vssd1 vccd1 vccd1 _17037_/A sky130_fd_sc_hd__nand2b_1
XFILLER_96_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15908_ _15908_/A vssd1 vssd1 vccd1 vccd1 _17556_/D sky130_fd_sc_hd__clkinv_2
X_16888_ _16888_/A _16888_/B _16888_/C vssd1 vssd1 vccd1 vccd1 _16890_/A sky130_fd_sc_hd__nand3_1
XFILLER_65_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15839_ _15841_/A _15841_/B vssd1 vssd1 vccd1 vccd1 _15839_/Y sky130_fd_sc_hd__nor2_1
XFILLER_64_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09360_ _09360_/A _09502_/B _09502_/C vssd1 vssd1 vccd1 vccd1 _09497_/A sky130_fd_sc_hd__and3_1
XFILLER_80_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17509_ fanout944/X _17509_/D vssd1 vssd1 vccd1 vccd1 _17509_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09291_ _09292_/A _09291_/B _09291_/C vssd1 vssd1 vccd1 vccd1 _09437_/A sky130_fd_sc_hd__nand3_1
XFILLER_36_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_13 _14758_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_24 _17529_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_35 _17435_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_46 _09299_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_57 _13966_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_68 _15151_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_79 _16880_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_824 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09627_ _09627_/A _09773_/A vssd1 vssd1 vccd1 vccd1 _09628_/C sky130_fd_sc_hd__nor2_1
XFILLER_16_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09558_ _09558_/A _09558_/B vssd1 vssd1 vccd1 vccd1 _09689_/A sky130_fd_sc_hd__xnor2_1
XFILLER_71_768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09489_ _09498_/A _09489_/B vssd1 vssd1 vccd1 vccd1 _09508_/A sky130_fd_sc_hd__xnor2_1
X_11520_ _11521_/A _11519_/Y _11520_/C _11561_/C vssd1 vssd1 vccd1 vccd1 _11565_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_12_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_194 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11451_ _11451_/A _11451_/B _11495_/A vssd1 vssd1 vccd1 vccd1 _11456_/A sky130_fd_sc_hd__nor3b_1
XFILLER_109_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_531 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10402_ _10402_/A _10402_/B _10402_/C vssd1 vssd1 vccd1 vccd1 _10402_/Y sky130_fd_sc_hd__nand3_1
X_14170_ _14170_/A _14245_/A _14170_/C vssd1 vssd1 vccd1 vccd1 _14245_/B sky130_fd_sc_hd__nor3_1
X_11382_ _11376_/A _11376_/C _11376_/B vssd1 vssd1 vccd1 vccd1 _11383_/C sky130_fd_sc_hd__a21o_1
XFILLER_125_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13121_ _13121_/A _13121_/B _13121_/C vssd1 vssd1 vccd1 vccd1 _13123_/A sky130_fd_sc_hd__nor3_1
X_10333_ _10333_/A _10333_/B vssd1 vssd1 vccd1 vccd1 _10334_/B sky130_fd_sc_hd__xnor2_1
XFILLER_139_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13052_ _13052_/A _13314_/A vssd1 vssd1 vccd1 vccd1 _13055_/A sky130_fd_sc_hd__or2_1
XFILLER_152_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10264_ _10249_/Y _10262_/X _10134_/Y _10231_/X vssd1 vssd1 vccd1 vccd1 _10283_/A
+ sky130_fd_sc_hd__o211ai_1
XFILLER_105_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_792 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12003_ _12200_/A _12001_/Y _09250_/Y _09255_/B vssd1 vssd1 vccd1 vccd1 _12004_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_87_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10195_ _10321_/B _10446_/B vssd1 vssd1 vccd1 vccd1 _10322_/A sky130_fd_sc_hd__nand2_1
XFILLER_105_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_98 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16811_ _16811_/A _16811_/B vssd1 vssd1 vccd1 vccd1 _16818_/A sky130_fd_sc_hd__xnor2_1
XFILLER_93_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout380 _17534_/Q vssd1 vssd1 vccd1 vccd1 fanout380/X sky130_fd_sc_hd__clkbuf_4
XFILLER_93_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout391 _12795_/A vssd1 vssd1 vccd1 vccd1 _17407_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_93_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16742_ _15658_/Y _16662_/C _16662_/D _16883_/A vssd1 vssd1 vccd1 vccd1 _16744_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_143_82 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13954_ _13954_/A _13954_/B _13954_/C vssd1 vssd1 vccd1 vccd1 _13955_/B sky130_fd_sc_hd__or3_1
XFILLER_93_359 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12905_ _13182_/A _13051_/B _13051_/D _13037_/B vssd1 vssd1 vccd1 vccd1 _12905_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_46_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16673_ _16673_/A _16673_/B vssd1 vssd1 vccd1 vccd1 _16674_/B sky130_fd_sc_hd__or2_1
X_13885_ _13885_/A _13885_/B vssd1 vssd1 vccd1 vccd1 _13888_/A sky130_fd_sc_hd__xor2_1
XFILLER_59_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12836_ _12651_/A _12655_/A _12833_/Y _12835_/X vssd1 vssd1 vccd1 vccd1 _13001_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_61_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15624_ _15624_/A _15624_/B vssd1 vssd1 vccd1 vccd1 _15624_/Y sky130_fd_sc_hd__nor2_1
XFILLER_34_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15555_ _15645_/B _15555_/B vssd1 vssd1 vccd1 vccd1 _15557_/A sky130_fd_sc_hd__xor2_1
XFILLER_15_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12767_ _12612_/A _12612_/Y _12765_/Y _12920_/B vssd1 vssd1 vccd1 vccd1 _12938_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_14_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14506_ _14565_/A _14506_/B vssd1 vssd1 vccd1 vccd1 _14508_/B sky130_fd_sc_hd__nor2_1
X_11718_ _11717_/A _16387_/C _11717_/X _16206_/A _11231_/X vssd1 vssd1 vccd1 vccd1
+ _16568_/A sky130_fd_sc_hd__a221o_2
X_15486_ _15486_/A _15486_/B vssd1 vssd1 vccd1 vccd1 _15489_/A sky130_fd_sc_hd__xnor2_1
XFILLER_14_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12698_ _13003_/A _12698_/B vssd1 vssd1 vccd1 vccd1 _12698_/Y sky130_fd_sc_hd__nor2_1
XFILLER_174_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17225_ _17584_/Q _17225_/A2 _17225_/B1 vssd1 vssd1 vccd1 vccd1 _17225_/X sky130_fd_sc_hd__a21o_1
X_14437_ _14554_/A _14641_/C _14437_/C vssd1 vssd1 vccd1 vccd1 _14438_/B sky130_fd_sc_hd__and3_1
X_11649_ _11649_/A _11649_/B vssd1 vssd1 vccd1 vccd1 _11657_/A sky130_fd_sc_hd__xor2_1
Xinput11 i_wb_addr[17] vssd1 vssd1 vccd1 vccd1 input11/X sky130_fd_sc_hd__clkbuf_1
XFILLER_128_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput22 i_wb_addr[27] vssd1 vssd1 vccd1 vccd1 input22/X sky130_fd_sc_hd__clkbuf_1
XFILLER_128_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput33 i_wb_addr[8] vssd1 vssd1 vccd1 vccd1 input33/X sky130_fd_sc_hd__clkbuf_1
XFILLER_174_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput44 i_wb_data[17] vssd1 vssd1 vccd1 vccd1 input44/X sky130_fd_sc_hd__clkbuf_1
X_17156_ _17156_/A _17156_/B _17154_/X vssd1 vssd1 vccd1 vccd1 _17156_/X sky130_fd_sc_hd__or3b_1
XFILLER_7_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput55 i_wb_data[27] vssd1 vssd1 vccd1 vccd1 input55/X sky130_fd_sc_hd__clkbuf_1
X_14368_ _14554_/A _14641_/D _14368_/C vssd1 vssd1 vccd1 vccd1 _14370_/A sky130_fd_sc_hd__and3_1
Xinput66 i_wb_data[8] vssd1 vssd1 vccd1 vccd1 input66/X sky130_fd_sc_hd__clkbuf_1
XFILLER_128_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16107_ _16108_/C _16644_/B _16114_/A vssd1 vssd1 vccd1 vccd1 _16107_/Y sky130_fd_sc_hd__a21boi_2
X_13319_ _13316_/Y _13431_/B _13189_/A _13189_/Y vssd1 vssd1 vccd1 vccd1 _13329_/B
+ sky130_fd_sc_hd__o211ai_1
X_17087_ _17088_/A _17088_/B _17088_/C vssd1 vssd1 vccd1 vccd1 _17089_/A sky130_fd_sc_hd__o21a_1
XFILLER_115_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14299_ _14599_/B _14301_/C _14485_/D _14680_/A vssd1 vssd1 vccd1 vccd1 _14302_/A
+ sky130_fd_sc_hd__a22oi_1
X_16038_ _15647_/A _16591_/B _15916_/X _15918_/X vssd1 vssd1 vccd1 vccd1 _16044_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_131_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08860_ _17381_/A _08860_/B vssd1 vssd1 vccd1 vccd1 _08861_/B sky130_fd_sc_hd__nand2_1
XFILLER_69_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08791_ _08791_/A _08791_/B _09319_/D _09058_/C vssd1 vssd1 vccd1 vccd1 _11878_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_85_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_998 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09412_ _09412_/A _10933_/C vssd1 vssd1 vccd1 vccd1 _16983_/A sky130_fd_sc_hd__nand2_8
XFILLER_25_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09343_ _09344_/A _09344_/B _09344_/C vssd1 vssd1 vccd1 vccd1 _09343_/X sky130_fd_sc_hd__o21a_2
XFILLER_52_278 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09274_ _16982_/A _09274_/B vssd1 vssd1 vccd1 vccd1 _09404_/A sky130_fd_sc_hd__xnor2_1
XFILLER_165_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_364 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08989_ _08989_/A _08989_/B vssd1 vssd1 vccd1 vccd1 _08991_/A sky130_fd_sc_hd__nor2_1
XFILLER_57_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_186 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10951_ _10951_/A _11065_/A vssd1 vssd1 vccd1 vccd1 _10953_/B sky130_fd_sc_hd__and2_1
XFILLER_90_329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13670_ _13671_/A _13671_/B _13671_/C vssd1 vssd1 vccd1 vccd1 _13670_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_43_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10882_ _10883_/B _10883_/C _10883_/A vssd1 vssd1 vccd1 vccd1 _10893_/A sky130_fd_sc_hd__a21o_1
XFILLER_16_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12621_ _12621_/A _12621_/B vssd1 vssd1 vccd1 vccd1 _12623_/B sky130_fd_sc_hd__xnor2_1
XFILLER_19_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15340_ _16315_/C _15493_/A _15755_/B _15081_/A vssd1 vssd1 vccd1 vccd1 _15340_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_12_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12552_ _13516_/S _12552_/B vssd1 vssd1 vccd1 vccd1 _12553_/B sky130_fd_sc_hd__or2_1
XFILLER_12_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11503_ _11502_/B _11502_/C _11502_/A vssd1 vssd1 vccd1 vccd1 _11543_/B sky130_fd_sc_hd__o21a_1
XFILLER_106_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15271_ _15207_/X _15270_/X _11437_/D vssd1 vssd1 vccd1 vccd1 _16505_/A sky130_fd_sc_hd__a21boi_4
XFILLER_156_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12483_ _12479_/Y _12480_/X _12312_/A _12314_/A vssd1 vssd1 vccd1 vccd1 _12522_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_7_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_840 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17010_ _17037_/B _17010_/B vssd1 vssd1 vccd1 vccd1 _17014_/B sky130_fd_sc_hd__xor2_1
X_14222_ _14222_/A _14222_/B vssd1 vssd1 vccd1 vccd1 _14262_/A sky130_fd_sc_hd__nand2_1
X_11434_ _11433_/B _11433_/C _11433_/A vssd1 vssd1 vccd1 vccd1 _11435_/C sky130_fd_sc_hd__a21bo_1
XFILLER_144_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14153_ _14153_/A _14153_/B _14426_/D _14360_/D vssd1 vssd1 vccd1 vccd1 _14154_/B
+ sky130_fd_sc_hd__and4_1
X_11365_ _11447_/A _11447_/B vssd1 vssd1 vccd1 vccd1 _11448_/A sky130_fd_sc_hd__or2_1
XFILLER_138_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13104_ _12964_/A _12966_/B _12964_/B vssd1 vssd1 vccd1 vccd1 _13106_/B sky130_fd_sc_hd__o21ba_1
XFILLER_4_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10316_ _10303_/Y _10315_/X _10330_/A _10287_/Y vssd1 vssd1 vccd1 vccd1 _10330_/B
+ sky130_fd_sc_hd__o211ai_4
X_14084_ _14084_/A _14084_/B vssd1 vssd1 vccd1 vccd1 _14087_/B sky130_fd_sc_hd__xnor2_1
XFILLER_98_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11296_ _11345_/A _11345_/B vssd1 vssd1 vccd1 vccd1 _11296_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_106_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13035_ _13035_/A _13414_/B _13035_/C _13908_/B vssd1 vssd1 vccd1 vccd1 _13036_/B
+ sky130_fd_sc_hd__and4_1
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10247_ _10358_/A _10358_/B vssd1 vssd1 vccd1 vccd1 _10261_/C sky130_fd_sc_hd__nand2_1
XFILLER_67_805 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10178_ _10182_/C _10180_/B _09929_/A _09927_/Y vssd1 vssd1 vccd1 vccd1 _10184_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_120_272 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14986_ _15100_/A _14986_/B vssd1 vssd1 vccd1 vccd1 _14986_/Y sky130_fd_sc_hd__nand2_1
XFILLER_81_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16725_ _16791_/A _16723_/Y _16643_/A _16648_/C vssd1 vssd1 vccd1 vccd1 _16725_/X
+ sky130_fd_sc_hd__a211o_1
X_13937_ _13727_/A _13825_/Y _13826_/Y _13936_/Y vssd1 vssd1 vccd1 vccd1 _13937_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_62_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13868_ _14215_/A _14050_/D vssd1 vssd1 vccd1 vccd1 _13869_/B sky130_fd_sc_hd__nand2_1
X_16656_ _17164_/C _15246_/X _16653_/X _16655_/X vssd1 vssd1 vccd1 vccd1 _16656_/X
+ sky130_fd_sc_hd__o211a_1
X_12819_ _12820_/A _12820_/B _12820_/C vssd1 vssd1 vccd1 vccd1 _12819_/X sky130_fd_sc_hd__a21o_1
XFILLER_62_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15607_ _15607_/A _15607_/B vssd1 vssd1 vccd1 vccd1 _15609_/C sky130_fd_sc_hd__xor2_1
X_16587_ _16566_/A _16566_/B _16560_/A vssd1 vssd1 vccd1 vccd1 _16639_/A sky130_fd_sc_hd__o21ai_1
XFILLER_16_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13799_ _13800_/A _13800_/B _13800_/C vssd1 vssd1 vccd1 vccd1 _13801_/A sky130_fd_sc_hd__a21oi_1
XFILLER_97_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15538_ _15538_/A _15538_/B vssd1 vssd1 vccd1 vccd1 _15538_/X sky130_fd_sc_hd__or2_1
XFILLER_147_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15469_ _15463_/A _16494_/B1 _15468_/X vssd1 vssd1 vccd1 vccd1 _17551_/D sky130_fd_sc_hd__a21oi_2
XFILLER_147_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17208_ _17546_/Q _17274_/B vssd1 vssd1 vccd1 vccd1 _17208_/X sky130_fd_sc_hd__and2_1
XFILLER_163_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17139_ _17139_/A _17139_/B vssd1 vssd1 vccd1 vccd1 _17140_/C sky130_fd_sc_hd__nor2_1
XFILLER_171_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_556 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09961_ _09960_/A _09960_/Y _09813_/X _09829_/Y vssd1 vssd1 vccd1 vccd1 _09964_/A
+ sky130_fd_sc_hd__a211oi_2
XFILLER_116_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08912_ _08912_/A _08912_/B vssd1 vssd1 vccd1 vccd1 _08918_/A sky130_fd_sc_hd__nor2_1
XFILLER_131_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09892_ _09892_/A _09892_/B _10421_/D _10534_/D vssd1 vssd1 vccd1 vccd1 _09895_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_134_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08843_ _08843_/A _08912_/A vssd1 vssd1 vccd1 vccd1 _08845_/B sky130_fd_sc_hd__nor2_1
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08774_ _08780_/B _08780_/A vssd1 vssd1 vccd1 vccd1 _08783_/B sky130_fd_sc_hd__and2b_1
XFILLER_57_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_562 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09326_ _09325_/B _09926_/B _10180_/B _12471_/A vssd1 vssd1 vccd1 vccd1 _09326_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_166_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09257_ _09257_/A _09257_/B vssd1 vssd1 vccd1 vccd1 _09391_/A sky130_fd_sc_hd__xnor2_1
XFILLER_126_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09188_ _09189_/A _09221_/A _09189_/C vssd1 vssd1 vccd1 vccd1 _09190_/A sky130_fd_sc_hd__o21a_1
XFILLER_5_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11150_ _11145_/A _11145_/B _11145_/C vssd1 vssd1 vccd1 vccd1 _11151_/C sky130_fd_sc_hd__a21oi_1
XFILLER_135_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_1047 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10101_ _10101_/A _10101_/B vssd1 vssd1 vccd1 vccd1 _10223_/A sky130_fd_sc_hd__nor2_1
XFILLER_89_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11081_ _11080_/B _11145_/A _11064_/X _11071_/Y vssd1 vssd1 vccd1 vccd1 _11084_/A
+ sky130_fd_sc_hd__a211oi_2
XFILLER_88_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10032_ _09910_/B _10030_/Y _10027_/C _10010_/A vssd1 vssd1 vccd1 vccd1 _10033_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_48_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_495 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_272 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14840_ _17371_/A _14840_/B vssd1 vssd1 vccd1 vccd1 _14840_/Y sky130_fd_sc_hd__nor2_1
XFILLER_75_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14771_ _17409_/A _14863_/A vssd1 vssd1 vccd1 vccd1 _16796_/B sky130_fd_sc_hd__or2_1
X_11983_ _11984_/A _11984_/B vssd1 vssd1 vccd1 vccd1 _12183_/B sky130_fd_sc_hd__and2b_1
XFILLER_44_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16510_ _16616_/A _16510_/B vssd1 vssd1 vccd1 vccd1 _16524_/A sky130_fd_sc_hd__or2_1
XFILLER_1_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13722_ _13723_/A _13723_/B vssd1 vssd1 vccd1 vccd1 _13824_/B sky130_fd_sc_hd__or2_1
X_10934_ _11122_/B _10933_/C _10933_/D _10933_/A vssd1 vssd1 vccd1 vccd1 _10935_/B
+ sky130_fd_sc_hd__a22oi_1
X_17490_ fanout942/X _17490_/D vssd1 vssd1 vccd1 vccd1 _17490_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16441_ _16442_/A _16442_/B vssd1 vssd1 vccd1 vccd1 _16550_/A sky130_fd_sc_hd__nand2_1
X_13653_ _13543_/A _13543_/B _13537_/Y vssd1 vssd1 vccd1 vccd1 _13654_/B sky130_fd_sc_hd__o21bai_1
X_10865_ _10865_/A _10865_/B vssd1 vssd1 vccd1 vccd1 _10883_/A sky130_fd_sc_hd__xnor2_1
XFILLER_140_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12604_ _12605_/A _12605_/B vssd1 vssd1 vccd1 vccd1 _12764_/B sky130_fd_sc_hd__nand2b_1
XPHY_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16372_ _16372_/A _16372_/B vssd1 vssd1 vccd1 vccd1 _16375_/A sky130_fd_sc_hd__xnor2_2
XPHY_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13584_ _13584_/A _13584_/B vssd1 vssd1 vccd1 vccd1 _13586_/C sky130_fd_sc_hd__xnor2_1
X_10796_ _10901_/B _10796_/B _10860_/B vssd1 vssd1 vccd1 vccd1 _11082_/A sky130_fd_sc_hd__or3_1
XPHY_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_412 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15323_ _15314_/A _16494_/B1 _15322_/X vssd1 vssd1 vccd1 vccd1 _17549_/D sky130_fd_sc_hd__a21oi_2
XFILLER_157_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12535_ _12331_/Y _12333_/B _12336_/A vssd1 vssd1 vccd1 vccd1 _12536_/B sky130_fd_sc_hd__a21oi_2
XFILLER_158_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_927 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15254_ _14992_/Y _14998_/Y _15254_/S vssd1 vssd1 vccd1 vccd1 _15254_/X sky130_fd_sc_hd__mux2_1
X_12466_ _12467_/A _12467_/B vssd1 vssd1 vccd1 vccd1 _12662_/B sky130_fd_sc_hd__nor2_1
XFILLER_144_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14205_ _14279_/A _14205_/B vssd1 vssd1 vccd1 vccd1 _14207_/B sky130_fd_sc_hd__and2b_1
X_11417_ _11418_/A _11418_/B vssd1 vssd1 vccd1 vccd1 _11713_/A sky130_fd_sc_hd__and2b_1
X_15185_ _15175_/B _14848_/C _16015_/A vssd1 vssd1 vccd1 vccd1 _15185_/Y sky130_fd_sc_hd__a21oi_1
X_12397_ _15095_/B _12397_/B vssd1 vssd1 vccd1 vccd1 _13837_/C sky130_fd_sc_hd__or2_1
XFILLER_153_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14136_ _14218_/B _14136_/B vssd1 vssd1 vccd1 vccd1 _14138_/B sky130_fd_sc_hd__or2_1
X_11348_ _11348_/A _11348_/B vssd1 vssd1 vccd1 vccd1 _11349_/C sky130_fd_sc_hd__and2_1
XFILLER_99_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14067_ _14068_/A _14068_/B vssd1 vssd1 vccd1 vccd1 _14162_/A sky130_fd_sc_hd__and2b_1
XFILLER_98_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11279_ _11518_/B _14893_/B _15208_/A _11561_/A vssd1 vssd1 vccd1 vccd1 _11280_/B
+ sky130_fd_sc_hd__a22oi_1
X_13018_ _13735_/A _13632_/B _14063_/C _14213_/D vssd1 vssd1 vccd1 vccd1 _13019_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_79_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14969_ _14899_/X _14968_/X _11675_/B vssd1 vssd1 vccd1 vccd1 _14969_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_63_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16708_ _16709_/B _16709_/A vssd1 vssd1 vccd1 vccd1 _16784_/B sky130_fd_sc_hd__nand2b_1
XFILLER_62_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16639_ _16639_/A _16854_/C vssd1 vssd1 vccd1 vccd1 _16639_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_62_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09111_ _09153_/B _09111_/B vssd1 vssd1 vccd1 vccd1 _09314_/B sky130_fd_sc_hd__or2_1
XFILLER_31_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09042_ _17387_/A _09042_/B vssd1 vssd1 vccd1 vccd1 _09279_/A sky130_fd_sc_hd__nand2_1
XFILLER_108_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_684 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09944_ _09945_/A _09943_/Y _10321_/A _10446_/B vssd1 vssd1 vccd1 vccd1 _10064_/A
+ sky130_fd_sc_hd__and4bb_1
Xfanout902 fanout904/X vssd1 vssd1 vccd1 vccd1 _11027_/C sky130_fd_sc_hd__buf_4
Xfanout913 _17273_/B1 vssd1 vssd1 vccd1 vccd1 _17291_/B1 sky130_fd_sc_hd__buf_2
XFILLER_104_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout924 _17428_/B vssd1 vssd1 vccd1 vccd1 _17364_/C1 sky130_fd_sc_hd__clkbuf_4
XFILLER_86_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout935 fanout936/X vssd1 vssd1 vccd1 vccd1 fanout935/X sky130_fd_sc_hd__clkbuf_2
XFILLER_86_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout946 fanout947/X vssd1 vssd1 vccd1 vccd1 fanout946/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_86_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout957 input2/X vssd1 vssd1 vccd1 vccd1 fanout957/X sky130_fd_sc_hd__buf_6
X_09875_ _09876_/A _09874_/Y _10271_/A _10036_/D vssd1 vssd1 vccd1 vccd1 _10018_/A
+ sky130_fd_sc_hd__and4bb_1
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08826_ _08826_/A _08826_/B vssd1 vssd1 vccd1 vccd1 _08893_/B sky130_fd_sc_hd__nor2_1
XFILLER_86_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08757_ _08757_/A _08757_/B vssd1 vssd1 vccd1 vccd1 _08766_/A sky130_fd_sc_hd__xor2_4
XTAP_2605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_649 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10650_ _10735_/A _10735_/B vssd1 vssd1 vccd1 vccd1 _10653_/C sky130_fd_sc_hd__nand2_1
XFILLER_13_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09309_ _09303_/X _09439_/A _09316_/A _09296_/Y vssd1 vssd1 vccd1 vccd1 _09316_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_10_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10581_ _10581_/A _10581_/B _10581_/C vssd1 vssd1 vccd1 vccd1 _11771_/B sky130_fd_sc_hd__or3_1
XFILLER_16_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12320_ _17413_/A _12787_/B _12487_/D _12320_/D vssd1 vssd1 vccd1 vccd1 _12492_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_139_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12251_ _12252_/A _12252_/B _12252_/C vssd1 vssd1 vccd1 vccd1 _12437_/A sky130_fd_sc_hd__o21ai_1
XFILLER_79_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11202_ _11202_/A _11202_/B vssd1 vssd1 vccd1 vccd1 _11204_/B sky130_fd_sc_hd__and2_1
XFILLER_135_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12182_ _12182_/A _12182_/B vssd1 vssd1 vccd1 vccd1 _12351_/A sky130_fd_sc_hd__xor2_1
XFILLER_134_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11133_ _11132_/B _11132_/C _11281_/B _11561_/A vssd1 vssd1 vccd1 vccd1 _11134_/B
+ sky130_fd_sc_hd__a22oi_1
XFILLER_122_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16990_ _16990_/A _16990_/B vssd1 vssd1 vccd1 vccd1 _16991_/D sky130_fd_sc_hd__nand2_2
XFILLER_135_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_676 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11064_ _11065_/A _11065_/B _11065_/C _11065_/D vssd1 vssd1 vccd1 vccd1 _11064_/X
+ sky130_fd_sc_hd__and4_1
X_15941_ _15941_/A _15941_/B vssd1 vssd1 vccd1 vccd1 _15944_/A sky130_fd_sc_hd__xnor2_1
XFILLER_122_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_94 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_635 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10015_ _14784_/A _10146_/B _10014_/D _10142_/A vssd1 vssd1 vccd1 vccd1 _10015_/Y
+ sky130_fd_sc_hd__a22oi_1
X_15872_ _16281_/A _16259_/B _15872_/C vssd1 vssd1 vccd1 vccd1 _15989_/B sky130_fd_sc_hd__and3_1
XFILLER_92_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17611_ fanout954/X _17611_/D vssd1 vssd1 vccd1 vccd1 _17611_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14823_ _16918_/B _16918_/C _14080_/C vssd1 vssd1 vccd1 vccd1 _16971_/A sky130_fd_sc_hd__a21oi_1
XFILLER_48_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17542_ fanout941/X _17542_/D vssd1 vssd1 vccd1 vccd1 _17542_/Q sky130_fd_sc_hd__dfxtp_1
X_11966_ _11965_/B _11966_/B vssd1 vssd1 vccd1 vccd1 _11967_/B sky130_fd_sc_hd__nand2b_1
X_14754_ _14755_/A _14755_/B vssd1 vssd1 vccd1 vccd1 _14754_/Y sky130_fd_sc_hd__nand2_1
XFILLER_44_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10917_ _10918_/B _10918_/A vssd1 vssd1 vccd1 vccd1 _11049_/A sky130_fd_sc_hd__and2b_1
XFILLER_32_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13705_ _13705_/A _13705_/B vssd1 vssd1 vccd1 vccd1 _13707_/B sky130_fd_sc_hd__xnor2_1
XFILLER_44_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17473_ fanout955/X _17546_/Q vssd1 vssd1 vccd1 vccd1 _17473_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14685_ _14710_/C _14710_/B _14684_/A vssd1 vssd1 vccd1 vccd1 _14686_/B sky130_fd_sc_hd__a21oi_1
X_11897_ _17375_/A _12447_/B _11894_/Y _12138_/A vssd1 vssd1 vccd1 vccd1 _11898_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_16424_ _16425_/A _16425_/B _16423_/A _16509_/B vssd1 vssd1 vccd1 vccd1 _16527_/A
+ sky130_fd_sc_hd__o211a_1
X_13636_ _13635_/A _13741_/A _13635_/C vssd1 vssd1 vccd1 vccd1 _13638_/B sky130_fd_sc_hd__o21ai_1
XFILLER_60_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10848_ _15116_/A _15206_/A _10836_/A _10834_/Y vssd1 vssd1 vccd1 vccd1 _10850_/C
+ sky130_fd_sc_hd__o22a_1
XFILLER_20_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16355_ _16355_/A _16355_/B vssd1 vssd1 vccd1 vccd1 _16356_/B sky130_fd_sc_hd__nand2_1
XFILLER_158_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13567_ _13897_/A _13691_/C _13568_/A vssd1 vssd1 vccd1 vccd1 _13695_/B sky130_fd_sc_hd__and3_1
X_10779_ _10779_/A _10779_/B vssd1 vssd1 vccd1 vccd1 _11749_/B sky130_fd_sc_hd__xnor2_1
XFILLER_118_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_702 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12518_ _12518_/A _12518_/B vssd1 vssd1 vccd1 vccd1 _12519_/B sky130_fd_sc_hd__xnor2_1
X_15306_ _15241_/B _15241_/C _15241_/A vssd1 vssd1 vccd1 vccd1 _15307_/C sky130_fd_sc_hd__a21boi_1
X_16286_ _16189_/B _16191_/B _16187_/Y vssd1 vssd1 vccd1 vccd1 _16288_/B sky130_fd_sc_hd__o21a_1
X_13498_ _13498_/A _13498_/B vssd1 vssd1 vccd1 vccd1 _13500_/C sky130_fd_sc_hd__xnor2_1
XFILLER_60_90 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12449_ _12276_/A _12278_/B _12276_/B vssd1 vssd1 vccd1 vccd1 _12451_/B sky130_fd_sc_hd__o21ba_1
X_15237_ _15237_/A1 _15373_/B _15238_/A vssd1 vssd1 vccd1 vccd1 _15241_/A sky130_fd_sc_hd__a21bo_1
XFILLER_172_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15168_ _15169_/A _15169_/B vssd1 vssd1 vccd1 vccd1 _15168_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_119_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1023 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_846 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14119_ _14119_/A _14119_/B _14117_/X vssd1 vssd1 vccd1 vccd1 _14120_/B sky130_fd_sc_hd__or3b_1
XFILLER_4_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15099_ _14863_/A _14864_/A _11808_/B _12025_/B _09925_/A _15095_/B vssd1 vssd1 vccd1
+ vccd1 _15100_/B sky130_fd_sc_hd__mux4_1
XFILLER_86_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09660_ _09499_/Y _09500_/X _09658_/A _09789_/A vssd1 vssd1 vccd1 vccd1 _09662_/A
+ sky130_fd_sc_hd__a211oi_1
XFILLER_95_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09591_ _09591_/A _09591_/B vssd1 vssd1 vccd1 vccd1 _09722_/B sky130_fd_sc_hd__nor2_1
XFILLER_83_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09025_ _09026_/A _09024_/Y _12070_/A _12338_/C vssd1 vssd1 vccd1 vccd1 _09269_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_156_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_8 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_868 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout710 _13968_/B vssd1 vssd1 vccd1 vccd1 _13450_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_49_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout721 _12077_/C vssd1 vssd1 vccd1 vccd1 _09058_/C sky130_fd_sc_hd__buf_2
XFILLER_132_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout732 _17496_/Q vssd1 vssd1 vccd1 vccd1 _12054_/B sky130_fd_sc_hd__buf_4
XFILLER_77_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09927_ _15254_/S _10309_/B _09652_/C vssd1 vssd1 vccd1 vccd1 _09927_/Y sky130_fd_sc_hd__a21oi_1
Xfanout743 _14778_/B vssd1 vssd1 vccd1 vccd1 _13764_/D sky130_fd_sc_hd__buf_2
XFILLER_58_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout754 _16760_/A vssd1 vssd1 vccd1 vccd1 _16935_/A sky130_fd_sc_hd__buf_2
XFILLER_58_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout765 _15204_/B vssd1 vssd1 vccd1 vccd1 _16880_/A sky130_fd_sc_hd__buf_2
Xfanout776 _17491_/Q vssd1 vssd1 vccd1 vccd1 _12166_/B sky130_fd_sc_hd__buf_4
XFILLER_58_443 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09858_ _11005_/A _10933_/C vssd1 vssd1 vccd1 vccd1 _16809_/B sky130_fd_sc_hd__and2_4
Xfanout787 fanout795/X vssd1 vssd1 vccd1 vccd1 _09229_/B sky130_fd_sc_hd__clkbuf_4
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout798 fanout805/X vssd1 vssd1 vccd1 vccd1 _09272_/D sky130_fd_sc_hd__buf_4
XTAP_3103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08809_ _08815_/B _08815_/A vssd1 vssd1 vccd1 vccd1 _08831_/B sky130_fd_sc_hd__and2b_1
XTAP_3136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09789_ _09789_/A _09789_/B vssd1 vssd1 vccd1 vccd1 _09790_/B sky130_fd_sc_hd__nor2_1
XTAP_3147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11820_ _11820_/A vssd1 vssd1 vccd1 vccd1 _11820_/Y sky130_fd_sc_hd__clkinv_2
XTAP_3169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_863 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11751_ _11739_/B _11739_/C _11739_/A vssd1 vssd1 vccd1 vccd1 _11753_/B sky130_fd_sc_hd__o21ai_1
XFILLER_26_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10702_ _10954_/A _10904_/A _11005_/B _10805_/D vssd1 vssd1 vccd1 vccd1 _10705_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_42_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14470_ _14471_/A _14471_/B vssd1 vssd1 vccd1 vccd1 _14531_/B sky130_fd_sc_hd__nor2_1
XTAP_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11682_ _11681_/A _11678_/A _11681_/B _11662_/B _11680_/Y vssd1 vssd1 vccd1 vccd1
+ _11683_/B sky130_fd_sc_hd__a311o_1
XFILLER_14_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13421_ _13545_/A _13423_/B _13423_/C vssd1 vssd1 vccd1 vccd1 _13421_/Y sky130_fd_sc_hd__a21oi_1
X_10633_ _10632_/A _10632_/Y _10519_/Y _10588_/X vssd1 vssd1 vccd1 vccd1 _10667_/A
+ sky130_fd_sc_hd__a211oi_4
XFILLER_14_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16140_ _16140_/A _16140_/B vssd1 vssd1 vccd1 vccd1 _16142_/B sky130_fd_sc_hd__xor2_1
XFILLER_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13352_ _14153_/A _13352_/B _13764_/D _13664_/D vssd1 vssd1 vccd1 vccd1 _13353_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_6_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10564_ _10564_/A _10564_/B vssd1 vssd1 vccd1 vccd1 _10566_/C sky130_fd_sc_hd__nand2_1
X_12303_ _12303_/A _12303_/B vssd1 vssd1 vccd1 vccd1 _12305_/C sky130_fd_sc_hd__xnor2_1
X_16071_ _16072_/A _16072_/B _16072_/C vssd1 vssd1 vccd1 vccd1 _16188_/A sky130_fd_sc_hd__o21a_1
X_13283_ _13149_/A _13151_/B _13149_/B vssd1 vssd1 vccd1 vccd1 _13285_/B sky130_fd_sc_hd__o21ba_1
X_10495_ _10496_/B _10496_/A vssd1 vssd1 vccd1 vccd1 _10503_/B sky130_fd_sc_hd__nand2b_1
XFILLER_136_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15022_ _16127_/A _15278_/A _16226_/B _15846_/A vssd1 vssd1 vccd1 vccd1 _15030_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_154_278 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12234_ _12714_/A _13080_/D _12235_/C vssd1 vssd1 vccd1 vccd1 _12236_/A sky130_fd_sc_hd__a21oi_1
XFILLER_108_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_930 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12165_ _12165_/A _12165_/B vssd1 vssd1 vccd1 vccd1 _12167_/A sky130_fd_sc_hd__nor2_1
XFILLER_150_440 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11116_ _11115_/B _11115_/C _17469_/D _11115_/A vssd1 vssd1 vccd1 vccd1 _11116_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_68_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12096_ _12096_/A _12096_/B vssd1 vssd1 vccd1 vccd1 _12098_/C sky130_fd_sc_hd__xnor2_1
X_16973_ _13993_/B _16868_/A _16974_/A vssd1 vssd1 vccd1 vccd1 _16973_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_111_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11047_ _11048_/A _11048_/B vssd1 vssd1 vccd1 vccd1 _11047_/Y sky130_fd_sc_hd__nor2_1
X_15924_ _16036_/A _15924_/B vssd1 vssd1 vccd1 vccd1 _15926_/B sky130_fd_sc_hd__or2_1
XFILLER_77_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput9 i_wb_addr[15] vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__clkbuf_1
X_15855_ _15855_/A _15855_/B vssd1 vssd1 vccd1 vccd1 _15858_/A sky130_fd_sc_hd__xnor2_1
X_14806_ _14806_/A _15456_/A vssd1 vssd1 vccd1 vccd1 _14806_/X sky130_fd_sc_hd__or2_1
X_15786_ _15786_/A _15786_/B vssd1 vssd1 vccd1 vccd1 _15788_/B sky130_fd_sc_hd__or2_1
X_12998_ _12997_/A _12997_/B _12997_/C vssd1 vssd1 vccd1 vccd1 _12999_/B sky130_fd_sc_hd__o21ai_1
XFILLER_45_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17525_ fanout943/X _17525_/D vssd1 vssd1 vccd1 vccd1 _17525_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14737_ _17167_/A _14739_/B vssd1 vssd1 vccd1 vccd1 _14737_/X sky130_fd_sc_hd__or2_1
X_11949_ _09016_/A _09016_/Y _11947_/X _11948_/Y vssd1 vssd1 vccd1 vccd1 _11998_/A
+ sky130_fd_sc_hd__a211oi_2
XTAP_2980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17456_ fanout953/X _17456_/D vssd1 vssd1 vccd1 vccd1 _17456_/Q sky130_fd_sc_hd__dfxtp_1
X_14668_ _14735_/A1 _12394_/A _13625_/Y _12853_/X vssd1 vssd1 vccd1 vccd1 _14668_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_32_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16407_ _16407_/A vssd1 vssd1 vccd1 vccd1 _17561_/D sky130_fd_sc_hd__inv_2
X_13619_ _13619_/A _13619_/B vssd1 vssd1 vccd1 vccd1 _13621_/B sky130_fd_sc_hd__nand2_1
X_17387_ _17387_/A _17389_/B vssd1 vssd1 vccd1 vccd1 _17387_/X sky130_fd_sc_hd__or2_1
X_14599_ _14680_/A _14599_/B _14738_/B _14708_/D vssd1 vssd1 vccd1 vccd1 _14600_/B
+ sky130_fd_sc_hd__and4_1
X_16338_ _16339_/A _16339_/B _16339_/C vssd1 vssd1 vccd1 vccd1 _16444_/A sky130_fd_sc_hd__a21oi_1
XFILLER_9_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_938 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16269_ _16270_/A _16270_/B _16270_/C vssd1 vssd1 vccd1 vccd1 _16271_/A sky130_fd_sc_hd__o21a_1
XFILLER_173_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_930 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_621 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_142 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_527 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09712_ _10255_/A _10932_/B vssd1 vssd1 vccd1 vccd1 _09852_/A sky130_fd_sc_hd__nand2_2
XFILLER_142_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09643_ _10560_/A _09937_/B _09643_/C vssd1 vssd1 vccd1 vccd1 _09793_/A sky130_fd_sc_hd__and3_1
XFILLER_55_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09574_ _09574_/A _09574_/B _09574_/C vssd1 vssd1 vccd1 vccd1 _09575_/C sky130_fd_sc_hd__or3_1
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_276 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09008_ _09009_/A _09009_/B vssd1 vssd1 vccd1 vccd1 _09010_/A sky130_fd_sc_hd__or2_1
XFILLER_3_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10280_ _10266_/X _10267_/Y _10275_/X _10388_/A vssd1 vssd1 vccd1 vccd1 _10283_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_117_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_974 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout540 _15237_/A1 vssd1 vssd1 vccd1 vccd1 _11506_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout551 _09755_/B vssd1 vssd1 vccd1 vccd1 _11930_/B sky130_fd_sc_hd__buf_2
XFILLER_116_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout562 _13516_/S vssd1 vssd1 vccd1 vccd1 _13831_/S sky130_fd_sc_hd__buf_2
X_13970_ _13971_/A _13971_/B vssd1 vssd1 vccd1 vccd1 _14058_/B sky130_fd_sc_hd__nand2_1
Xfanout573 fanout578/X vssd1 vssd1 vccd1 vccd1 _11470_/A sky130_fd_sc_hd__clkbuf_2
Xfanout584 _17512_/Q vssd1 vssd1 vccd1 vccd1 _17164_/B sky130_fd_sc_hd__buf_2
XFILLER_59_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout595 _14954_/A vssd1 vssd1 vccd1 vccd1 _14958_/A sky130_fd_sc_hd__buf_2
XFILLER_18_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12921_ _12920_/A _12920_/B _12920_/C vssd1 vssd1 vccd1 vccd1 _12933_/B sky130_fd_sc_hd__a21oi_2
XFILLER_73_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15640_ _16812_/A _16591_/B vssd1 vssd1 vccd1 vccd1 _16419_/A sky130_fd_sc_hd__nand2_1
XFILLER_62_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12852_ _13831_/S _12852_/B vssd1 vssd1 vccd1 vccd1 _12852_/X sky130_fd_sc_hd__or2_2
XTAP_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11803_ _12054_/A _10431_/B _10309_/C vssd1 vssd1 vccd1 vccd1 _11804_/B sky130_fd_sc_hd__a21o_1
X_15571_ _15486_/A _15486_/B _15483_/Y vssd1 vssd1 vccd1 vccd1 _15573_/B sky130_fd_sc_hd__o21a_1
X_12783_ _12631_/A _12631_/Y _12781_/X _12938_/B vssd1 vssd1 vccd1 vccd1 _12825_/A
+ sky130_fd_sc_hd__o211a_1
XTAP_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17310_ _12129_/B _17322_/A2 _17309_/X _17358_/C1 vssd1 vssd1 vccd1 vccd1 _17484_/D
+ sky130_fd_sc_hd__o211a_1
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11734_ _11731_/B _11729_/C _11729_/B vssd1 vssd1 vccd1 vccd1 _11736_/B sky130_fd_sc_hd__o21a_1
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14522_ _14519_/X _14520_/Y _14463_/B _14465_/A vssd1 vssd1 vccd1 vccd1 _14523_/B
+ sky130_fd_sc_hd__o211ai_1
XTAP_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17241_ _17557_/Q _17292_/B vssd1 vssd1 vccd1 vccd1 _17241_/X sky130_fd_sc_hd__and2_1
X_11665_ _11673_/A _11673_/B vssd1 vssd1 vccd1 vccd1 _11674_/A sky130_fd_sc_hd__and2_1
X_14453_ _14454_/A _14454_/B vssd1 vssd1 vccd1 vccd1 _14509_/C sky130_fd_sc_hd__nand2_1
XFILLER_30_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10616_ _10719_/C _10508_/D _10509_/A _10507_/Y vssd1 vssd1 vccd1 vccd1 _10617_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_13404_ _13745_/B _13738_/B _13735_/D _13852_/A vssd1 vssd1 vccd1 vccd1 _13406_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_168_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17172_ input69/X input68/X input35/X vssd1 vssd1 vccd1 vccd1 _17172_/Y sky130_fd_sc_hd__nand3b_4
X_14384_ _16913_/C _14385_/B _14509_/A vssd1 vssd1 vccd1 vccd1 _14386_/A sky130_fd_sc_hd__a21oi_1
X_11596_ _11630_/A _15116_/B _11628_/B _11593_/Y vssd1 vssd1 vccd1 vccd1 _11598_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_128_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13335_ _13897_/A _13968_/B vssd1 vssd1 vccd1 vccd1 _13337_/C sky130_fd_sc_hd__nand2_1
X_16123_ _16304_/A _16112_/X _16113_/Y _16122_/X _16111_/X vssd1 vssd1 vccd1 vccd1
+ _16123_/X sky130_fd_sc_hd__o311a_1
X_10547_ _10547_/A _10547_/B _10547_/C vssd1 vssd1 vccd1 vccd1 _10671_/A sky130_fd_sc_hd__or3_1
XFILLER_6_553 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16054_ _16760_/A _16054_/B vssd1 vssd1 vccd1 vccd1 _16827_/D sky130_fd_sc_hd__nand2_2
X_13266_ _13266_/A _13266_/B vssd1 vssd1 vccd1 vccd1 _13271_/A sky130_fd_sc_hd__xnor2_1
X_10478_ _10478_/A _10478_/B vssd1 vssd1 vccd1 vccd1 _10480_/A sky130_fd_sc_hd__nor2_1
XFILLER_6_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12217_ _12848_/S _12217_/B vssd1 vssd1 vccd1 vccd1 _12218_/A sky130_fd_sc_hd__nor2_2
X_15005_ _14941_/X _15002_/X _15003_/X _15004_/Y _17156_/B vssd1 vssd1 vccd1 vccd1
+ _15005_/X sky130_fd_sc_hd__a311o_1
X_13197_ _13197_/A _13197_/B vssd1 vssd1 vccd1 vccd1 _13199_/C sky130_fd_sc_hd__xnor2_1
XFILLER_97_803 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12148_ _12148_/A _12148_/B _12148_/C vssd1 vssd1 vccd1 vccd1 _12149_/B sky130_fd_sc_hd__and3_1
XFILLER_111_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16956_ _16900_/A _16900_/C _16900_/B vssd1 vssd1 vccd1 vccd1 _16958_/B sky130_fd_sc_hd__a21bo_1
X_12079_ _17393_/A _12079_/B vssd1 vssd1 vccd1 vccd1 _12080_/B sky130_fd_sc_hd__nand2_1
XFILLER_38_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15907_ _15898_/A _16806_/A2 _15887_/Y _15906_/X vssd1 vssd1 vccd1 vccd1 _15908_/A
+ sky130_fd_sc_hd__a22o_1
X_16887_ _16887_/A _16887_/B vssd1 vssd1 vccd1 vccd1 _16888_/C sky130_fd_sc_hd__or2_1
XFILLER_2_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15838_ _15741_/A _15741_/B _15731_/X vssd1 vssd1 vccd1 vccd1 _15841_/B sky130_fd_sc_hd__o21a_1
XFILLER_24_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15769_ _15769_/A _15769_/B _15769_/C vssd1 vssd1 vccd1 vccd1 _15776_/B sky130_fd_sc_hd__nor3_1
XFILLER_33_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17508_ fanout944/X _17508_/D vssd1 vssd1 vccd1 vccd1 _17508_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_61_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09290_ _09290_/A _09290_/B _09290_/C vssd1 vssd1 vccd1 vccd1 _09291_/C sky130_fd_sc_hd__nand3_1
XFILLER_162_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17439_ fanout937/X _17439_/D vssd1 vssd1 vccd1 vccd1 _17439_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_14 _17081_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_25 _17531_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_36 _17442_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_47 _17381_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_58 fanout772/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_69 _15151_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput110 _17438_/Q vssd1 vssd1 vccd1 vccd1 o_wb_data[4] sky130_fd_sc_hd__clkbuf_1
XFILLER_133_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_988 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_446 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09626_ _09626_/A _09629_/B _09626_/C vssd1 vssd1 vccd1 vccd1 _09773_/A sky130_fd_sc_hd__and3_1
XFILLER_56_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09557_ _17393_/A _09557_/B vssd1 vssd1 vccd1 vccd1 _09558_/B sky130_fd_sc_hd__nand2_1
XFILLER_43_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09488_ _09388_/A _09486_/Y _09484_/B _09460_/X vssd1 vssd1 vccd1 vccd1 _09488_/Y
+ sky130_fd_sc_hd__o211ai_1
XFILLER_62_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11450_ _11403_/B _11400_/B _11400_/C vssd1 vssd1 vccd1 vccd1 _11451_/B sky130_fd_sc_hd__a21oi_1
Xwire215 wire215/A vssd1 vssd1 vccd1 vccd1 wire215/X sky130_fd_sc_hd__clkbuf_1
XFILLER_137_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10401_ _10402_/A _10402_/B _10402_/C vssd1 vssd1 vccd1 vccd1 _10405_/B sky130_fd_sc_hd__and3_1
X_11381_ _11380_/A _11426_/A vssd1 vssd1 vccd1 vccd1 _11383_/B sky130_fd_sc_hd__nand2b_1
XFILLER_109_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13120_ _13120_/A _13120_/B vssd1 vssd1 vccd1 vccd1 _13121_/C sky130_fd_sc_hd__xor2_1
XFILLER_109_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10332_ _10333_/B _10333_/A vssd1 vssd1 vccd1 vccd1 _10332_/X sky130_fd_sc_hd__and2b_1
XFILLER_3_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13051_ _13182_/A _13051_/B _13948_/C _13051_/D vssd1 vssd1 vccd1 vccd1 _13314_/A
+ sky130_fd_sc_hd__and4_1
X_10263_ _10249_/Y _10262_/X _10134_/Y _10231_/X vssd1 vssd1 vccd1 vccd1 _10263_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_87_22 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12002_ _09250_/Y _09255_/B _12200_/A _12001_/Y vssd1 vssd1 vccd1 vccd1 _12200_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_127_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10194_ _10194_/A _10194_/B _10194_/C vssd1 vssd1 vccd1 vccd1 _10214_/A sky130_fd_sc_hd__nor3_1
X_16810_ _15801_/A _15658_/Y _16662_/D _16808_/X vssd1 vssd1 vccd1 vccd1 _16811_/B
+ sky130_fd_sc_hd__o31a_1
Xfanout370 _12487_/A vssd1 vssd1 vccd1 vccd1 _09797_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_94_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout381 _12788_/A vssd1 vssd1 vccd1 vccd1 _13897_/A sky130_fd_sc_hd__buf_2
XFILLER_47_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16741_ _16715_/Y _16717_/Y _16853_/A vssd1 vssd1 vccd1 vccd1 _16787_/A sky130_fd_sc_hd__o21ai_1
Xfanout392 _14772_/A vssd1 vssd1 vccd1 vccd1 _12795_/A sky130_fd_sc_hd__buf_4
XFILLER_98_1010 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13953_ _14044_/A vssd1 vssd1 vccd1 vccd1 _14134_/A sky130_fd_sc_hd__inv_2
XFILLER_46_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_94 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12904_ _13051_/B _13051_/D vssd1 vssd1 vccd1 vccd1 _13182_/C sky130_fd_sc_hd__nand2_1
XFILLER_59_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16672_ _16673_/A _16673_/B vssd1 vssd1 vccd1 vccd1 _16751_/B sky130_fd_sc_hd__nand2_1
XFILLER_35_928 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13884_ _13885_/B _13885_/A vssd1 vssd1 vccd1 vccd1 _13986_/B sky130_fd_sc_hd__and2b_1
XTAP_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15623_ _15623_/A _15623_/B vssd1 vssd1 vccd1 vccd1 _15623_/X sky130_fd_sc_hd__xor2_1
X_12835_ _12991_/B _12834_/B _12834_/C vssd1 vssd1 vccd1 vccd1 _12835_/X sky130_fd_sc_hd__o21a_1
XTAP_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15554_ _15645_/B _15555_/B vssd1 vssd1 vccd1 vccd1 _15554_/Y sky130_fd_sc_hd__nor2_1
XFILLER_43_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12766_ _12766_/A _12928_/B _12766_/C vssd1 vssd1 vccd1 vccd1 _12920_/B sky130_fd_sc_hd__or3_2
XTAP_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14505_ _14505_/A _14505_/B vssd1 vssd1 vccd1 vccd1 _14506_/B sky130_fd_sc_hd__and2_1
X_11717_ _11717_/A _16295_/A _16206_/B vssd1 vssd1 vccd1 vccd1 _11717_/X sky130_fd_sc_hd__and3_1
XTAP_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15485_ _16317_/B _16536_/A vssd1 vssd1 vccd1 vccd1 _15486_/B sky130_fd_sc_hd__nand2_1
X_12697_ _12379_/B _13004_/A _12695_/X vssd1 vssd1 vccd1 vccd1 _12698_/B sky130_fd_sc_hd__o21a_1
X_17224_ _17442_/Q _17275_/A2 _17222_/X _17223_/X _17364_/C1 vssd1 vssd1 vccd1 vccd1
+ _17442_/D sky130_fd_sc_hd__o221a_1
X_11648_ _11648_/A _11648_/B vssd1 vssd1 vccd1 vccd1 _11686_/A sky130_fd_sc_hd__xnor2_1
X_14436_ _14554_/A _14641_/C _14437_/C vssd1 vssd1 vccd1 vccd1 _14438_/A sky130_fd_sc_hd__a21oi_1
XFILLER_174_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput12 i_wb_addr[18] vssd1 vssd1 vccd1 vccd1 input12/X sky130_fd_sc_hd__clkbuf_1
Xinput23 i_wb_addr[28] vssd1 vssd1 vccd1 vccd1 input23/X sky130_fd_sc_hd__clkbuf_1
XFILLER_174_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput34 i_wb_addr[9] vssd1 vssd1 vccd1 vccd1 input34/X sky130_fd_sc_hd__clkbuf_1
Xinput45 i_wb_data[18] vssd1 vssd1 vccd1 vccd1 input45/X sky130_fd_sc_hd__clkbuf_1
X_17155_ _17152_/Y _17153_/X _17133_/A _17136_/X vssd1 vssd1 vccd1 vccd1 _17156_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_171_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11579_ _11579_/A _11579_/B _11579_/C vssd1 vssd1 vccd1 vccd1 _11614_/A sky130_fd_sc_hd__nand3_1
X_14367_ _14367_/A _17023_/A vssd1 vssd1 vccd1 vccd1 _14368_/C sky130_fd_sc_hd__xor2_1
Xinput56 i_wb_data[28] vssd1 vssd1 vccd1 vccd1 input56/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput67 i_wb_data[9] vssd1 vssd1 vccd1 vccd1 input67/X sky130_fd_sc_hd__clkbuf_1
X_16106_ _16106_/A _16106_/B vssd1 vssd1 vccd1 vccd1 _16106_/Y sky130_fd_sc_hd__nand2_1
XFILLER_115_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13318_ _13189_/A _13189_/Y _13316_/Y _13431_/B vssd1 vssd1 vccd1 vccd1 _13329_/A
+ sky130_fd_sc_hd__a211o_1
X_17086_ _17086_/A _17086_/B vssd1 vssd1 vccd1 vccd1 _17088_/C sky130_fd_sc_hd__and2_1
X_14298_ _14214_/A _14216_/B _14214_/B vssd1 vssd1 vccd1 vccd1 _14306_/A sky130_fd_sc_hd__o21ba_1
X_16037_ _16416_/A _16041_/B _15935_/A _15933_/B vssd1 vssd1 vccd1 vccd1 _16046_/A
+ sky130_fd_sc_hd__o31a_1
XFILLER_171_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13249_ _13249_/A _13249_/B _13249_/C _13249_/D vssd1 vssd1 vccd1 vccd1 _13249_/Y
+ sky130_fd_sc_hd__nand4_2
XFILLER_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_302 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08790_ _08792_/D vssd1 vssd1 vccd1 vccd1 _08790_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_96_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16939_ _16983_/A _16939_/B vssd1 vssd1 vccd1 vccd1 _16986_/A sky130_fd_sc_hd__or2_1
XFILLER_84_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09411_ _09411_/A _09411_/B _09417_/B vssd1 vssd1 vccd1 vccd1 _09434_/B sky130_fd_sc_hd__or3_1
XFILLER_16_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09342_ _09342_/A _09342_/B vssd1 vssd1 vccd1 vccd1 _09344_/C sky130_fd_sc_hd__nor2_1
XFILLER_21_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09273_ _09273_/A _09273_/B vssd1 vssd1 vccd1 vccd1 _09274_/B sky130_fd_sc_hd__nor2_1
XFILLER_21_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_863 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08988_ _17425_/A _08988_/B _11920_/D _09362_/D vssd1 vssd1 vccd1 vccd1 _08989_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_87_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10950_ _10857_/Y _10863_/B _10951_/A _10949_/Y vssd1 vssd1 vccd1 vccd1 _11065_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_28_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09609_ _09610_/A _09610_/C vssd1 vssd1 vccd1 vccd1 _09614_/B sky130_fd_sc_hd__nor2_1
X_10881_ _10883_/B _10883_/C _10883_/A vssd1 vssd1 vccd1 vccd1 _10881_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_83_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12620_ _17421_/A _12923_/D vssd1 vssd1 vccd1 vccd1 _12621_/B sky130_fd_sc_hd__nand2_1
XFILLER_19_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12551_ _11827_/X _11854_/C _12845_/S vssd1 vssd1 vccd1 vccd1 _12552_/B sky130_fd_sc_hd__mux2_1
XFILLER_8_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11502_ _11502_/A _11502_/B _11502_/C vssd1 vssd1 vccd1 vccd1 _11543_/A sky130_fd_sc_hd__nor3_2
XFILLER_129_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15270_ _15270_/A _15270_/B _15270_/C vssd1 vssd1 vccd1 vccd1 _15270_/X sky130_fd_sc_hd__or3_1
X_12482_ _12312_/A _12314_/A _12479_/Y _12480_/X vssd1 vssd1 vccd1 vccd1 _12522_/A
+ sky130_fd_sc_hd__a211oi_1
XFILLER_40_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11433_ _11433_/A _11433_/B _11433_/C vssd1 vssd1 vccd1 vccd1 _11477_/A sky130_fd_sc_hd__nand3_1
X_14221_ _14221_/A _14221_/B _14221_/C vssd1 vssd1 vccd1 vccd1 _14222_/B sky130_fd_sc_hd__or3_1
XFILLER_22_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14152_ _14153_/B _14426_/D _14360_/D _14153_/A vssd1 vssd1 vccd1 vccd1 _14154_/A
+ sky130_fd_sc_hd__a22oi_1
X_11364_ _11364_/A _11364_/B vssd1 vssd1 vccd1 vccd1 _11447_/B sky130_fd_sc_hd__xnor2_1
XFILLER_99_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13103_ _13103_/A _13103_/B vssd1 vssd1 vccd1 vccd1 _13106_/A sky130_fd_sc_hd__xnor2_1
XFILLER_98_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10315_ _10315_/A _10315_/B _10315_/C vssd1 vssd1 vccd1 vccd1 _10315_/X sky130_fd_sc_hd__and3_1
X_14083_ _14387_/A _14366_/B _14084_/A vssd1 vssd1 vccd1 vccd1 _14173_/B sky130_fd_sc_hd__and3_1
X_11295_ _11295_/A _11295_/B vssd1 vssd1 vccd1 vccd1 _11345_/B sky130_fd_sc_hd__xnor2_1
XFILLER_152_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13034_ _13414_/B _13035_/C _13908_/B _13035_/A vssd1 vssd1 vccd1 vccd1 _13036_/A
+ sky130_fd_sc_hd__a22oi_1
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10246_ _10246_/A _10246_/B vssd1 vssd1 vccd1 vccd1 _10358_/B sky130_fd_sc_hd__xor2_1
XFILLER_3_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10177_ _10177_/A _10177_/B _10289_/A vssd1 vssd1 vccd1 vccd1 _10188_/B sky130_fd_sc_hd__nand3_1
XFILLER_121_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_338 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14985_ _10431_/B _14863_/B _14863_/A _14864_/A _09925_/A _15095_/B vssd1 vssd1 vccd1
+ vccd1 _14986_/B sky130_fd_sc_hd__mux4_1
X_16724_ _16643_/Y _16647_/A _16723_/B _16723_/A _16721_/Y vssd1 vssd1 vccd1 vccd1
+ _16791_/B sky130_fd_sc_hd__a221o_1
X_13936_ _13936_/A _13936_/B _13728_/Y vssd1 vssd1 vccd1 vccd1 _13936_/Y sky130_fd_sc_hd__nor3b_1
XFILLER_75_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16655_ _16649_/A _17163_/A2 _16654_/X vssd1 vssd1 vccd1 vccd1 _16655_/X sky130_fd_sc_hd__o21ba_1
X_13867_ _13867_/A _13867_/B vssd1 vssd1 vccd1 vccd1 _13869_/A sky130_fd_sc_hd__nor2_1
XFILLER_62_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_717 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15606_ _15607_/A _15607_/B vssd1 vssd1 vccd1 vccd1 _15606_/Y sky130_fd_sc_hd__nand2_1
XFILLER_16_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12818_ _12820_/A _12820_/B _12820_/C vssd1 vssd1 vccd1 vccd1 _12821_/A sky130_fd_sc_hd__a21oi_1
X_16586_ _16571_/A _17170_/B1 _16575_/X _16585_/X vssd1 vssd1 vccd1 vccd1 _17563_/D
+ sky130_fd_sc_hd__a22oi_1
X_13798_ _13906_/B _13798_/B vssd1 vssd1 vccd1 vccd1 _13800_/C sky130_fd_sc_hd__nand2_1
XFILLER_31_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15537_ _16011_/A _15537_/B vssd1 vssd1 vccd1 vccd1 _15537_/X sky130_fd_sc_hd__or2_1
X_12749_ _13182_/A _13037_/B vssd1 vssd1 vccd1 vccd1 _12749_/Y sky130_fd_sc_hd__nand2_1
XFILLER_31_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1046 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15468_ _15446_/Y _15447_/X _15467_/X _15445_/X vssd1 vssd1 vccd1 vccd1 _15468_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_147_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_852 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17207_ _17578_/Q _17273_/A2 _17273_/B1 vssd1 vssd1 vccd1 vccd1 _17207_/X sky130_fd_sc_hd__a21o_1
XFILLER_8_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14419_ _14533_/A _14419_/B vssd1 vssd1 vccd1 vccd1 _14419_/Y sky130_fd_sc_hd__nand2_1
X_15399_ _16315_/B _16410_/A _16041_/B _15820_/A vssd1 vssd1 vccd1 vccd1 _15400_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_128_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17138_ _17138_/A _17138_/B vssd1 vssd1 vccd1 vccd1 _17138_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_7_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17069_ _14434_/Y _14764_/Y _14825_/Y _17023_/A vssd1 vssd1 vccd1 vccd1 _17069_/Y
+ sky130_fd_sc_hd__o211ai_1
X_09960_ _09960_/A _09960_/B _09960_/C vssd1 vssd1 vccd1 vccd1 _09960_/Y sky130_fd_sc_hd__nand3_1
XFILLER_89_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08911_ _17381_/A _09321_/D _08843_/A _08841_/Y vssd1 vssd1 vccd1 vccd1 _08912_/B
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09891_ _09891_/A _09891_/B vssd1 vssd1 vccd1 vccd1 _09906_/A sky130_fd_sc_hd__nand2_1
XFILLER_97_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08842_ _08843_/A _08841_/Y _17381_/A _09321_/D vssd1 vssd1 vccd1 vccd1 _08912_/A
+ sky130_fd_sc_hd__and4bb_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08773_ _08773_/A _08804_/A vssd1 vssd1 vccd1 vccd1 _08780_/B sky130_fd_sc_hd__nor2_1
XFILLER_69_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_820 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_522 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_780 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09325_ _09755_/A _09325_/B _09926_/B _10180_/B vssd1 vssd1 vccd1 vccd1 _09462_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_138_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09256_ _09256_/A _09256_/B vssd1 vssd1 vccd1 vccd1 _09395_/A sky130_fd_sc_hd__xnor2_1
XFILLER_138_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09187_ _17409_/A _09555_/D vssd1 vssd1 vccd1 vccd1 _09189_/C sky130_fd_sc_hd__nand2_1
XFILLER_153_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10100_ _10090_/A _10088_/X _10081_/A _10084_/A vssd1 vssd1 vccd1 vccd1 _10101_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_68_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11080_ _11080_/A _11080_/B _11080_/C _11080_/D vssd1 vssd1 vccd1 vccd1 _11145_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_89_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10031_ _10010_/A _10027_/C _10030_/Y _09910_/B vssd1 vssd1 vccd1 vccd1 _10033_/A
+ sky130_fd_sc_hd__a211oi_1
XFILLER_88_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14770_ _14770_/A _14864_/A vssd1 vssd1 vccd1 vccd1 _16864_/B sky130_fd_sc_hd__or2_1
X_11982_ _11982_/A _11982_/B vssd1 vssd1 vccd1 vccd1 _11984_/B sky130_fd_sc_hd__xnor2_1
XFILLER_56_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_820 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13721_ _13577_/B _13579_/B _13577_/A vssd1 vssd1 vccd1 vccd1 _13723_/B sky130_fd_sc_hd__o21ba_1
X_10933_ _10933_/A _11122_/B _10933_/C _10933_/D vssd1 vssd1 vccd1 vccd1 _10935_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_17_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1046 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16440_ _16331_/A _16331_/B _16345_/A vssd1 vssd1 vccd1 vccd1 _16442_/B sky130_fd_sc_hd__a21o_1
X_10864_ _10863_/B _10863_/C _10863_/A vssd1 vssd1 vccd1 vccd1 _10864_/Y sky130_fd_sc_hd__o21ai_1
X_13652_ _13652_/A _13652_/B vssd1 vssd1 vccd1 vccd1 _13655_/B sky130_fd_sc_hd__xnor2_1
XFILLER_31_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12603_ _12603_/A _12603_/B vssd1 vssd1 vccd1 vccd1 _12605_/B sky130_fd_sc_hd__xnor2_1
XPHY_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16371_ _16372_/B _16372_/A vssd1 vssd1 vccd1 vccd1 _16371_/Y sky130_fd_sc_hd__nand2b_1
XPHY_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10795_ _10884_/A _10794_/B _10794_/A vssd1 vssd1 vccd1 vccd1 _10860_/B sky130_fd_sc_hd__o21ba_1
XPHY_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13583_ _14155_/A _14050_/D vssd1 vssd1 vccd1 vccd1 _13584_/B sky130_fd_sc_hd__nand2_1
XFILLER_13_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15322_ _16207_/B _15303_/Y _15321_/X _15301_/Y vssd1 vssd1 vccd1 vccd1 _15322_/X
+ sky130_fd_sc_hd__o211a_1
XPHY_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12534_ _12534_/A _12534_/B vssd1 vssd1 vccd1 vccd1 _12536_/A sky130_fd_sc_hd__xnor2_1
XPHY_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15253_ _14988_/Y _14999_/Y _15384_/S vssd1 vssd1 vccd1 vccd1 _15253_/X sky130_fd_sc_hd__mux2_1
X_12465_ _17421_/A _12770_/D vssd1 vssd1 vccd1 vccd1 _12467_/B sky130_fd_sc_hd__nand2_1
XFILLER_173_939 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_8 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14204_ _14204_/A _14279_/B vssd1 vssd1 vccd1 vccd1 _14278_/B sky130_fd_sc_hd__or2_1
X_11416_ _11416_/A _11416_/B vssd1 vssd1 vccd1 vccd1 _11418_/B sky130_fd_sc_hd__or2_1
XFILLER_126_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15184_ _14790_/Y _14929_/X _15713_/B1 _15175_/B vssd1 vssd1 vccd1 vccd1 _15184_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_12396_ _12388_/X _14210_/A _17371_/A vssd1 vssd1 vccd1 vccd1 _12396_/X sky130_fd_sc_hd__mux2_1
XFILLER_126_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11347_ _11347_/A _11347_/B vssd1 vssd1 vccd1 vccd1 _11348_/B sky130_fd_sc_hd__nand2_1
XFILLER_141_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14135_ _14134_/A _14134_/B _14134_/C vssd1 vssd1 vccd1 vccd1 _14136_/B sky130_fd_sc_hd__o21a_1
XFILLER_4_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11278_ _11561_/A _14893_/B _11387_/C vssd1 vssd1 vccd1 vccd1 _11283_/B sky130_fd_sc_hd__and3_1
X_14066_ _14066_/A _14066_/B vssd1 vssd1 vccd1 vccd1 _14068_/B sky130_fd_sc_hd__xnor2_1
X_13017_ _13632_/B _14063_/C _14213_/D _13735_/A vssd1 vssd1 vccd1 vccd1 _13019_/A
+ sky130_fd_sc_hd__a22oi_1
X_10229_ _10192_/B _10207_/B _10192_/D _10193_/A vssd1 vssd1 vccd1 vccd1 _10229_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_140_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14968_ _14966_/X _14967_/X _15147_/D vssd1 vssd1 vccd1 vccd1 _14968_/X sky130_fd_sc_hd__a21o_1
XFILLER_81_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16707_ _16542_/A _16626_/B _16624_/X vssd1 vssd1 vccd1 vccd1 _16709_/B sky130_fd_sc_hd__a21oi_1
X_13919_ _14018_/B _13919_/B vssd1 vssd1 vccd1 vccd1 _13921_/C sky130_fd_sc_hd__nand2_1
XFILLER_47_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14899_ _15314_/A _14906_/B _14899_/C vssd1 vssd1 vccd1 vccd1 _14899_/X sky130_fd_sc_hd__or3_2
X_16638_ _16638_/A _16638_/B vssd1 vssd1 vccd1 vccd1 _16854_/C sky130_fd_sc_hd__xnor2_2
XFILLER_63_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16569_ _16568_/A _16568_/B _16207_/B _16568_/Y vssd1 vssd1 vccd1 vccd1 _16569_/X
+ sky130_fd_sc_hd__a211o_1
X_09110_ _09110_/A _09110_/B vssd1 vssd1 vccd1 vccd1 _09111_/B sky130_fd_sc_hd__nor2_1
XFILLER_13_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_958 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09041_ _09043_/A _17081_/B vssd1 vssd1 vccd1 vccd1 _09041_/Y sky130_fd_sc_hd__nor2_1
XFILLER_159_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xmax_cap120 _13492_/A vssd1 vssd1 vccd1 vccd1 _13607_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_172_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09943_ _09942_/A _10062_/B _10062_/C vssd1 vssd1 vccd1 vccd1 _09943_/Y sky130_fd_sc_hd__a21oi_1
Xfanout903 fanout904/X vssd1 vssd1 vccd1 vccd1 _10954_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_132_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout914 _17273_/B1 vssd1 vssd1 vccd1 vccd1 _17282_/B1 sky130_fd_sc_hd__clkbuf_2
Xfanout925 _17358_/C1 vssd1 vssd1 vccd1 vccd1 _17388_/C1 sky130_fd_sc_hd__buf_2
Xfanout936 fanout937/X vssd1 vssd1 vccd1 vccd1 fanout936/X sky130_fd_sc_hd__clkbuf_2
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout947 fanout948/X vssd1 vssd1 vccd1 vccd1 fanout947/X sky130_fd_sc_hd__clkbuf_2
X_09874_ _14784_/A _10016_/D _10146_/B _09873_/A vssd1 vssd1 vccd1 vccd1 _09874_/Y
+ sky130_fd_sc_hd__a22oi_1
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_934 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08825_ _17389_/A _09446_/D _09042_/B _17391_/A vssd1 vssd1 vccd1 vccd1 _08826_/B
+ sky130_fd_sc_hd__a22oi_1
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08756_ _08757_/B _08757_/A vssd1 vssd1 vccd1 vccd1 _11877_/A sky130_fd_sc_hd__nand2b_1
XTAP_2606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_1000 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09308_ _09316_/A _09296_/Y _09303_/X _09439_/A vssd1 vssd1 vccd1 vccd1 _09311_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_70_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10580_ _10582_/A _10582_/B vssd1 vssd1 vccd1 vccd1 _10583_/A sky130_fd_sc_hd__or2_1
XFILLER_103_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09239_ _09239_/A _09239_/B vssd1 vssd1 vccd1 vccd1 _09240_/B sky130_fd_sc_hd__nor2_1
XFILLER_108_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12250_ _12250_/A _12250_/B vssd1 vssd1 vccd1 vccd1 _12252_/C sky130_fd_sc_hd__xnor2_1
XFILLER_119_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11201_ _11201_/A _11201_/B vssd1 vssd1 vccd1 vccd1 _16387_/A sky130_fd_sc_hd__xnor2_1
XFILLER_107_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12181_ _11978_/A _11980_/B _11978_/B vssd1 vssd1 vccd1 vccd1 _12182_/B sky130_fd_sc_hd__o21ba_1
XFILLER_119_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11132_ _11561_/A _11132_/B _11132_/C _15624_/A vssd1 vssd1 vccd1 vccd1 _11137_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_150_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11063_ _11061_/A _11061_/C _11077_/A vssd1 vssd1 vccd1 vccd1 _11065_/D sky130_fd_sc_hd__a21o_1
X_15940_ _16072_/B _15940_/B vssd1 vssd1 vccd1 vccd1 _15941_/B sky130_fd_sc_hd__nor2_1
XFILLER_95_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10014_ _10142_/A _14784_/A _10146_/B _10014_/D vssd1 vssd1 vccd1 vccd1 _10017_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_49_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15871_ _15871_/A _15871_/B vssd1 vssd1 vccd1 vccd1 _15872_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_444 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17610_ fanout950/X _17610_/D vssd1 vssd1 vccd1 vccd1 _17610_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_64_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14822_ _16864_/B _16865_/A _16864_/A vssd1 vssd1 vccd1 vccd1 _16918_/C sky130_fd_sc_hd__a21bo_1
XFILLER_76_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17541_ fanout944/X _17541_/D vssd1 vssd1 vccd1 vccd1 _17541_/Q sky130_fd_sc_hd__dfxtp_2
X_14753_ _14701_/A _14701_/B _14725_/Y _14752_/Y vssd1 vssd1 vccd1 vccd1 _14755_/B
+ sky130_fd_sc_hd__o31a_1
X_11965_ _11966_/B _11965_/B vssd1 vssd1 vccd1 vccd1 _11967_/A sky130_fd_sc_hd__nand2b_1
XFILLER_45_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13704_ _13908_/A _13704_/B vssd1 vssd1 vccd1 vccd1 _13705_/B sky130_fd_sc_hd__nand2_1
X_17472_ fanout955/X _17545_/Q vssd1 vssd1 vccd1 vccd1 _17472_/Q sky130_fd_sc_hd__dfxtp_1
X_10916_ _10808_/A _10807_/B _10807_/A vssd1 vssd1 vccd1 vccd1 _10918_/B sky130_fd_sc_hd__o21ba_1
XFILLER_45_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_823 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14684_ _14684_/A vssd1 vssd1 vccd1 vccd1 _14719_/B sky130_fd_sc_hd__inv_2
X_11896_ _11894_/Y _12138_/A _17375_/A _12447_/B vssd1 vssd1 vccd1 vccd1 _12138_/B
+ sky130_fd_sc_hd__and4bb_1
XFILLER_17_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16423_ _16423_/A _16509_/B vssd1 vssd1 vccd1 vccd1 _16423_/Y sky130_fd_sc_hd__nand2_1
XFILLER_60_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13635_ _13635_/A _13741_/A _13635_/C vssd1 vssd1 vccd1 vccd1 _13638_/A sky130_fd_sc_hd__or3_1
X_10847_ _10828_/A _10827_/B _10827_/A vssd1 vssd1 vccd1 vccd1 _10855_/A sky130_fd_sc_hd__o21ba_1
X_16354_ _16354_/A _16354_/B vssd1 vssd1 vccd1 vccd1 _16356_/A sky130_fd_sc_hd__nor2_1
X_13566_ _13897_/A _13691_/C vssd1 vssd1 vccd1 vccd1 _13568_/B sky130_fd_sc_hd__nand2_1
X_10778_ _10778_/A _11742_/A vssd1 vssd1 vccd1 vccd1 _10779_/B sky130_fd_sc_hd__nor2_1
XFILLER_12_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15305_ _15314_/A _15373_/B _15305_/C vssd1 vssd1 vccd1 vccd1 _15307_/B sky130_fd_sc_hd__and3b_1
X_12517_ _12517_/A _12517_/B vssd1 vssd1 vccd1 vccd1 _12518_/B sky130_fd_sc_hd__xnor2_1
XFILLER_173_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16285_ _16285_/A _16285_/B vssd1 vssd1 vccd1 vccd1 _16288_/A sky130_fd_sc_hd__xor2_1
XFILLER_145_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_416 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13497_ _13498_/B _13498_/A vssd1 vssd1 vccd1 vccd1 _13497_/X sky130_fd_sc_hd__and2b_1
XFILLER_9_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15236_ _15235_/B _15235_/C _15235_/A vssd1 vssd1 vccd1 vccd1 _15236_/X sky130_fd_sc_hd__a21o_1
XFILLER_161_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12448_ _12448_/A _12448_/B vssd1 vssd1 vccd1 vccd1 _12451_/A sky130_fd_sc_hd__xnor2_1
XFILLER_160_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15167_ _15089_/S _15687_/A _15170_/B vssd1 vssd1 vccd1 vccd1 _15169_/B sky130_fd_sc_hd__o21ai_1
XFILLER_141_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12379_ _12696_/A _12379_/B vssd1 vssd1 vccd1 vccd1 _12380_/B sky130_fd_sc_hd__or2_1
XFILLER_114_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_525 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14118_ _14119_/A _14119_/B _14117_/X vssd1 vssd1 vccd1 vccd1 _14279_/A sky130_fd_sc_hd__o21ba_1
XFILLER_119_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15098_ _17164_/D _15097_/X _15103_/S vssd1 vssd1 vccd1 vccd1 _15715_/B sky130_fd_sc_hd__mux2_1
XFILLER_113_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14049_ _14050_/B _14141_/D _14050_/D _13966_/A vssd1 vssd1 vccd1 vccd1 _14051_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_68_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09590_ _09894_/C _10311_/D _09473_/A _09465_/Y vssd1 vssd1 vccd1 vccd1 _09591_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_36_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_694 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_580 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09024_ _12068_/B _12340_/B _09267_/D _17403_/A vssd1 vssd1 vccd1 vccd1 _09024_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_129_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout700 _16654_/B2 vssd1 vssd1 vccd1 vccd1 _12871_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_104_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout711 _16571_/A vssd1 vssd1 vccd1 vccd1 _13968_/B sky130_fd_sc_hd__buf_4
Xfanout722 _17497_/Q vssd1 vssd1 vccd1 vccd1 _12077_/C sky130_fd_sc_hd__clkbuf_4
X_09926_ _15254_/S _09926_/B _09926_/C vssd1 vssd1 vccd1 vccd1 _09929_/A sky130_fd_sc_hd__and3_1
Xfanout733 _16298_/A vssd1 vssd1 vccd1 vccd1 _13208_/D sky130_fd_sc_hd__buf_4
Xfanout744 _14859_/B vssd1 vssd1 vccd1 vccd1 _14778_/B sky130_fd_sc_hd__buf_6
XFILLER_59_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_880 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout755 _17119_/A vssd1 vssd1 vccd1 vccd1 _16760_/A sky130_fd_sc_hd__clkbuf_2
Xfanout766 _16014_/A vssd1 vssd1 vccd1 vccd1 _15204_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout777 _16758_/A vssd1 vssd1 vccd1 vccd1 _16807_/A sky130_fd_sc_hd__clkbuf_4
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09857_ _09710_/Y _09856_/Y _09855_/X vssd1 vssd1 vccd1 vccd1 _09994_/A sky130_fd_sc_hd__a21o_1
Xfanout788 _11132_/C vssd1 vssd1 vccd1 vccd1 _16938_/A sky130_fd_sc_hd__clkbuf_4
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout799 fanout805/X vssd1 vssd1 vccd1 vccd1 _09557_/B sky130_fd_sc_hd__buf_2
XFILLER_105_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08808_ _08808_/A _08883_/A vssd1 vssd1 vccd1 vccd1 _08815_/B sky130_fd_sc_hd__nor2_1
XFILLER_58_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09788_ _09788_/A _09788_/B vssd1 vssd1 vccd1 vccd1 _09789_/B sky130_fd_sc_hd__and2_1
XTAP_3137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08739_ _17607_/Q _17608_/Q vssd1 vssd1 vccd1 vccd1 _14933_/A sky130_fd_sc_hd__nand2b_2
XFILLER_38_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_31 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11750_ _11750_/A _11750_/B vssd1 vssd1 vccd1 vccd1 _16795_/A sky130_fd_sc_hd__xor2_2
XFILLER_53_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_311 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10701_ _10701_/A _10701_/B vssd1 vssd1 vccd1 vccd1 _10708_/A sky130_fd_sc_hd__xor2_2
XTAP_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11681_ _11681_/A _11681_/B vssd1 vssd1 vccd1 vccd1 _15235_/B sky130_fd_sc_hd__or2_1
XTAP_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13420_ _13420_/A _13420_/B vssd1 vssd1 vccd1 vccd1 _13423_/C sky130_fd_sc_hd__xnor2_1
XFILLER_41_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10632_ _10632_/A _10632_/B _10632_/C _10632_/D vssd1 vssd1 vccd1 vccd1 _10632_/Y
+ sky130_fd_sc_hd__nand4_2
X_13351_ _14153_/B _13764_/D _13664_/D _13227_/A vssd1 vssd1 vccd1 vccd1 _13353_/A
+ sky130_fd_sc_hd__a22oi_1
X_10563_ _10563_/A _10563_/B vssd1 vssd1 vccd1 vccd1 _10564_/B sky130_fd_sc_hd__or2_1
XFILLER_155_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12302_ _17373_/A _12592_/C _12470_/B vssd1 vssd1 vccd1 vccd1 _12303_/B sky130_fd_sc_hd__and3_1
X_16070_ _16070_/A _16070_/B vssd1 vssd1 vccd1 vccd1 _16072_/C sky130_fd_sc_hd__xnor2_1
XFILLER_127_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10494_ _10601_/A _10493_/B _10493_/A vssd1 vssd1 vccd1 vccd1 _10496_/B sky130_fd_sc_hd__o21ba_1
XFILLER_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13282_ _13282_/A _13282_/B vssd1 vssd1 vccd1 vccd1 _13285_/A sky130_fd_sc_hd__xnor2_1
XFILLER_6_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15021_ _15402_/A _15402_/B vssd1 vssd1 vccd1 vccd1 _15734_/A sky130_fd_sc_hd__nand2_2
X_12233_ _12869_/A _13208_/C vssd1 vssd1 vccd1 vccd1 _12235_/C sky130_fd_sc_hd__and2_4
XFILLER_135_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12164_ _12163_/A _12163_/B _12163_/C vssd1 vssd1 vccd1 vccd1 _12165_/B sky130_fd_sc_hd__o21a_1
XFILLER_151_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11115_ _11115_/A _11115_/B _11115_/C _17469_/D vssd1 vssd1 vccd1 vccd1 _11118_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_68_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12095_ _12096_/A _12096_/B vssd1 vssd1 vccd1 vccd1 _12286_/B sky130_fd_sc_hd__nand2b_1
X_16972_ _16972_/A _16972_/B vssd1 vssd1 vccd1 vccd1 _16972_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_111_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_891 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11046_ _11046_/A _11046_/B vssd1 vssd1 vccd1 vccd1 _11048_/B sky130_fd_sc_hd__nand2_1
X_15923_ _15923_/A _15923_/B vssd1 vssd1 vccd1 vccd1 _15924_/B sky130_fd_sc_hd__and2_1
XFILLER_110_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15854_ _16536_/A _15854_/B vssd1 vssd1 vccd1 vccd1 _15855_/B sky130_fd_sc_hd__nand2_1
XFILLER_77_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_639 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_959 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14805_ _14805_/A _14805_/B _14805_/C vssd1 vssd1 vccd1 vccd1 _15456_/A sky130_fd_sc_hd__and3_1
XFILLER_80_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15785_ _15883_/B _15787_/B vssd1 vssd1 vccd1 vccd1 _15788_/A sky130_fd_sc_hd__or2_1
XFILLER_17_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12997_ _12997_/A _12997_/B _12997_/C vssd1 vssd1 vccd1 vccd1 _12999_/A sky130_fd_sc_hd__or3_1
X_17524_ fanout943/X _17524_/D vssd1 vssd1 vccd1 vccd1 _17524_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_55_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14736_ _14736_/A _14744_/A vssd1 vssd1 vccd1 vccd1 _14739_/B sky130_fd_sc_hd__nand2_1
X_11948_ _11917_/X _11918_/Y _12156_/B _11947_/D vssd1 vssd1 vccd1 vccd1 _11948_/Y
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_17_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_299 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17455_ fanout953/X _17455_/D vssd1 vssd1 vccd1 vccd1 _17455_/Q sky130_fd_sc_hd__dfxtp_1
X_14667_ _14734_/A _14667_/B vssd1 vssd1 vccd1 vccd1 _14667_/Y sky130_fd_sc_hd__nand2_1
X_11879_ _08760_/Y _16302_/A _08764_/A _08764_/B vssd1 vssd1 vccd1 vccd1 _11886_/A
+ sky130_fd_sc_hd__o22ai_4
XFILLER_33_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16406_ _16386_/Y _16389_/Y _16405_/X _17170_/B1 _16399_/A vssd1 vssd1 vccd1 vccd1
+ _16407_/A sky130_fd_sc_hd__a32o_1
X_13618_ _13618_/A _13618_/B vssd1 vssd1 vccd1 vccd1 _13729_/B sky130_fd_sc_hd__xnor2_1
XFILLER_158_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17386_ input38/X _17426_/A2 _17385_/X _17426_/C1 vssd1 vssd1 vccd1 vccd1 _17521_/D
+ sky130_fd_sc_hd__o211a_1
X_14598_ _14599_/B _14738_/B _14708_/D _14680_/A vssd1 vssd1 vccd1 vccd1 _14600_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_158_563 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16337_ _16337_/A _16337_/B vssd1 vssd1 vccd1 vccd1 _16339_/C sky130_fd_sc_hd__xnor2_1
X_13549_ _13662_/B _13547_/X _13425_/Y _13430_/A vssd1 vssd1 vccd1 vccd1 _13558_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_72_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16268_ _16268_/A _16268_/B vssd1 vssd1 vccd1 vccd1 _16270_/C sky130_fd_sc_hd__xnor2_1
X_15219_ _15220_/A _15220_/B vssd1 vssd1 vccd1 vccd1 _15287_/A sky130_fd_sc_hd__nand2b_1
X_16199_ _16200_/A _16200_/B _16200_/C vssd1 vssd1 vccd1 vccd1 _16382_/A sky130_fd_sc_hd__a21oi_1
XFILLER_142_942 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09711_ _10255_/A _10932_/B vssd1 vssd1 vccd1 vccd1 _09711_/X sky130_fd_sc_hd__and2_1
XFILLER_132_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09642_ _09642_/A _09642_/B vssd1 vssd1 vccd1 vccd1 _09643_/C sky130_fd_sc_hd__xnor2_1
XFILLER_56_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09573_ _09573_/A _09573_/B vssd1 vssd1 vccd1 vccd1 _09575_/B sky130_fd_sc_hd__xnor2_1
XFILLER_36_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_661 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_878 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_1000 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09007_ _09007_/A _09007_/B vssd1 vssd1 vccd1 vccd1 _09009_/B sky130_fd_sc_hd__xnor2_1
XFILLER_152_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_986 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout530 _17516_/Q vssd1 vssd1 vccd1 vccd1 _10970_/A sky130_fd_sc_hd__clkbuf_4
Xfanout541 _09899_/A vssd1 vssd1 vccd1 vccd1 _15237_/A1 sky130_fd_sc_hd__buf_2
Xfanout552 _17514_/Q vssd1 vssd1 vccd1 vccd1 _09755_/B sky130_fd_sc_hd__clkbuf_4
X_09909_ _09909_/A _09909_/B _09909_/C vssd1 vssd1 vccd1 vccd1 _09910_/B sky130_fd_sc_hd__and3_1
XFILLER_59_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout563 _17112_/A1 vssd1 vssd1 vccd1 vccd1 _13516_/S sky130_fd_sc_hd__clkbuf_4
Xfanout574 fanout578/X vssd1 vssd1 vccd1 vccd1 _15805_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_47_915 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout585 _15126_/A vssd1 vssd1 vccd1 vccd1 _10753_/A sky130_fd_sc_hd__buf_2
X_12920_ _12920_/A _12920_/B _12920_/C vssd1 vssd1 vccd1 vccd1 _12933_/A sky130_fd_sc_hd__and3_1
Xfanout596 _14982_/A vssd1 vssd1 vccd1 vccd1 _14954_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_101_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12851_ _12220_/X _12229_/C _17164_/B vssd1 vssd1 vccd1 vccd1 _12852_/B sky130_fd_sc_hd__mux2_1
XTAP_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_34 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11802_ _11837_/A _11802_/B vssd1 vssd1 vccd1 vccd1 _11802_/Y sky130_fd_sc_hd__nand2_1
XTAP_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15570_ _15570_/A _15570_/B vssd1 vssd1 vccd1 vccd1 _15573_/A sky130_fd_sc_hd__xor2_1
XTAP_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12782_ _12938_/A _12782_/B _12782_/C vssd1 vssd1 vccd1 vccd1 _12938_/B sky130_fd_sc_hd__nand3_2
XTAP_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14521_ _14463_/B _14465_/A _14519_/X _14520_/Y vssd1 vssd1 vccd1 vccd1 _14577_/A
+ sky130_fd_sc_hd__a211o_1
XTAP_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11733_ _11732_/B _11732_/C _11732_/A vssd1 vssd1 vccd1 vccd1 _11733_/X sky130_fd_sc_hd__o21a_1
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17240_ _17589_/Q _17273_/A2 _17273_/B1 vssd1 vssd1 vccd1 vccd1 _17240_/X sky130_fd_sc_hd__a21o_1
XFILLER_30_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14452_ _14387_/A _14450_/B _14388_/A _14386_/B vssd1 vssd1 vccd1 vccd1 _14454_/B
+ sky130_fd_sc_hd__a31o_1
X_11664_ _11664_/A _11664_/B vssd1 vssd1 vccd1 vccd1 _11673_/B sky130_fd_sc_hd__nor2_1
XFILLER_168_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13403_ _13403_/A _13403_/B vssd1 vssd1 vccd1 vccd1 _13409_/A sky130_fd_sc_hd__nand2_1
X_10615_ _10615_/A _10615_/B _10615_/C vssd1 vssd1 vccd1 vccd1 _10615_/Y sky130_fd_sc_hd__nand3_1
X_17171_ input69/X input68/X input35/X vssd1 vssd1 vccd1 vccd1 _17171_/X sky130_fd_sc_hd__and3b_2
X_14383_ _14383_/A _14383_/B vssd1 vssd1 vccd1 vccd1 _14509_/A sky130_fd_sc_hd__and2_1
X_11595_ _11595_/A _11595_/B vssd1 vssd1 vccd1 vccd1 _11628_/B sky130_fd_sc_hd__xnor2_1
XFILLER_10_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16122_ _16122_/A _16122_/B _16122_/C vssd1 vssd1 vccd1 vccd1 _16122_/X sky130_fd_sc_hd__and3_1
X_13334_ _14769_/A _13450_/B _13334_/C _13966_/D vssd1 vssd1 vccd1 vccd1 _13455_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_128_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10546_ _10546_/A _10655_/A vssd1 vssd1 vccd1 vccd1 _10547_/C sky130_fd_sc_hd__nor2_1
XFILLER_6_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_577 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_565 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16053_ _16935_/A _16054_/B vssd1 vssd1 vccd1 vccd1 _16695_/B sky130_fd_sc_hd__and2_2
XFILLER_142_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_983 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13265_ _13266_/A _13266_/B vssd1 vssd1 vccd1 vccd1 _13509_/A sky130_fd_sc_hd__or2_1
X_10477_ _10591_/A _11027_/A _10594_/B _11006_/C vssd1 vssd1 vccd1 vccd1 _10478_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_6_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15004_ _15002_/X _15003_/X _14941_/X vssd1 vssd1 vccd1 vccd1 _15004_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_170_558 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12216_ _12216_/A vssd1 vssd1 vccd1 vccd1 _12217_/B sky130_fd_sc_hd__inv_2
XFILLER_155_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13196_ _14215_/A _13434_/D vssd1 vssd1 vccd1 vccd1 _13197_/B sky130_fd_sc_hd__nand2_1
XFILLER_29_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_997 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12147_ _12148_/A _12148_/B _12148_/C vssd1 vssd1 vccd1 vccd1 _12149_/A sky130_fd_sc_hd__a21oi_1
XFILLER_173_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16955_ _16955_/A _16955_/B vssd1 vssd1 vccd1 vccd1 _16958_/A sky130_fd_sc_hd__xnor2_1
X_12078_ _12078_/A _12078_/B vssd1 vssd1 vccd1 vccd1 _12080_/A sky130_fd_sc_hd__nor2_1
XFILLER_110_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_168 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11029_ _11032_/A _11029_/B _11025_/Y vssd1 vssd1 vccd1 vccd1 _11046_/A sky130_fd_sc_hd__or3b_1
X_15906_ _16207_/B _15889_/Y _15894_/X _15905_/X vssd1 vssd1 vccd1 vccd1 _15906_/X
+ sky130_fd_sc_hd__o211a_1
X_16886_ _16886_/A _16886_/B vssd1 vssd1 vccd1 vccd1 _16887_/B sky130_fd_sc_hd__and2_1
XFILLER_38_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15837_ _15837_/A _15837_/B vssd1 vssd1 vccd1 vccd1 _15841_/A sky130_fd_sc_hd__xnor2_2
XFILLER_65_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15768_ _15769_/A _15769_/B _15769_/C vssd1 vssd1 vccd1 vccd1 _15877_/A sky130_fd_sc_hd__o21a_1
XTAP_3490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_642 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17507_ fanout945/X _17507_/D vssd1 vssd1 vccd1 vccd1 _17507_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14719_ _14719_/A _14719_/B _14719_/C vssd1 vssd1 vccd1 vccd1 _14747_/B sky130_fd_sc_hd__or3_1
XFILLER_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_973 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15699_ _15610_/Y _15611_/X _15610_/A vssd1 vssd1 vccd1 vccd1 _15700_/B sky130_fd_sc_hd__a21oi_1
XFILLER_32_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17438_ fanout939/X _17438_/D vssd1 vssd1 vccd1 vccd1 _17438_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_123_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_15 _16641_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_336 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_26 _17536_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_37 _08988_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_48 _12442_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17369_ _17369_/A _17377_/B vssd1 vssd1 vccd1 vccd1 _17369_/Y sky130_fd_sc_hd__nand2_1
XANTENNA_59 _10146_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_363 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput100 _17458_/Q vssd1 vssd1 vccd1 vccd1 o_wb_data[24] sky130_fd_sc_hd__clkbuf_1
XFILLER_161_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput111 _17439_/Q vssd1 vssd1 vccd1 vccd1 o_wb_data[5] sky130_fd_sc_hd__clkbuf_1
XFILLER_115_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09625_ _09627_/A _09625_/B vssd1 vssd1 vccd1 vccd1 _09626_/C sky130_fd_sc_hd__nor2_1
XFILLER_102_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09556_ _09556_/A _09556_/B vssd1 vssd1 vccd1 vccd1 _09558_/A sky130_fd_sc_hd__nor2_1
XFILLER_71_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09487_ _09460_/X _09484_/B _09486_/Y _09388_/A vssd1 vssd1 vccd1 vccd1 _09487_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_23_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10400_ _10501_/A _10501_/B _10396_/X vssd1 vssd1 vccd1 vccd1 _10402_/C sky130_fd_sc_hd__a21o_1
XFILLER_165_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11380_ _11380_/A _11380_/B _11380_/C vssd1 vssd1 vccd1 vccd1 _11426_/A sky130_fd_sc_hd__or3_1
XFILLER_164_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10331_ _10331_/A _10331_/B vssd1 vssd1 vccd1 vccd1 _10333_/B sky130_fd_sc_hd__xor2_1
XFILLER_139_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_780 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1038 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13050_ _13051_/B _13948_/C _13051_/D _13182_/A vssd1 vssd1 vccd1 vccd1 _13052_/A
+ sky130_fd_sc_hd__a22oi_1
X_10262_ _10262_/A _10262_/B _10262_/C vssd1 vssd1 vccd1 vccd1 _10262_/X sky130_fd_sc_hd__and3_1
XFILLER_140_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12001_ _11998_/X _11999_/Y _09122_/A _09255_/X vssd1 vssd1 vccd1 vccd1 _12001_/Y
+ sky130_fd_sc_hd__a211oi_1
XFILLER_79_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_34 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10193_ _10193_/A _10193_/B vssd1 vssd1 vccd1 vccd1 _10194_/C sky130_fd_sc_hd__nor2_1
XFILLER_160_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_848 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout360 _17536_/Q vssd1 vssd1 vccd1 vccd1 _16965_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_120_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout371 _17535_/Q vssd1 vssd1 vccd1 vccd1 _12487_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_59_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout382 _13689_/A vssd1 vssd1 vccd1 vccd1 _14387_/A sky130_fd_sc_hd__buf_2
X_16740_ _16722_/A _16806_/A2 _16719_/Y _16739_/X vssd1 vssd1 vccd1 vccd1 _17565_/D
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_19_414 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13952_ _13954_/A _13954_/B _13954_/C vssd1 vssd1 vccd1 vccd1 _14044_/A sky130_fd_sc_hd__o21a_1
Xfanout393 _14772_/A vssd1 vssd1 vccd1 vccd1 _10560_/A sky130_fd_sc_hd__buf_2
XFILLER_120_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1022 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12903_ _12903_/A _12903_/B vssd1 vssd1 vccd1 vccd1 _12913_/A sky130_fd_sc_hd__or2_1
X_16671_ _16671_/A _16671_/B vssd1 vssd1 vccd1 vccd1 _16673_/B sky130_fd_sc_hd__nor2_1
XFILLER_100_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13883_ _13774_/A _13776_/B _13774_/B vssd1 vssd1 vccd1 vccd1 _13885_/B sky130_fd_sc_hd__o21ba_1
XFILLER_28_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15622_ _15622_/A _15622_/B vssd1 vssd1 vccd1 vccd1 _15623_/B sky130_fd_sc_hd__nand2_1
X_12834_ _12991_/B _12834_/B _12834_/C vssd1 vssd1 vccd1 vccd1 _13001_/A sky130_fd_sc_hd__or3_1
XTAP_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15553_ _15553_/A _15553_/B _16514_/A vssd1 vssd1 vccd1 vccd1 _15555_/B sky130_fd_sc_hd__or3_1
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12765_ _12928_/B _12766_/C _12766_/A vssd1 vssd1 vccd1 vccd1 _12765_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_15_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14504_ _14505_/A _14505_/B vssd1 vssd1 vccd1 vccd1 _14565_/A sky130_fd_sc_hd__nor2_1
X_11716_ _11302_/B _16294_/A _11302_/A vssd1 vssd1 vccd1 vccd1 _16387_/C sky130_fd_sc_hd__o21a_1
XTAP_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15484_ _15484_/A _15567_/A vssd1 vssd1 vccd1 vccd1 _15486_/A sky130_fd_sc_hd__xnor2_1
XTAP_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12696_ _12696_/A _12696_/B vssd1 vssd1 vccd1 vccd1 _13004_/A sky130_fd_sc_hd__or2_1
XFILLER_30_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17223_ _17551_/Q _17274_/B vssd1 vssd1 vccd1 vccd1 _17223_/X sky130_fd_sc_hd__and2_1
XFILLER_174_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14435_ _17023_/A _14492_/A _14432_/X vssd1 vssd1 vccd1 vccd1 _14437_/C sky130_fd_sc_hd__o21a_1
X_11647_ _11624_/A _11624_/B _15524_/B _15524_/C vssd1 vssd1 vccd1 vccd1 _15525_/A
+ sky130_fd_sc_hd__a22o_1
Xinput13 i_wb_addr[19] vssd1 vssd1 vccd1 vccd1 input13/X sky130_fd_sc_hd__clkbuf_1
XFILLER_128_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput24 i_wb_addr[29] vssd1 vssd1 vccd1 vccd1 input24/X sky130_fd_sc_hd__clkbuf_1
X_17154_ _17133_/A _17136_/X _17152_/Y _17153_/X vssd1 vssd1 vccd1 vccd1 _17154_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_155_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput35 i_wb_cyc vssd1 vssd1 vccd1 vccd1 input35/X sky130_fd_sc_hd__clkbuf_2
X_14366_ _14599_/B _14366_/B vssd1 vssd1 vccd1 vccd1 _17023_/A sky130_fd_sc_hd__nand2_4
X_11578_ _11574_/A _11574_/C _11607_/A vssd1 vssd1 vccd1 vccd1 _11579_/C sky130_fd_sc_hd__o21ai_1
Xinput46 i_wb_data[19] vssd1 vssd1 vccd1 vccd1 input46/X sky130_fd_sc_hd__clkbuf_1
XFILLER_156_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput57 i_wb_data[29] vssd1 vssd1 vccd1 vccd1 input57/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_156_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16105_ _16105_/A _16105_/B vssd1 vssd1 vccd1 vccd1 _16106_/B sky130_fd_sc_hd__xor2_2
XFILLER_143_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput68 i_wb_stb vssd1 vssd1 vccd1 vccd1 input68/X sky130_fd_sc_hd__clkbuf_2
XFILLER_156_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13317_ _13317_/A _13317_/B _13317_/C vssd1 vssd1 vccd1 vccd1 _13431_/B sky130_fd_sc_hd__and3_1
X_10529_ _15805_/A _10421_/D _10422_/A _10420_/Y vssd1 vssd1 vccd1 vccd1 _10531_/C
+ sky130_fd_sc_hd__o2bb2a_1
X_17085_ _17085_/A _17085_/B _17085_/C vssd1 vssd1 vccd1 vccd1 _17086_/B sky130_fd_sc_hd__or3_1
X_14297_ _14297_/A _14297_/B vssd1 vssd1 vccd1 vccd1 _14337_/A sky130_fd_sc_hd__xor2_1
XFILLER_143_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16036_ _16036_/A _16036_/B vssd1 vssd1 vccd1 vccd1 _16048_/A sky130_fd_sc_hd__xnor2_1
X_13248_ _13248_/A _13248_/B _13248_/C vssd1 vssd1 vccd1 vccd1 _13249_/D sky130_fd_sc_hd__or3_1
XFILLER_112_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13179_ _13046_/A _13047_/B _13177_/Y _13312_/B vssd1 vssd1 vccd1 vccd1 _13189_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16938_ _16938_/A _16938_/B _16939_/B _16938_/D vssd1 vssd1 vccd1 vccd1 _16994_/A
+ sky130_fd_sc_hd__or4_1
XFILLER_37_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16869_ _16864_/B _17162_/A2 _16974_/B _14864_/A _16869_/C1 vssd1 vssd1 vccd1 vccd1
+ _16869_/X sky130_fd_sc_hd__a221o_1
XFILLER_25_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09410_ _09410_/A _09548_/A vssd1 vssd1 vccd1 vccd1 _09417_/B sky130_fd_sc_hd__nor2_1
XFILLER_53_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09341_ _09214_/A _09214_/B _09214_/C vssd1 vssd1 vccd1 vccd1 _09342_/B sky130_fd_sc_hd__a21oi_1
XFILLER_33_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09272_ _09414_/A _12077_/B _11961_/B _09272_/D vssd1 vssd1 vccd1 vccd1 _09273_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_61_792 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_280 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_820 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_875 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_823 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08987_ _12770_/B _11920_/D _09362_/D _17425_/A vssd1 vssd1 vccd1 vccd1 _08989_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_103_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_786 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09608_ _15538_/A _14864_/A _09602_/A _09471_/Y vssd1 vssd1 vccd1 vccd1 _09610_/C
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_113_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_523 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10880_ _11114_/A _11114_/B vssd1 vssd1 vccd1 vccd1 _10883_/C sky130_fd_sc_hd__nand2_1
XFILLER_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09539_ _09531_/X _09532_/Y _09487_/X _09530_/B vssd1 vssd1 vccd1 vccd1 _09540_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_25_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_910 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12550_ _12545_/X _12549_/X _17371_/A vssd1 vssd1 vccd1 vccd1 _12550_/X sky130_fd_sc_hd__mux2_1
XFILLER_12_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11501_ _11456_/X _11490_/Y _11499_/A _11539_/A vssd1 vssd1 vccd1 vccd1 _11502_/C
+ sky130_fd_sc_hd__a211oi_1
XFILLER_11_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12481_ _12481_/A _12481_/B _12481_/C vssd1 vssd1 vccd1 vccd1 _12481_/Y sky130_fd_sc_hd__nand3_1
XFILLER_12_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14220_ _14221_/A _14221_/B _14221_/C vssd1 vssd1 vccd1 vccd1 _14222_/A sky130_fd_sc_hd__o21ai_1
X_11432_ _11426_/A _11426_/C _11426_/B vssd1 vssd1 vccd1 vccd1 _11433_/C sky130_fd_sc_hd__a21o_1
XFILLER_156_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_188 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_51 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14151_ _14151_/A _14151_/B vssd1 vssd1 vccd1 vccd1 _14190_/A sky130_fd_sc_hd__nor2_1
X_11363_ _11492_/A _11492_/B vssd1 vssd1 vccd1 vccd1 _11447_/A sky130_fd_sc_hd__nand2b_1
X_13102_ _13103_/A _13103_/B vssd1 vssd1 vccd1 vccd1 _13236_/A sky130_fd_sc_hd__and2b_1
X_10314_ _10314_/A _10314_/B vssd1 vssd1 vccd1 vccd1 _10315_/C sky130_fd_sc_hd__xnor2_1
XFILLER_125_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14082_ _14387_/A _14366_/B vssd1 vssd1 vccd1 vccd1 _14084_/B sky130_fd_sc_hd__nand2_1
X_11294_ _11299_/A _11294_/B vssd1 vssd1 vccd1 vccd1 _11345_/A sky130_fd_sc_hd__nand2_1
XFILLER_4_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13033_ _13033_/A _13033_/B _13033_/C vssd1 vssd1 vccd1 vccd1 _13046_/B sky130_fd_sc_hd__nand3_1
XFILLER_79_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10245_ _10245_/A _10245_/B vssd1 vssd1 vccd1 vccd1 _10358_/A sky130_fd_sc_hd__xnor2_1
XFILLER_78_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10176_ _10177_/B _10289_/A _10177_/A vssd1 vssd1 vccd1 vccd1 _10188_/A sky130_fd_sc_hd__a21o_1
XFILLER_154_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14984_ _15252_/B _14983_/X _15384_/S vssd1 vssd1 vccd1 vccd1 _15537_/B sky130_fd_sc_hd__mux2_1
XFILLER_120_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout190 _16138_/A vssd1 vssd1 vccd1 vccd1 _16410_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_19_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13935_ _13935_/A _13935_/B _13510_/X vssd1 vssd1 vccd1 vccd1 _13935_/Y sky130_fd_sc_hd__nor3b_1
X_16723_ _16723_/A _16723_/B vssd1 vssd1 vccd1 vccd1 _16723_/Y sky130_fd_sc_hd__nand2_1
XFILLER_93_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16654_ _16649_/B _17162_/A2 _16974_/B _16654_/B2 _17162_/C1 vssd1 vssd1 vccd1 vccd1
+ _16654_/X sky130_fd_sc_hd__a221o_1
XFILLER_19_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13866_ _13966_/A _14213_/B _13866_/C _13866_/D vssd1 vssd1 vccd1 vccd1 _13867_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_16_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15605_ _15507_/A _15507_/B _15509_/Y vssd1 vssd1 vccd1 vccd1 _15607_/B sky130_fd_sc_hd__a21o_1
X_12817_ _12817_/A _12817_/B vssd1 vssd1 vccd1 vccd1 _12820_/C sky130_fd_sc_hd__xnor2_1
X_16585_ _16566_/Y _16567_/X _16579_/X _16584_/X vssd1 vssd1 vccd1 vccd1 _16585_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_50_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13797_ _14176_/A _13993_/B _13796_/C vssd1 vssd1 vccd1 vccd1 _13798_/B sky130_fd_sc_hd__a21o_1
XFILLER_62_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_1014 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15536_ _10716_/A _14785_/X _14806_/X _15535_/Y vssd1 vssd1 vccd1 vccd1 _15536_/X
+ sky130_fd_sc_hd__a31o_1
X_12748_ _13051_/B _13037_/B _13035_/C _13182_/A vssd1 vssd1 vccd1 vccd1 _12751_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_31_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15467_ _15454_/X _15467_/B _15467_/C _15467_/D vssd1 vssd1 vccd1 vccd1 _15467_/X
+ sky130_fd_sc_hd__and4b_1
XFILLER_129_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12679_ _12679_/A _12679_/B vssd1 vssd1 vccd1 vccd1 _12682_/A sky130_fd_sc_hd__nand2_1
XFILLER_8_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17206_ _17436_/Q _17275_/A2 _17204_/X _17205_/X _17364_/C1 vssd1 vssd1 vccd1 vccd1
+ _17436_/D sky130_fd_sc_hd__o221a_1
XFILLER_147_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14418_ _14533_/A _14419_/B vssd1 vssd1 vccd1 vccd1 _14418_/X sky130_fd_sc_hd__or2_1
XFILLER_129_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15398_ _15913_/A _15832_/A vssd1 vssd1 vccd1 vccd1 _15481_/A sky130_fd_sc_hd__nor2_1
XFILLER_8_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17137_ _17167_/A _14829_/X _14828_/Y _14597_/B vssd1 vssd1 vccd1 vccd1 _17137_/X
+ sky130_fd_sc_hd__a211o_1
X_14349_ _14350_/A _14350_/B _14350_/C vssd1 vssd1 vccd1 vccd1 _14349_/X sky130_fd_sc_hd__o21a_1
XFILLER_144_834 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17068_ _17064_/X _17065_/X _17066_/X _17018_/Y vssd1 vssd1 vccd1 vccd1 _17068_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_170_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08910_ _08910_/A _08910_/B _08910_/C vssd1 vssd1 vccd1 vccd1 _08910_/Y sky130_fd_sc_hd__nand3_1
X_16019_ _16019_/A vssd1 vssd1 vccd1 vccd1 _17557_/D sky130_fd_sc_hd__clkinv_2
XFILLER_98_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09890_ _09890_/A _09898_/A _09890_/C vssd1 vssd1 vccd1 vccd1 _09891_/B sky130_fd_sc_hd__or3_1
XFILLER_112_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08841_ _17383_/A _09319_/C _09319_/D _08913_/A vssd1 vssd1 vccd1 vccd1 _08841_/Y
+ sky130_fd_sc_hd__a22oi_1
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_998 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_786 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08772_ _17401_/A _09229_/B _08772_/C _08772_/D vssd1 vssd1 vccd1 vccd1 _08804_/A
+ sky130_fd_sc_hd__and4_1
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_386 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09324_ _09328_/A _09451_/A _09328_/C vssd1 vssd1 vccd1 vccd1 _09332_/B sky130_fd_sc_hd__o21ai_1
XFILLER_34_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09255_ _09256_/A _09255_/B _09255_/C vssd1 vssd1 vccd1 vccd1 _09255_/X sky130_fd_sc_hd__and3_1
XFILLER_21_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09186_ _17535_/Q _17411_/A _09267_/D _12174_/D vssd1 vssd1 vccd1 vccd1 _09221_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_88_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10030_ _09909_/A _09909_/B _09909_/C vssd1 vssd1 vccd1 vccd1 _10030_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_89_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11981_ _11982_/A _11982_/B vssd1 vssd1 vccd1 vccd1 _12183_/A sky130_fd_sc_hd__and2b_1
XFILLER_75_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13720_ _13720_/A _13720_/B vssd1 vssd1 vccd1 vccd1 _13723_/A sky130_fd_sc_hd__xnor2_1
XFILLER_84_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10932_ _11124_/C _10932_/B vssd1 vssd1 vccd1 vccd1 _10936_/A sky130_fd_sc_hd__nand2_1
XFILLER_44_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13651_ _13643_/A _13844_/C _13534_/A _13532_/B vssd1 vssd1 vccd1 vccd1 _13652_/B
+ sky130_fd_sc_hd__a31o_1
X_10863_ _10863_/A _10863_/B _10863_/C vssd1 vssd1 vccd1 vccd1 _10895_/A sky130_fd_sc_hd__or3_1
XFILLER_44_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12602_ _12603_/B _12603_/A vssd1 vssd1 vccd1 vccd1 _12764_/A sky130_fd_sc_hd__nand2b_1
XPHY_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16370_ _16272_/A _16271_/B _16271_/A vssd1 vssd1 vccd1 vccd1 _16372_/B sky130_fd_sc_hd__o21ba_1
XFILLER_13_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13582_ _13582_/A _13582_/B vssd1 vssd1 vccd1 vccd1 _13584_/A sky130_fd_sc_hd__nor2_1
X_10794_ _10794_/A _10794_/B vssd1 vssd1 vccd1 vccd1 _10884_/B sky130_fd_sc_hd__nor2_1
XPHY_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15321_ _15321_/A _15321_/B _15321_/C _15321_/D vssd1 vssd1 vccd1 vccd1 _15321_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_169_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12533_ _12534_/B _12534_/A vssd1 vssd1 vccd1 vccd1 _12533_/X sky130_fd_sc_hd__and2b_1
XPHY_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15252_ _16011_/B _15252_/B vssd1 vssd1 vccd1 vccd1 _15252_/X sky130_fd_sc_hd__or2_1
X_12464_ _12464_/A _12662_/A vssd1 vssd1 vccd1 vccd1 _12467_/A sky130_fd_sc_hd__or2_1
XFILLER_32_1042 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_94 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14203_ _14202_/A _14202_/B _14202_/C vssd1 vssd1 vccd1 vccd1 _14279_/B sky130_fd_sc_hd__a21oi_1
X_11415_ _11415_/A _11415_/B vssd1 vssd1 vccd1 vccd1 _11418_/A sky130_fd_sc_hd__nand2_1
X_15183_ _11321_/X _14790_/Y _14798_/Y _16485_/A _15182_/Y vssd1 vssd1 vccd1 vccd1
+ _15188_/A sky130_fd_sc_hd__o311a_1
X_12395_ _12391_/X _12394_/Y _13840_/S vssd1 vssd1 vccd1 vccd1 _14210_/A sky130_fd_sc_hd__mux2_1
XFILLER_137_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14134_ _14134_/A _14134_/B _14134_/C vssd1 vssd1 vccd1 vccd1 _14218_/B sky130_fd_sc_hd__nor3_1
X_11346_ _11343_/A _11312_/Y _11329_/Y _11367_/A vssd1 vssd1 vccd1 vccd1 _11349_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_152_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14065_ _14155_/A _14065_/B vssd1 vssd1 vccd1 vccd1 _14066_/B sky130_fd_sc_hd__nand2_1
XFILLER_165_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11277_ _11518_/B _15208_/A vssd1 vssd1 vccd1 vccd1 _11387_/C sky130_fd_sc_hd__and2_1
XFILLER_79_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13016_ _17371_/A _13831_/S _11820_/A _13015_/Y _15457_/A vssd1 vssd1 vccd1 vccd1
+ _13016_/X sky130_fd_sc_hd__a311o_1
XFILLER_79_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10228_ _10214_/A _10214_/C _10214_/B vssd1 vssd1 vccd1 vccd1 _10228_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_121_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10159_ _10053_/A _10053_/B _10053_/C vssd1 vssd1 vccd1 vccd1 _10159_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_94_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14967_ _15617_/A _15208_/A _14967_/C _14967_/D vssd1 vssd1 vccd1 vccd1 _14967_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_54_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16706_ _16784_/A _16706_/B vssd1 vssd1 vccd1 vccd1 _16709_/A sky130_fd_sc_hd__and2_1
XFILLER_63_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13918_ _13918_/A _13918_/B vssd1 vssd1 vccd1 vccd1 _13919_/B sky130_fd_sc_hd__or2_1
X_14898_ _14899_/C vssd1 vssd1 vccd1 vccd1 _14898_/Y sky130_fd_sc_hd__inv_2
XFILLER_74_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16637_ _16714_/A _16637_/B vssd1 vssd1 vccd1 vccd1 _16638_/B sky130_fd_sc_hd__or2_1
X_13849_ _13849_/A _13849_/B _13849_/C vssd1 vssd1 vccd1 vccd1 _13851_/A sky130_fd_sc_hd__nor3_1
XFILLER_35_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16568_ _16568_/A _16568_/B vssd1 vssd1 vccd1 vccd1 _16568_/Y sky130_fd_sc_hd__nor2_1
XFILLER_31_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15519_ _15520_/A _15520_/B _15520_/C vssd1 vssd1 vccd1 vccd1 _15519_/X sky130_fd_sc_hd__o21a_1
X_16499_ _16747_/A _16499_/B _16499_/C vssd1 vssd1 vccd1 vccd1 _16609_/B sky130_fd_sc_hd__or3_1
XFILLER_148_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09040_ _14873_/B _10647_/D vssd1 vssd1 vccd1 vccd1 _17081_/B sky130_fd_sc_hd__nand2_4
XFILLER_30_283 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmax_cap121 _11586_/B vssd1 vssd1 vccd1 vccd1 _11620_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_144_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09942_ _09942_/A _10062_/B _10062_/C vssd1 vssd1 vccd1 vccd1 _09945_/A sky130_fd_sc_hd__and3_1
Xfanout904 _17479_/Q vssd1 vssd1 vccd1 vccd1 fanout904/X sky130_fd_sc_hd__clkbuf_4
Xfanout915 _17225_/B1 vssd1 vssd1 vccd1 vccd1 _17273_/B1 sky130_fd_sc_hd__clkbuf_4
Xfanout926 _17358_/C1 vssd1 vssd1 vccd1 vccd1 _17426_/C1 sky130_fd_sc_hd__buf_2
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout937 fanout941/X vssd1 vssd1 vccd1 vccd1 fanout937/X sky130_fd_sc_hd__clkbuf_2
X_09873_ _09873_/A _14784_/A _10016_/D _10146_/B vssd1 vssd1 vccd1 vccd1 _09876_/A
+ sky130_fd_sc_hd__and4_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout948 fanout957/X vssd1 vssd1 vccd1 vccd1 fanout948/X sky130_fd_sc_hd__clkbuf_2
XFILLER_100_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08824_ _17387_/A _09058_/C vssd1 vssd1 vccd1 vccd1 _08893_/A sky130_fd_sc_hd__nand2_1
XFILLER_58_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_946 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08755_ _08755_/A _08768_/A vssd1 vssd1 vccd1 vccd1 _08757_/B sky130_fd_sc_hd__nor2_2
XFILLER_57_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_1012 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09307_ _09438_/A _09438_/B vssd1 vssd1 vccd1 vccd1 _09439_/A sky130_fd_sc_hd__and2_1
XFILLER_16_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_907 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09238_ _09238_/A _09238_/B _09238_/C vssd1 vssd1 vccd1 vccd1 _09239_/B sky130_fd_sc_hd__nor3_1
XFILLER_139_469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09169_ _09333_/A _09333_/B vssd1 vssd1 vccd1 vccd1 _09178_/B sky130_fd_sc_hd__nand2b_1
XFILLER_108_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11200_ _11201_/A _11201_/B vssd1 vssd1 vccd1 vccd1 _11200_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_135_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12180_ _12180_/A _12180_/B vssd1 vssd1 vccd1 vccd1 _12182_/A sky130_fd_sc_hd__nor2_1
XFILLER_79_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11131_ _11131_/A _11131_/B vssd1 vssd1 vccd1 vccd1 _11137_/A sky130_fd_sc_hd__xnor2_1
XFILLER_1_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11062_ _10951_/A _10949_/Y _10857_/Y _10863_/B vssd1 vssd1 vccd1 vccd1 _11065_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_49_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10013_ _14784_/A _10014_/D vssd1 vssd1 vccd1 vccd1 _10145_/A sky130_fd_sc_hd__nand2_1
X_15870_ _15868_/A _15868_/B _15871_/B vssd1 vssd1 vccd1 vccd1 _15989_/A sky130_fd_sc_hd__o21ba_1
XFILLER_95_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_391 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14821_ _16796_/B _16797_/A _16796_/A vssd1 vssd1 vccd1 vccd1 _16865_/A sky130_fd_sc_hd__a21bo_1
XFILLER_36_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_62 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17540_ fanout944/X _17540_/D vssd1 vssd1 vccd1 vccd1 _17540_/Q sky130_fd_sc_hd__dfxtp_1
X_14752_ _14729_/A _14726_/X _14728_/B vssd1 vssd1 vccd1 vccd1 _14752_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_17_534 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11964_ _17407_/A _09557_/B _09225_/A _09223_/B vssd1 vssd1 vccd1 vccd1 _11965_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_91_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13703_ _13703_/A _13703_/B vssd1 vssd1 vccd1 vccd1 _13705_/A sky130_fd_sc_hd__nor2_1
X_17471_ fanout955/X _17544_/Q vssd1 vssd1 vccd1 vccd1 _17471_/Q sky130_fd_sc_hd__dfxtp_1
X_10915_ _10915_/A _10915_/B vssd1 vssd1 vccd1 vccd1 _10918_/A sky130_fd_sc_hd__xnor2_1
XFILLER_60_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14683_ _14683_/A _14693_/B vssd1 vssd1 vccd1 vccd1 _14684_/A sky130_fd_sc_hd__and2_1
X_11895_ _17379_/A _11895_/B _11895_/C _11895_/D vssd1 vssd1 vccd1 vccd1 _12138_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_32_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16422_ _16422_/A _16422_/B vssd1 vssd1 vccd1 vccd1 _16509_/B sky130_fd_sc_hd__nand2_1
X_13634_ _13635_/A _13741_/A _13635_/C vssd1 vssd1 vccd1 vccd1 _13741_/B sky130_fd_sc_hd__nor3_1
X_10846_ _10846_/A _10846_/B vssd1 vssd1 vccd1 vccd1 _10859_/A sky130_fd_sc_hd__xnor2_1
XFILLER_158_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16353_ _16619_/A _15658_/Y _16681_/C _16446_/A vssd1 vssd1 vccd1 vccd1 _16354_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_13_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13565_ _13565_/A _13695_/A vssd1 vssd1 vccd1 vccd1 _13568_/A sky130_fd_sc_hd__nor2_1
X_10777_ _10777_/A _10778_/A _10777_/C vssd1 vssd1 vccd1 vccd1 _11742_/A sky130_fd_sc_hd__nor3_1
XFILLER_12_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15304_ _15305_/C _15373_/B _15314_/A vssd1 vssd1 vccd1 vccd1 _15307_/A sky130_fd_sc_hd__a21boi_1
X_12516_ _12517_/A _12517_/B vssd1 vssd1 vccd1 vccd1 _12516_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_157_255 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16284_ _16192_/A _16192_/B _16184_/A vssd1 vssd1 vccd1 vccd1 _16285_/B sky130_fd_sc_hd__a21o_1
XFILLER_8_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13496_ _13496_/A _13496_/B vssd1 vssd1 vccd1 vccd1 _13498_/B sky130_fd_sc_hd__nor2_1
XFILLER_173_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15235_ _15235_/A _15235_/B _15235_/C vssd1 vssd1 vccd1 vccd1 _15235_/Y sky130_fd_sc_hd__nand3_1
XFILLER_8_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12447_ _12907_/A _12447_/B vssd1 vssd1 vccd1 vccd1 _12448_/B sky130_fd_sc_hd__nand2_1
XFILLER_126_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15166_ _15166_/A _15166_/B vssd1 vssd1 vccd1 vccd1 _15169_/A sky130_fd_sc_hd__xnor2_1
X_12378_ _11781_/B _12377_/Y _13005_/A vssd1 vssd1 vccd1 vccd1 _12379_/B sky130_fd_sc_hd__a21oi_1
XFILLER_99_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14117_ _14117_/A _14117_/B vssd1 vssd1 vccd1 vccd1 _14117_/X sky130_fd_sc_hd__xor2_1
XFILLER_99_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11329_ _11331_/B _11331_/C _11331_/A vssd1 vssd1 vccd1 vccd1 _11329_/Y sky130_fd_sc_hd__a21oi_1
X_15097_ _15097_/A _15097_/B vssd1 vssd1 vccd1 vccd1 _15097_/X sky130_fd_sc_hd__or2_1
XFILLER_99_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14048_ _14150_/A _14048_/B vssd1 vssd1 vccd1 vccd1 _14057_/A sky130_fd_sc_hd__or2_1
XFILLER_79_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15999_ _16317_/A _16644_/B _16014_/A vssd1 vssd1 vccd1 vccd1 _16001_/A sky130_fd_sc_hd__a21bo_1
XFILLER_35_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_592 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09023_ _12068_/A _12068_/B _12340_/B _09267_/D vssd1 vssd1 vccd1 vccd1 _09026_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_40_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout701 _16654_/B2 vssd1 vssd1 vccd1 vccd1 _13564_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_172_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout712 _17498_/Q vssd1 vssd1 vccd1 vccd1 _16571_/A sky130_fd_sc_hd__clkbuf_4
X_09925_ _09925_/A _14863_/B vssd1 vssd1 vccd1 vccd1 _09926_/C sky130_fd_sc_hd__and2_1
Xfanout723 _10657_/B vssd1 vssd1 vccd1 vccd1 _10545_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_131_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_829 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout734 _16298_/A vssd1 vssd1 vccd1 vccd1 _13080_/C sky130_fd_sc_hd__clkbuf_2
Xfanout745 _10297_/D vssd1 vssd1 vccd1 vccd1 _12500_/B sky130_fd_sc_hd__buf_4
Xfanout756 _16114_/A vssd1 vssd1 vccd1 vccd1 _17119_/A sky130_fd_sc_hd__buf_2
XFILLER_105_22 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout767 fanout772/X vssd1 vssd1 vccd1 vccd1 _16014_/A sky130_fd_sc_hd__buf_2
X_09856_ _10254_/A _10270_/B vssd1 vssd1 vccd1 vccd1 _09856_/Y sky130_fd_sc_hd__nand2_1
Xfanout778 _10743_/C vssd1 vssd1 vccd1 vccd1 _16758_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout789 _11132_/C vssd1 vssd1 vccd1 vccd1 _16745_/A sky130_fd_sc_hd__clkbuf_2
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08807_ _08808_/A _08806_/Y _17401_/A _09272_/D vssd1 vssd1 vccd1 vccd1 _08883_/A
+ sky130_fd_sc_hd__and4bb_1
XTAP_3105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09787_ _09932_/A _09932_/B vssd1 vssd1 vccd1 vccd1 _09933_/A sky130_fd_sc_hd__or2_1
XTAP_3127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_88 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08738_ _17614_/Q _08737_/Y _17131_/A vssd1 vssd1 vccd1 vccd1 _17614_/D sky130_fd_sc_hd__mux2_1
XTAP_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10700_ _10701_/A _10701_/B vssd1 vssd1 vccd1 vccd1 _10715_/A sky130_fd_sc_hd__nand2_1
XTAP_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11680_ _11681_/A _11681_/B vssd1 vssd1 vccd1 vccd1 _11680_/Y sky130_fd_sc_hd__nor2_1
XTAP_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10631_ _10632_/A _10632_/B _10632_/C _10632_/D vssd1 vssd1 vccd1 vccd1 _10631_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_139_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13350_ _13195_/A _13197_/B _13195_/B vssd1 vssd1 vccd1 vccd1 _13357_/A sky130_fd_sc_hd__o21ba_1
XFILLER_14_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10562_ _10671_/A _10671_/B vssd1 vssd1 vccd1 vccd1 _10672_/A sky130_fd_sc_hd__or2_1
XFILLER_155_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12301_ _17375_/A _12439_/D _12105_/A _12103_/B vssd1 vssd1 vccd1 vccd1 _12303_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_154_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13281_ _13846_/A _14065_/B vssd1 vssd1 vccd1 vccd1 _13282_/B sky130_fd_sc_hd__nand2_1
X_10493_ _10493_/A _10493_/B vssd1 vssd1 vccd1 vccd1 _10601_/B sky130_fd_sc_hd__nor2_1
X_15020_ _15402_/A _15402_/B vssd1 vssd1 vccd1 vccd1 _15020_/X sky130_fd_sc_hd__and2_1
XFILLER_108_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12232_ _15998_/A _12210_/Y _12231_/X vssd1 vssd1 vccd1 vccd1 _17578_/D sky130_fd_sc_hd__o21ai_1
XFILLER_108_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12163_ _12163_/A _12163_/B _12163_/C vssd1 vssd1 vccd1 vccd1 _12165_/A sky130_fd_sc_hd__nor3_1
XFILLER_107_185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11114_ _11114_/A _11114_/B vssd1 vssd1 vccd1 vccd1 _11130_/A sky130_fd_sc_hd__xnor2_1
XFILLER_96_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12094_ _12286_/A _12094_/B vssd1 vssd1 vccd1 vccd1 _12096_/B sky130_fd_sc_hd__and2_1
X_16971_ _16971_/A _16971_/B vssd1 vssd1 vccd1 vccd1 _16971_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_7_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11045_ _11032_/A _11029_/B _11025_/Y vssd1 vssd1 vccd1 vccd1 _11046_/B sky130_fd_sc_hd__o21bai_1
X_15922_ _15923_/A _15923_/B vssd1 vssd1 vccd1 vccd1 _16036_/A sky130_fd_sc_hd__nor2_1
XFILLER_7_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15853_ _15853_/A _15853_/B vssd1 vssd1 vccd1 vccd1 _15855_/A sky130_fd_sc_hd__xnor2_1
XFILLER_92_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14804_ _14803_/A _14803_/B _10799_/Y vssd1 vssd1 vccd1 vccd1 _14805_/C sky130_fd_sc_hd__o21ai_1
XFILLER_36_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12996_ _12996_/A vssd1 vssd1 vccd1 vccd1 _12997_/C sky130_fd_sc_hd__inv_2
X_15784_ _15784_/A _15784_/B vssd1 vssd1 vccd1 vccd1 _15787_/B sky130_fd_sc_hd__nor2_1
XFILLER_29_191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17523_ fanout943/X _17523_/D vssd1 vssd1 vccd1 vccd1 _17523_/Q sky130_fd_sc_hd__dfxtp_4
X_11947_ _11917_/X _11918_/Y _12156_/B _11947_/D vssd1 vssd1 vccd1 vccd1 _11947_/X
+ sky130_fd_sc_hd__and4bb_1
XFILLER_33_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14735_ _14735_/A1 _13628_/B _13625_/Y _12853_/X vssd1 vssd1 vccd1 vccd1 _14735_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_18_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14666_ _13390_/X _13393_/B _14757_/S vssd1 vssd1 vccd1 vccd1 _14667_/B sky130_fd_sc_hd__mux2_1
X_17454_ fanout951/X _17454_/D vssd1 vssd1 vccd1 vccd1 _17454_/Q sky130_fd_sc_hd__dfxtp_1
X_11878_ _11878_/A _11878_/B vssd1 vssd1 vccd1 vccd1 _11888_/A sky130_fd_sc_hd__or2_1
X_13617_ _13618_/A _13618_/B vssd1 vssd1 vccd1 vccd1 _13617_/X sky130_fd_sc_hd__and2b_1
X_16405_ _16111_/A _16396_/Y _16398_/X _16304_/A _16404_/X vssd1 vssd1 vccd1 vccd1
+ _16405_/X sky130_fd_sc_hd__o221a_1
X_10829_ _10829_/A _10829_/B vssd1 vssd1 vccd1 vccd1 _11092_/B sky130_fd_sc_hd__xnor2_1
XFILLER_60_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17385_ _17385_/A _17389_/B vssd1 vssd1 vccd1 vccd1 _17385_/X sky130_fd_sc_hd__or2_1
X_14597_ _14597_/A _14597_/B vssd1 vssd1 vccd1 vccd1 _14618_/A sky130_fd_sc_hd__xnor2_1
XFILLER_158_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16336_ _16760_/B _16814_/B vssd1 vssd1 vccd1 vccd1 _16337_/B sky130_fd_sc_hd__nand2_1
X_13548_ _13425_/Y _13430_/A _13662_/B _13547_/X vssd1 vssd1 vccd1 vccd1 _13558_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_158_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16267_ _16268_/A _16268_/B vssd1 vssd1 vccd1 vccd1 _16267_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_145_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13479_ _13479_/A _13479_/B vssd1 vssd1 vccd1 vccd1 _13480_/B sky130_fd_sc_hd__nand2_1
XFILLER_65_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15218_ _15218_/A _15218_/B vssd1 vssd1 vccd1 vccd1 _15220_/B sky130_fd_sc_hd__xor2_1
XFILLER_133_409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16198_ _16290_/B _16198_/B vssd1 vssd1 vccd1 vccd1 _16200_/C sky130_fd_sc_hd__nand2b_1
XFILLER_127_984 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_770 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15149_ _16935_/A _15204_/B _16807_/A _16938_/A _15147_/A vssd1 vssd1 vccd1 vccd1
+ _15149_/X sky130_fd_sc_hd__o41a_1
XFILLER_142_954 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09710_ _10126_/B _10142_/B vssd1 vssd1 vccd1 vccd1 _09710_/Y sky130_fd_sc_hd__nand2_1
XFILLER_68_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09641_ _09642_/B _09642_/A vssd1 vssd1 vccd1 vccd1 _09645_/B sky130_fd_sc_hd__and2b_1
XFILLER_56_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09572_ _09573_/B _09573_/A vssd1 vssd1 vccd1 vccd1 _09581_/B sky130_fd_sc_hd__nand2b_1
XFILLER_83_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1012 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09006_ _09007_/A _09007_/B vssd1 vssd1 vccd1 vccd1 _09006_/X sky130_fd_sc_hd__or2_1
XFILLER_118_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout520 _10638_/B vssd1 vssd1 vccd1 vccd1 _11115_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_132_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout531 _14734_/A vssd1 vssd1 vccd1 vccd1 _14636_/A sky130_fd_sc_hd__buf_2
Xfanout542 _09899_/A vssd1 vssd1 vccd1 vccd1 _14789_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_116_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09908_ _09932_/A _09908_/B vssd1 vssd1 vccd1 vccd1 _09909_/C sky130_fd_sc_hd__and2_1
Xfanout553 _14889_/C vssd1 vssd1 vccd1 vccd1 _15628_/A sky130_fd_sc_hd__clkbuf_4
Xfanout564 _13627_/S vssd1 vssd1 vccd1 vccd1 _16011_/A sky130_fd_sc_hd__buf_2
Xfanout575 fanout578/X vssd1 vssd1 vccd1 vccd1 _10045_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout586 _17512_/Q vssd1 vssd1 vccd1 vccd1 _15126_/A sky130_fd_sc_hd__clkbuf_2
X_09839_ _10109_/B _10072_/B _09981_/D _09979_/A vssd1 vssd1 vccd1 vccd1 _09839_/Y
+ sky130_fd_sc_hd__a22oi_1
Xfanout597 _14794_/A vssd1 vssd1 vccd1 vccd1 _10545_/C sky130_fd_sc_hd__buf_2
XFILLER_47_938 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12850_ _17371_/A _12849_/X _12847_/X _16653_/A vssd1 vssd1 vccd1 vccd1 _12850_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_74_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11801_ _12025_/A _10657_/B _10543_/C vssd1 vssd1 vccd1 vccd1 _11802_/B sky130_fd_sc_hd__a21o_1
XTAP_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12781_ _12938_/A _12782_/B _12782_/C vssd1 vssd1 vccd1 vccd1 _12781_/X sky130_fd_sc_hd__a21o_1
XTAP_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14520_ _14519_/B _14519_/C _14519_/A vssd1 vssd1 vccd1 vccd1 _14520_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11732_ _11732_/A _11732_/B _11732_/C vssd1 vssd1 vccd1 vccd1 _11732_/Y sky130_fd_sc_hd__nor3_1
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14451_ _14451_/A _14567_/A vssd1 vssd1 vccd1 vccd1 _14454_/A sky130_fd_sc_hd__nor2_1
X_11663_ _11663_/A _11663_/B vssd1 vssd1 vccd1 vccd1 _11664_/B sky130_fd_sc_hd__and2_1
XTAP_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13402_ _13526_/B _13401_/B _13401_/C vssd1 vssd1 vccd1 vccd1 _13403_/B sky130_fd_sc_hd__a21o_1
XFILLER_174_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10614_ _10615_/A _10615_/B _10615_/C vssd1 vssd1 vccd1 vccd1 _10614_/X sky130_fd_sc_hd__a21o_2
X_17170_ _17150_/X _17156_/X _17169_/X _17170_/B1 _17153_/A vssd1 vssd1 vccd1 vccd1
+ _17574_/D sky130_fd_sc_hd__a32oi_2
X_14382_ _14382_/A _14382_/B vssd1 vssd1 vccd1 vccd1 _14396_/A sky130_fd_sc_hd__or2_1
X_11594_ _11630_/A _15116_/B vssd1 vssd1 vccd1 vccd1 _11628_/A sky130_fd_sc_hd__nand2_1
X_16121_ _11848_/Y _13832_/Y _16120_/X vssd1 vssd1 vccd1 vccd1 _16122_/C sky130_fd_sc_hd__a21oi_1
X_13333_ _13450_/B _13334_/C _13966_/D _14769_/A vssd1 vssd1 vccd1 vccd1 _13337_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_127_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10545_ _10546_/A _10544_/Y _10545_/C _10545_/D vssd1 vssd1 vccd1 vccd1 _10655_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_6_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16052_ _15964_/A _15964_/B _15962_/Y vssd1 vssd1 vccd1 vccd1 _16075_/A sky130_fd_sc_hd__a21oi_1
X_13264_ _13264_/A _13264_/B vssd1 vssd1 vccd1 vccd1 _13266_/B sky130_fd_sc_hd__nor2_1
XFILLER_155_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10476_ _11027_/A _10594_/B _11006_/C _10591_/A vssd1 vssd1 vccd1 vccd1 _10478_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_6_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_995 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15003_ _15056_/A _15003_/B _15450_/B vssd1 vssd1 vccd1 vccd1 _15003_/X sky130_fd_sc_hd__or3_1
X_12215_ _12700_/B _11816_/Y _12214_/Y vssd1 vssd1 vccd1 vccd1 _12216_/A sky130_fd_sc_hd__a21oi_1
X_13195_ _13195_/A _13195_/B vssd1 vssd1 vccd1 vccd1 _13197_/A sky130_fd_sc_hd__nor2_1
XFILLER_135_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12146_ _12146_/A _12146_/B vssd1 vssd1 vccd1 vccd1 _12148_/C sky130_fd_sc_hd__nand2_1
XFILLER_123_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16954_ _16758_/C _16893_/A _16935_/A _16758_/B vssd1 vssd1 vccd1 vccd1 _16955_/B
+ sky130_fd_sc_hd__o211a_1
X_12077_ _12077_/A _12077_/B _12077_/C _12077_/D vssd1 vssd1 vccd1 vccd1 _12078_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_49_242 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11028_ _11027_/B _10954_/D _11027_/D _11027_/A vssd1 vssd1 vccd1 vccd1 _11029_/B
+ sky130_fd_sc_hd__a22oi_1
X_15905_ _16015_/A _16014_/B _15898_/Y _15904_/X _15897_/X vssd1 vssd1 vccd1 vccd1
+ _15905_/X sky130_fd_sc_hd__o311a_1
XFILLER_37_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16885_ _16886_/A _16886_/B vssd1 vssd1 vccd1 vccd1 _16887_/A sky130_fd_sc_hd__nor2_1
XFILLER_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_415 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_223 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15836_ _15836_/A _15836_/B vssd1 vssd1 vccd1 vccd1 _15837_/B sky130_fd_sc_hd__xnor2_2
XFILLER_46_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15767_ _15866_/B _15767_/B vssd1 vssd1 vccd1 vccd1 _15769_/C sky130_fd_sc_hd__nor2_1
X_12979_ _12979_/A _12979_/B vssd1 vssd1 vccd1 vccd1 _12981_/B sky130_fd_sc_hd__xnor2_1
XFILLER_52_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17506_ fanout947/X _17506_/D vssd1 vssd1 vccd1 vccd1 _17506_/Q sky130_fd_sc_hd__dfxtp_1
X_14718_ _14747_/A _14718_/B vssd1 vssd1 vccd1 vccd1 _14719_/C sky130_fd_sc_hd__nand2_1
XFILLER_33_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15698_ _15698_/A _15698_/B vssd1 vssd1 vccd1 vccd1 _15700_/A sky130_fd_sc_hd__nor2_1
XFILLER_36_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17437_ fanout938/X _17437_/D vssd1 vssd1 vccd1 vccd1 _17437_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_21_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14649_ _14649_/A _14649_/B vssd1 vssd1 vccd1 vccd1 _14651_/B sky130_fd_sc_hd__xnor2_2
XFILLER_32_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_16 _16738_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_27 _17538_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_38 _14765_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17368_ input58/X _17377_/B _17367_/Y _17378_/C1 vssd1 vssd1 vccd1 vccd1 _17512_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA_49 _09899_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16319_ _16229_/A _16229_/B _16227_/B vssd1 vssd1 vccd1 vccd1 _16321_/B sky130_fd_sc_hd__a21o_1
XFILLER_9_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17299_ input47/X _17362_/C _17429_/C vssd1 vssd1 vccd1 vccd1 _17299_/X sky130_fd_sc_hd__or3_1
XFILLER_174_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_515 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput101 _17459_/Q vssd1 vssd1 vccd1 vccd1 o_wb_data[25] sky130_fd_sc_hd__clkbuf_1
XFILLER_127_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput112 _17440_/Q vssd1 vssd1 vccd1 vccd1 o_wb_data[6] sky130_fd_sc_hd__clkbuf_1
XFILLER_115_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_551 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09624_ _09624_/A _09624_/B _09624_/C vssd1 vssd1 vccd1 vccd1 _09625_/B sky130_fd_sc_hd__nor3_1
XFILLER_56_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09555_ _17397_/A _17395_/A _09555_/C _09555_/D vssd1 vssd1 vccd1 vccd1 _09556_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_71_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09486_ _09387_/A _09387_/B _09387_/C vssd1 vssd1 vccd1 vccd1 _09486_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_114 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10330_ _10330_/A _10330_/B vssd1 vssd1 vccd1 vccd1 _10333_/A sky130_fd_sc_hd__nand2_1
XFILLER_125_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_943 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10261_ _10261_/A _10261_/B _10261_/C vssd1 vssd1 vccd1 vccd1 _10262_/C sky130_fd_sc_hd__nand3_1
XFILLER_79_805 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12000_ _09122_/A _09255_/X _11998_/X _11999_/Y vssd1 vssd1 vccd1 vccd1 _12200_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_79_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10192_ _10193_/A _10192_/B _10207_/B _10192_/D vssd1 vssd1 vccd1 vccd1 _10193_/B
+ sky130_fd_sc_hd__nor4_2
XFILLER_105_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_79 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout350 _14153_/B vssd1 vssd1 vccd1 vccd1 _13977_/B sky130_fd_sc_hd__buf_2
Xfanout361 _09502_/A vssd1 vssd1 vccd1 vccd1 _17415_/A sky130_fd_sc_hd__buf_4
XFILLER_4_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout372 _13893_/A vssd1 vssd1 vccd1 vccd1 _14318_/B sky130_fd_sc_hd__clkbuf_2
X_13951_ _13951_/A _13951_/B vssd1 vssd1 vccd1 vccd1 _13954_/C sky130_fd_sc_hd__xnor2_1
Xfanout383 _12788_/A vssd1 vssd1 vccd1 vccd1 _13689_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_87_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout394 _14772_/A vssd1 vssd1 vccd1 vccd1 _10321_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_19_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12902_ _12902_/A _12902_/B _12902_/C vssd1 vssd1 vccd1 vccd1 _12918_/B sky130_fd_sc_hd__nand3_1
XFILLER_4_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16670_ _16670_/A _16670_/B _16670_/C vssd1 vssd1 vccd1 vccd1 _16751_/A sky130_fd_sc_hd__nand3_1
X_13882_ _13882_/A _13882_/B vssd1 vssd1 vccd1 vccd1 _13885_/A sky130_fd_sc_hd__xnor2_1
XFILLER_19_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12833_ _12991_/B _12834_/B _12834_/C vssd1 vssd1 vccd1 vccd1 _12833_/Y sky130_fd_sc_hd__nor3_1
XFILLER_74_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15621_ _15621_/A _15621_/B vssd1 vssd1 vccd1 vccd1 _15621_/Y sky130_fd_sc_hd__xnor2_1
XTAP_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_470 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15552_ _16315_/D _15552_/B vssd1 vssd1 vccd1 vccd1 _15552_/X sky130_fd_sc_hd__or2_1
X_12764_ _12764_/A _12764_/B _12764_/C vssd1 vssd1 vccd1 vccd1 _12766_/C sky130_fd_sc_hd__and3_1
XFILLER_14_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11715_ _16295_/A _16206_/A _16206_/B vssd1 vssd1 vccd1 vccd1 _16387_/B sky130_fd_sc_hd__and3_1
X_14503_ _14441_/B _14443_/B _14441_/A vssd1 vssd1 vccd1 vccd1 _14505_/B sky130_fd_sc_hd__o21ba_1
X_15483_ _15484_/A _15567_/A vssd1 vssd1 vccd1 vccd1 _15483_/Y sky130_fd_sc_hd__nand2_1
XFILLER_30_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12695_ _12372_/X _12538_/Y _12539_/Y vssd1 vssd1 vccd1 vccd1 _12695_/X sky130_fd_sc_hd__a21o_1
XTAP_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17222_ _17583_/Q _17225_/A2 _17225_/B1 vssd1 vssd1 vccd1 vccd1 _17222_/X sky130_fd_sc_hd__a21o_1
X_11646_ _11646_/A _11646_/B _11646_/C vssd1 vssd1 vccd1 vccd1 _15524_/C sky130_fd_sc_hd__and3_1
X_14434_ _14492_/A vssd1 vssd1 vccd1 vccd1 _14434_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_668 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput14 i_wb_addr[1] vssd1 vssd1 vccd1 vccd1 input14/X sky130_fd_sc_hd__clkbuf_1
XFILLER_122_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput25 i_wb_addr[2] vssd1 vssd1 vccd1 vccd1 input25/X sky130_fd_sc_hd__dlymetal6s2s_1
X_14365_ _14440_/B _14365_/B vssd1 vssd1 vccd1 vccd1 _14400_/A sky130_fd_sc_hd__nor2_1
X_17153_ _17153_/A _17153_/B vssd1 vssd1 vccd1 vccd1 _17153_/X sky130_fd_sc_hd__and2_1
X_11577_ _11582_/A _11577_/B vssd1 vssd1 vccd1 vccd1 _11579_/B sky130_fd_sc_hd__nor2_1
Xinput36 i_wb_data[0] vssd1 vssd1 vccd1 vccd1 input36/X sky130_fd_sc_hd__clkbuf_2
XFILLER_156_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput47 i_wb_data[1] vssd1 vssd1 vccd1 vccd1 input47/X sky130_fd_sc_hd__clkbuf_2
X_16104_ _11465_/A _11465_/B _11707_/Y vssd1 vssd1 vccd1 vccd1 _16105_/B sky130_fd_sc_hd__o21ai_1
X_13316_ _13317_/A _13317_/B _13317_/C vssd1 vssd1 vccd1 vccd1 _13316_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_10_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput58 i_wb_data[2] vssd1 vssd1 vccd1 vccd1 input58/X sky130_fd_sc_hd__clkbuf_2
X_10528_ _10528_/A _10626_/A vssd1 vssd1 vccd1 vccd1 _10536_/A sky130_fd_sc_hd__nor2_1
XFILLER_128_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17084_ _17085_/A _17085_/B _17085_/C vssd1 vssd1 vccd1 vccd1 _17086_/A sky130_fd_sc_hd__o21ai_1
Xinput69 i_wb_we vssd1 vssd1 vccd1 vccd1 input69/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_128_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14296_ _14297_/A _14297_/B vssd1 vssd1 vccd1 vccd1 _14296_/X sky130_fd_sc_hd__and2b_1
XFILLER_7_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16035_ _16035_/A _16035_/B vssd1 vssd1 vccd1 vccd1 _16036_/B sky130_fd_sc_hd__xor2_2
XFILLER_6_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13247_ _13248_/A _13248_/B _13248_/C vssd1 vssd1 vccd1 vccd1 _13249_/C sky130_fd_sc_hd__o21ai_2
XFILLER_171_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10459_ _10459_/A _10459_/B _10459_/C vssd1 vssd1 vccd1 vccd1 _10459_/Y sky130_fd_sc_hd__nand3_1
X_13178_ _13178_/A _13178_/B _13178_/C vssd1 vssd1 vccd1 vccd1 _13312_/B sky130_fd_sc_hd__and3_1
XFILLER_123_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12129_ _17421_/A _12129_/B vssd1 vssd1 vccd1 vccd1 _12131_/B sky130_fd_sc_hd__nand2_1
XFILLER_85_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16937_ _16937_/A _16937_/B vssd1 vssd1 vccd1 vccd1 _16943_/A sky130_fd_sc_hd__nor2_1
XFILLER_77_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16868_ _16868_/A _16868_/B vssd1 vssd1 vccd1 vccd1 _16872_/A sky130_fd_sc_hd__nor2_1
XFILLER_37_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15819_ _15918_/A _16743_/C _17043_/B _15726_/A vssd1 vssd1 vccd1 vccd1 _15821_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_80_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16799_ _16796_/B _16799_/A2 _16799_/B1 _14863_/A _16869_/C1 vssd1 vssd1 vccd1 vccd1
+ _16799_/X sky130_fd_sc_hd__a221o_1
X_09340_ _09391_/B _09391_/C _09391_/A vssd1 vssd1 vccd1 vccd1 _09395_/B sky130_fd_sc_hd__a21oi_2
XFILLER_61_760 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09271_ _12077_/B _11961_/B _09272_/D _09414_/A vssd1 vssd1 vccd1 vccd1 _09273_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_61_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_112 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_835 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08986_ _08985_/A _09074_/A vssd1 vssd1 vccd1 vccd1 _09014_/A sky130_fd_sc_hd__and2b_1
XFILLER_57_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_798 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09607_ _09607_/A _09735_/A vssd1 vssd1 vccd1 vccd1 _09614_/A sky130_fd_sc_hd__nor2_1
XFILLER_83_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_535 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09538_ _09538_/A _09538_/B vssd1 vssd1 vccd1 vccd1 _09678_/A sky130_fd_sc_hd__xor2_1
XFILLER_58_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09469_ _09473_/A _09591_/A _09473_/C vssd1 vssd1 vccd1 vccd1 _09478_/B sky130_fd_sc_hd__o21ai_1
XFILLER_24_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_495 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11500_ _11499_/A _11539_/A _11456_/X _11490_/Y vssd1 vssd1 vccd1 vccd1 _11502_/B
+ sky130_fd_sc_hd__o211a_2
XFILLER_157_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12480_ _12481_/A _12481_/B _12481_/C vssd1 vssd1 vccd1 vccd1 _12480_/X sky130_fd_sc_hd__and3_1
XFILLER_132_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11431_ _11430_/A _11475_/A vssd1 vssd1 vccd1 vccd1 _11433_/B sky130_fd_sc_hd__nand2b_1
XFILLER_22_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_651 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14150_ _14150_/A _14150_/B _14150_/C vssd1 vssd1 vccd1 vccd1 _14151_/B sky130_fd_sc_hd__nor3_1
X_11362_ _11362_/A _11362_/B vssd1 vssd1 vccd1 vccd1 _11492_/B sky130_fd_sc_hd__xnor2_1
XFILLER_165_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13101_ _13101_/A _13101_/B vssd1 vssd1 vccd1 vccd1 _13103_/B sky130_fd_sc_hd__xnor2_1
XFILLER_138_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10313_ _10314_/B _10314_/A vssd1 vssd1 vccd1 vccd1 _10450_/A sky130_fd_sc_hd__and2b_1
X_14081_ _14081_/A _14173_/A vssd1 vssd1 vccd1 vccd1 _14084_/A sky130_fd_sc_hd__nor2_1
X_11293_ _11293_/A _11293_/B vssd1 vssd1 vccd1 vccd1 _11294_/B sky130_fd_sc_hd__nand2_1
XFILLER_3_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13032_ _13033_/A _13033_/B _13033_/C vssd1 vssd1 vccd1 vccd1 _13046_/A sky130_fd_sc_hd__a21o_1
XFILLER_106_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10244_ _10244_/A _14788_/B vssd1 vssd1 vccd1 vccd1 _10245_/B sky130_fd_sc_hd__nand2_1
XFILLER_140_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10175_ _10288_/A _10296_/A _10288_/C vssd1 vssd1 vccd1 vccd1 _10289_/A sky130_fd_sc_hd__o21ai_1
XFILLER_120_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout180 _16334_/C vssd1 vssd1 vccd1 vccd1 _16747_/A sky130_fd_sc_hd__buf_4
XFILLER_59_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14983_ _10182_/C _14981_/Y _14982_/Y _15097_/A vssd1 vssd1 vccd1 vccd1 _14983_/X
+ sky130_fd_sc_hd__a211o_1
Xfanout191 _15151_/X vssd1 vssd1 vccd1 vccd1 _16317_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_75_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16722_ _16722_/A _17153_/B vssd1 vssd1 vccd1 vccd1 _16723_/B sky130_fd_sc_hd__nor2_1
X_13934_ _13935_/A _13935_/B vssd1 vssd1 vccd1 vccd1 _13934_/Y sky130_fd_sc_hd__nor2_1
XFILLER_47_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16653_ _16653_/A _16653_/B vssd1 vssd1 vccd1 vccd1 _16653_/X sky130_fd_sc_hd__or2_1
XFILLER_74_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13865_ _14213_/B _13866_/C _13866_/D _14213_/A vssd1 vssd1 vccd1 vccd1 _13867_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_34_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15604_ _15604_/A _15604_/B vssd1 vssd1 vccd1 vccd1 _15607_/A sky130_fd_sc_hd__xnor2_1
X_12816_ _12816_/A _12816_/B vssd1 vssd1 vccd1 vccd1 _12817_/B sky130_fd_sc_hd__xnor2_1
XFILLER_15_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16584_ _16304_/A _16577_/X _16583_/X _16569_/X vssd1 vssd1 vccd1 vccd1 _16584_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_43_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13796_ _14176_/A _13993_/B _13796_/C vssd1 vssd1 vccd1 vccd1 _13906_/B sky130_fd_sc_hd__nand3_1
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15535_ _16485_/A _15535_/B vssd1 vssd1 vccd1 vccd1 _15535_/Y sky130_fd_sc_hd__nand2_1
X_12747_ _12747_/A _12747_/B vssd1 vssd1 vccd1 vccd1 _12766_/A sky130_fd_sc_hd__xnor2_1
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12678_ _12676_/A _12676_/B _12676_/C vssd1 vssd1 vccd1 vccd1 _12679_/B sky130_fd_sc_hd__o21ai_1
X_15466_ _16015_/A _15541_/B _15463_/Y _15465_/Y _15462_/Y vssd1 vssd1 vccd1 vccd1
+ _15467_/D sky130_fd_sc_hd__o311a_1
X_17205_ _17545_/Q _17274_/B vssd1 vssd1 vccd1 vccd1 _17205_/X sky130_fd_sc_hd__and2_1
X_11629_ _11629_/A _11629_/B _15116_/B _11629_/D vssd1 vssd1 vccd1 vccd1 _11632_/A
+ sky130_fd_sc_hd__and4_1
X_14417_ _14284_/B _14534_/A _14415_/X vssd1 vssd1 vccd1 vccd1 _14419_/B sky130_fd_sc_hd__a21o_1
XFILLER_128_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15397_ _15397_/A _16152_/A vssd1 vssd1 vccd1 vccd1 _15832_/A sky130_fd_sc_hd__nand2_1
XFILLER_156_662 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17136_ _17099_/Y _17102_/X _17133_/Y _17134_/X vssd1 vssd1 vccd1 vccd1 _17136_/X
+ sky130_fd_sc_hd__a211o_1
X_14348_ _14348_/A _14348_/B vssd1 vssd1 vccd1 vccd1 _14350_/C sky130_fd_sc_hd__xnor2_1
XFILLER_155_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_846 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14279_ _14279_/A _14279_/B vssd1 vssd1 vccd1 vccd1 _14279_/Y sky130_fd_sc_hd__nor2_1
X_17067_ _17018_/Y _17066_/X _17065_/X _17064_/X vssd1 vssd1 vccd1 vccd1 _17067_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_144_879 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16018_ _15996_/Y _15998_/X _16017_/X _16494_/B1 _16014_/A vssd1 vssd1 vccd1 vccd1
+ _16019_/A sky130_fd_sc_hd__a32o_1
XFILLER_170_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08840_ _08913_/A _09728_/B _09319_/C _09319_/D vssd1 vssd1 vccd1 vccd1 _08843_/A
+ sky130_fd_sc_hd__and4_1
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08771_ _17399_/A _09030_/C _09272_/D _17403_/A vssd1 vssd1 vccd1 vccd1 _08772_/D
+ sky130_fd_sc_hd__a22o_1
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_798 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09323_ _09323_/A _09323_/B vssd1 vssd1 vccd1 vccd1 _09328_/C sky130_fd_sc_hd__nor2_1
XFILLER_21_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_966 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09254_ _09255_/B _09255_/C vssd1 vssd1 vccd1 vccd1 _09256_/B sky130_fd_sc_hd__nand2_1
X_09185_ _17411_/A _09267_/D _12174_/D _09942_/A vssd1 vssd1 vccd1 vccd1 _09189_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_88_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_857 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08969_ _09493_/A _11932_/B _08969_/C vssd1 vssd1 vccd1 vccd1 _08973_/B sky130_fd_sc_hd__and3_1
XFILLER_69_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11980_ _11980_/A _11980_/B vssd1 vssd1 vccd1 vccd1 _11982_/B sky130_fd_sc_hd__xnor2_1
XFILLER_56_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10931_ _14788_/A _10971_/B _10922_/X _14806_/A _10800_/C vssd1 vssd1 vccd1 vccd1
+ _10938_/A sky130_fd_sc_hd__a32o_1
XFILLER_17_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10862_ _10861_/A _10861_/B _10861_/C vssd1 vssd1 vccd1 vccd1 _10863_/C sky130_fd_sc_hd__a21oi_1
XFILLER_140_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13650_ _13648_/X _13650_/B vssd1 vssd1 vccd1 vccd1 _13652_/A sky130_fd_sc_hd__and2b_1
XFILLER_72_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12601_ _12446_/A _12448_/B _12446_/B vssd1 vssd1 vccd1 vccd1 _12603_/B sky130_fd_sc_hd__o21ba_1
XFILLER_140_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13581_ _13977_/A _13977_/B _13966_/D _13866_/D vssd1 vssd1 vccd1 vccd1 _13582_/B
+ sky130_fd_sc_hd__and4_1
XPHY_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10793_ _11132_/B _10897_/B _10933_/C _11629_/A vssd1 vssd1 vccd1 vccd1 _10794_/B
+ sky130_fd_sc_hd__a22oi_1
XPHY_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_730 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12532_ _12534_/A _12534_/B vssd1 vssd1 vccd1 vccd1 _12532_/Y sky130_fd_sc_hd__nand2b_1
X_15320_ _15386_/A _15313_/Y _15319_/X _16582_/A vssd1 vssd1 vccd1 vccd1 _15321_/D
+ sky130_fd_sc_hd__o2bb2a_1
XPHY_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_62 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15251_ _16485_/A _15243_/Y _15244_/X _15250_/X vssd1 vssd1 vccd1 vccd1 _15257_/C
+ sky130_fd_sc_hd__a31o_1
X_12463_ _12770_/A _12770_/B _12618_/D _12463_/D vssd1 vssd1 vccd1 vccd1 _12662_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_138_651 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11414_ _11299_/B _11299_/C _11299_/A vssd1 vssd1 vccd1 vccd1 _11415_/B sky130_fd_sc_hd__o21ai_1
XFILLER_126_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14202_ _14202_/A _14202_/B _14202_/C vssd1 vssd1 vccd1 vccd1 _14204_/A sky130_fd_sc_hd__and3_1
X_15182_ _11321_/X _14790_/Y _14798_/Y vssd1 vssd1 vccd1 vccd1 _15182_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_166_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12394_ _12394_/A vssd1 vssd1 vccd1 vccd1 _12394_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_126_846 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14133_ _13947_/Y _14042_/Y _14218_/A vssd1 vssd1 vccd1 vccd1 _14134_/C sky130_fd_sc_hd__a21o_1
X_11345_ _11345_/A _11345_/B vssd1 vssd1 vccd1 vccd1 _11357_/A sky130_fd_sc_hd__xor2_1
XFILLER_152_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14064_ _14064_/A _14064_/B vssd1 vssd1 vccd1 vccd1 _14066_/A sky130_fd_sc_hd__nor2_1
X_11276_ _11137_/C _11276_/B vssd1 vssd1 vccd1 vccd1 _11283_/A sky130_fd_sc_hd__and2b_1
XFILLER_98_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13015_ _17371_/A _13015_/B vssd1 vssd1 vccd1 vccd1 _13015_/Y sky130_fd_sc_hd__nor2_1
X_10227_ _10219_/A _10219_/C _10219_/B vssd1 vssd1 vccd1 vccd1 _10342_/B sky130_fd_sc_hd__o21ai_1
XFILLER_67_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10158_ _10157_/C _10157_/Y _10028_/B _10104_/X vssd1 vssd1 vccd1 vccd1 _10193_/A
+ sky130_fd_sc_hd__a211oi_2
X_14966_ _15147_/C _15208_/C _14877_/Y vssd1 vssd1 vccd1 vccd1 _14966_/X sky130_fd_sc_hd__a21o_1
X_10089_ _10081_/A _10084_/A _10090_/A _10088_/X vssd1 vssd1 vccd1 vccd1 _10101_/A
+ sky130_fd_sc_hd__a211oi_1
XFILLER_47_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16705_ _16705_/A _16705_/B vssd1 vssd1 vccd1 vccd1 _16706_/B sky130_fd_sc_hd__nand2_1
XFILLER_63_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13917_ _13918_/A _13918_/B vssd1 vssd1 vccd1 vccd1 _14018_/B sky130_fd_sc_hd__nand2_1
XFILLER_35_524 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14897_ _15463_/A _15208_/C _15208_/D _14897_/D vssd1 vssd1 vccd1 vccd1 _14899_/C
+ sky130_fd_sc_hd__or4_2
X_16636_ _16636_/A _16636_/B _16636_/C vssd1 vssd1 vccd1 vccd1 _16637_/B sky130_fd_sc_hd__and3_1
X_13848_ _13848_/A _13848_/B vssd1 vssd1 vccd1 vccd1 _13849_/C sky130_fd_sc_hd__xnor2_1
XFILLER_62_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16567_ _16566_/A _16566_/B _17063_/A vssd1 vssd1 vccd1 vccd1 _16567_/X sky130_fd_sc_hd__a21o_1
X_13779_ _13779_/A _13779_/B vssd1 vssd1 vccd1 vccd1 _13781_/A sky130_fd_sc_hd__nor2_1
XFILLER_95_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15518_ _15518_/A _15518_/B vssd1 vssd1 vccd1 vccd1 _15520_/C sky130_fd_sc_hd__xnor2_1
X_16498_ _16498_/A _16609_/A vssd1 vssd1 vccd1 vccd1 _16499_/C sky130_fd_sc_hd__nand2_1
XFILLER_149_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15449_ _15532_/A vssd1 vssd1 vccd1 vccd1 _15449_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_802 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_695 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_846 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17119_ _17119_/A _17119_/B _17119_/C vssd1 vssd1 vccd1 vccd1 _17121_/A sky130_fd_sc_hd__and3_1
Xmax_cap122 _14337_/Y vssd1 vssd1 vccd1 vccd1 _14404_/C1 sky130_fd_sc_hd__clkbuf_1
XFILLER_116_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09941_ _09941_/A _09941_/B vssd1 vssd1 vccd1 vccd1 _09948_/A sky130_fd_sc_hd__nor2_1
XFILLER_131_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout905 _10062_/B vssd1 vssd1 vccd1 vccd1 _09502_/B sky130_fd_sc_hd__buf_2
Xfanout916 _17172_/Y vssd1 vssd1 vccd1 vccd1 _17225_/B1 sky130_fd_sc_hd__clkbuf_4
Xfanout927 _17358_/C1 vssd1 vssd1 vccd1 vccd1 _17408_/C1 sky130_fd_sc_hd__clkbuf_2
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09872_ _09872_/A _09872_/B vssd1 vssd1 vccd1 vccd1 _09878_/A sky130_fd_sc_hd__nor2_1
XFILLER_140_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout938 fanout939/X vssd1 vssd1 vccd1 vccd1 fanout938/X sky130_fd_sc_hd__buf_2
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout949 fanout950/X vssd1 vssd1 vccd1 vccd1 fanout949/X sky130_fd_sc_hd__buf_2
XFILLER_85_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08823_ _17391_/A _17389_/A _09446_/D _09042_/B vssd1 vssd1 vccd1 vccd1 _08826_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_100_724 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08754_ _17401_/A _12166_/B _08754_/C _08754_/D vssd1 vssd1 vccd1 vccd1 _08768_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_57_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_8 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_527 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_45 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09306_ _09306_/A _09306_/B vssd1 vssd1 vccd1 vccd1 _09438_/B sky130_fd_sc_hd__nor2_1
XFILLER_167_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09237_ _09238_/A _09238_/B _09238_/C vssd1 vssd1 vccd1 vccd1 _09239_/A sky130_fd_sc_hd__o21a_1
XFILLER_155_919 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_278 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09168_ _09168_/A _09168_/B vssd1 vssd1 vccd1 vccd1 _09333_/B sky130_fd_sc_hd__xnor2_1
XFILLER_147_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09099_ _10180_/A _09350_/B _14978_/A vssd1 vssd1 vccd1 vccd1 _09099_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_134_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11130_ _11130_/A _11130_/B _11130_/C vssd1 vssd1 vccd1 vccd1 _11139_/B sky130_fd_sc_hd__nand3_1
XFILLER_122_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11061_ _11061_/A _11077_/A _11061_/C vssd1 vssd1 vccd1 vccd1 _11065_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10012_ _10018_/A _10018_/B vssd1 vssd1 vccd1 vccd1 _10019_/A sky130_fd_sc_hd__nor2_1
XFILLER_95_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14820_ _16729_/B _16730_/A _13459_/A vssd1 vssd1 vccd1 vccd1 _16797_/A sky130_fd_sc_hd__a21o_1
XFILLER_76_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14751_ _14751_/A _14751_/B vssd1 vssd1 vccd1 vccd1 _14755_/A sky130_fd_sc_hd__nand2_1
XFILLER_91_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11963_ _12169_/B _11963_/B vssd1 vssd1 vccd1 vccd1 _11966_/B sky130_fd_sc_hd__nand2_1
XFILLER_91_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13702_ _13702_/A _13702_/B _13702_/C vssd1 vssd1 vccd1 vccd1 _13703_/B sky130_fd_sc_hd__and3_1
X_17470_ fanout955/X _17543_/Q vssd1 vssd1 vccd1 vccd1 _17470_/Q sky130_fd_sc_hd__dfxtp_1
X_10914_ _10914_/A _10914_/B vssd1 vssd1 vccd1 vccd1 _10915_/B sky130_fd_sc_hd__nor2_1
X_11894_ _11895_/B _11895_/C _11895_/D _17379_/A vssd1 vssd1 vccd1 vccd1 _11894_/Y
+ sky130_fd_sc_hd__a22oi_1
X_14682_ _14682_/A _14682_/B vssd1 vssd1 vccd1 vccd1 _14719_/A sky130_fd_sc_hd__xnor2_2
XFILLER_32_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16421_ _16422_/A _16422_/B vssd1 vssd1 vccd1 vccd1 _16423_/A sky130_fd_sc_hd__or2_1
X_10845_ _10846_/A _10846_/B vssd1 vssd1 vccd1 vccd1 _10943_/B sky130_fd_sc_hd__nand2_1
X_13633_ _13846_/A _13735_/D vssd1 vssd1 vccd1 vccd1 _13635_/C sky130_fd_sc_hd__nand2_1
XFILLER_25_590 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16352_ _16352_/A _16809_/C _16352_/C vssd1 vssd1 vccd1 vccd1 _16354_/A sky130_fd_sc_hd__and3_1
X_10776_ _10678_/B _10691_/X _10774_/A _11722_/A vssd1 vssd1 vccd1 vccd1 _10777_/C
+ sky130_fd_sc_hd__a211oi_1
XFILLER_9_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13564_ _14167_/A _13893_/A _13564_/C _14141_/D vssd1 vssd1 vccd1 vccd1 _13695_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_40_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15303_ _15303_/A _15303_/B vssd1 vssd1 vccd1 vccd1 _15303_/Y sky130_fd_sc_hd__nand2_1
XFILLER_9_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12515_ _12670_/A _12515_/B vssd1 vssd1 vccd1 vccd1 _12517_/B sky130_fd_sc_hd__nor2_1
X_16283_ _16283_/A _16283_/B vssd1 vssd1 vccd1 vccd1 _16285_/A sky130_fd_sc_hd__xor2_1
X_13495_ _13495_/A _13495_/B vssd1 vssd1 vccd1 vccd1 _13498_/A sky130_fd_sc_hd__nor2_1
XFILLER_139_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12446_ _12446_/A _12446_/B vssd1 vssd1 vccd1 vccd1 _12448_/A sky130_fd_sc_hd__nor2_1
X_15234_ _15233_/A _15233_/B _08743_/A vssd1 vssd1 vccd1 vccd1 _15234_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_166_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12377_ _12377_/A _12377_/B vssd1 vssd1 vccd1 vccd1 _12377_/Y sky130_fd_sc_hd__nor2_1
X_15165_ _15165_/A _15230_/A vssd1 vssd1 vccd1 vccd1 _15166_/B sky130_fd_sc_hd__nand2_1
XFILLER_99_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11328_ _11369_/A _11369_/B vssd1 vssd1 vccd1 vccd1 _11331_/C sky130_fd_sc_hd__nand2_1
XFILLER_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14116_ _14117_/A _14117_/B vssd1 vssd1 vccd1 vccd1 _14202_/B sky130_fd_sc_hd__nand2b_1
XFILLER_113_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15096_ _14978_/Y _14981_/Y _15096_/S vssd1 vssd1 vccd1 vccd1 _15097_/B sky130_fd_sc_hd__mux2_1
XFILLER_153_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11259_ _15373_/C _11561_/D _11592_/B _15396_/A vssd1 vssd1 vccd1 vccd1 _11259_/Y
+ sky130_fd_sc_hd__a22oi_1
X_14047_ _14047_/A _14047_/B vssd1 vssd1 vccd1 vccd1 _14048_/B sky130_fd_sc_hd__and2_1
XFILLER_113_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15998_ _15998_/A _15998_/B _11707_/Y vssd1 vssd1 vccd1 vccd1 _15998_/X sky130_fd_sc_hd__or3b_2
XFILLER_94_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14949_ _14949_/A _14949_/B vssd1 vssd1 vccd1 vccd1 _14949_/Y sky130_fd_sc_hd__nor2_1
XFILLER_36_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16619_ _16619_/A _16827_/D _16695_/C vssd1 vssd1 vccd1 vccd1 _16774_/A sky130_fd_sc_hd__or3_2
XFILLER_62_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17599_ fanout936/X _17599_/D vssd1 vssd1 vccd1 vccd1 _17599_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09022_ _09027_/A _09027_/B vssd1 vssd1 vccd1 vccd1 _09033_/A sky130_fd_sc_hd__nor2_1
XFILLER_164_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout702 _16654_/B2 vssd1 vssd1 vccd1 vccd1 _14213_/D sky130_fd_sc_hd__clkbuf_4
X_09924_ _10182_/C _09926_/B _09783_/A _09781_/Y vssd1 vssd1 vccd1 vccd1 _09930_/B
+ sky130_fd_sc_hd__o2bb2a_1
Xfanout713 _12079_/B vssd1 vssd1 vccd1 vccd1 _09319_/D sky130_fd_sc_hd__buf_2
XFILLER_172_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout724 _17497_/Q vssd1 vssd1 vccd1 vccd1 _10657_/B sky130_fd_sc_hd__buf_4
Xfanout735 _16298_/A vssd1 vssd1 vccd1 vccd1 _13866_/D sky130_fd_sc_hd__buf_2
XFILLER_86_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout746 _10993_/D vssd1 vssd1 vccd1 vccd1 _10534_/D sky130_fd_sc_hd__buf_2
XFILLER_98_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_722 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout757 _17493_/Q vssd1 vssd1 vccd1 vccd1 _16114_/A sky130_fd_sc_hd__buf_2
X_09855_ _10254_/A _10126_/B _10142_/B _10270_/B vssd1 vssd1 vccd1 vccd1 _09855_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_140_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout768 _10532_/D vssd1 vssd1 vccd1 vccd1 _10016_/D sky130_fd_sc_hd__buf_4
XFILLER_85_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_34 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout779 _10743_/C vssd1 vssd1 vccd1 vccd1 _15898_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_86_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08806_ _17399_/A _11961_/B _12340_/B _17403_/A vssd1 vssd1 vccd1 vccd1 _08806_/Y
+ sky130_fd_sc_hd__a22oi_1
XTAP_3106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09786_ _09786_/A _09786_/B vssd1 vssd1 vccd1 vccd1 _09932_/B sky130_fd_sc_hd__or2_1
XTAP_3117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_980 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08737_ _14929_/A vssd1 vssd1 vccd1 vccd1 _08737_/Y sky130_fd_sc_hd__inv_2
XTAP_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10630_ _10499_/Y _10589_/X _10598_/X _10611_/Y vssd1 vssd1 vccd1 vccd1 _10632_/D
+ sky130_fd_sc_hd__o211ai_4
XFILLER_167_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10561_ _10561_/A _11749_/A vssd1 vssd1 vccd1 vccd1 _10671_/B sky130_fd_sc_hd__or2_1
XFILLER_155_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12300_ _12508_/B _12300_/B vssd1 vssd1 vccd1 vccd1 _12307_/A sky130_fd_sc_hd__nor2_1
XFILLER_14_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13280_ _13280_/A _13280_/B vssd1 vssd1 vccd1 vccd1 _13282_/A sky130_fd_sc_hd__nor2_1
X_10492_ _11006_/B _14849_/A _10703_/B _10954_/A vssd1 vssd1 vccd1 vccd1 _10493_/B
+ sky130_fd_sc_hd__a22oi_1
XFILLER_10_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12231_ _11849_/A _12227_/X _12230_/X _16735_/A vssd1 vssd1 vccd1 vccd1 _12231_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_30_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12162_ _12162_/A _12325_/B vssd1 vssd1 vccd1 vccd1 _12163_/C sky130_fd_sc_hd__nor2_1
XFILLER_108_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11113_ _11112_/A _11112_/C _11112_/B vssd1 vssd1 vccd1 vccd1 _11113_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_146_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12093_ _12093_/A _12093_/B _12093_/C vssd1 vssd1 vccd1 vccd1 _12094_/B sky130_fd_sc_hd__or3_1
XFILLER_1_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16970_ _16970_/A _16970_/B vssd1 vssd1 vccd1 vccd1 _16971_/B sky130_fd_sc_hd__nand2_1
XFILLER_111_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11044_ _11058_/A _11058_/B vssd1 vssd1 vccd1 vccd1 _11048_/A sky130_fd_sc_hd__nand2b_1
X_15921_ _15921_/A _15921_/B vssd1 vssd1 vccd1 vccd1 _15923_/B sky130_fd_sc_hd__xnor2_1
XFILLER_89_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15852_ _15853_/A _15853_/B vssd1 vssd1 vccd1 vccd1 _15852_/Y sky130_fd_sc_hd__nand2_1
XFILLER_36_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14803_ _14803_/A _14803_/B vssd1 vssd1 vccd1 vccd1 _14803_/Y sky130_fd_sc_hd__nor2_1
X_15783_ _15784_/A _15784_/B vssd1 vssd1 vccd1 vccd1 _15883_/B sky130_fd_sc_hd__and2_1
X_12995_ _17405_/A _13208_/C _12801_/A _12799_/A vssd1 vssd1 vccd1 vccd1 _12996_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_57_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17522_ fanout942/X _17522_/D vssd1 vssd1 vccd1 vccd1 _17522_/Q sky130_fd_sc_hd__dfxtp_4
X_14734_ _14734_/A _14734_/B vssd1 vssd1 vccd1 vccd1 _14734_/Y sky130_fd_sc_hd__nand2_1
X_11946_ _11943_/Y _11944_/X _09006_/X _09010_/A vssd1 vssd1 vccd1 vccd1 _11947_/D
+ sky130_fd_sc_hd__o211ai_1
XFILLER_91_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17453_ fanout951/X _17453_/D vssd1 vssd1 vccd1 vccd1 _17453_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14665_ _14763_/S _14663_/Y _14664_/X _14636_/Y _14637_/X vssd1 vssd1 vccd1 vccd1
+ _17602_/D sky130_fd_sc_hd__a32o_1
XTAP_2994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11877_ _11877_/A _11877_/B _11877_/C vssd1 vssd1 vccd1 vccd1 _11891_/B sky130_fd_sc_hd__and3_1
XFILLER_60_655 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16404_ _16404_/A _16404_/B _16404_/C vssd1 vssd1 vccd1 vccd1 _16404_/X sky130_fd_sc_hd__and3_1
X_13616_ _13618_/B _13618_/A vssd1 vssd1 vccd1 vccd1 _13616_/Y sky130_fd_sc_hd__nand2b_1
X_10828_ _10828_/A _10828_/B vssd1 vssd1 vccd1 vccd1 _11092_/A sky130_fd_sc_hd__xnor2_1
XFILLER_158_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17384_ input37/X _17426_/A2 _17383_/X _17388_/C1 vssd1 vssd1 vccd1 vccd1 _17520_/D
+ sky130_fd_sc_hd__o211a_1
X_14596_ _14676_/A _14641_/C vssd1 vssd1 vccd1 vccd1 _14596_/Y sky130_fd_sc_hd__nand2_1
XFILLER_60_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16335_ _16333_/X _16335_/B vssd1 vssd1 vccd1 vccd1 _16337_/A sky130_fd_sc_hd__nand2b_1
X_13547_ _13662_/A _13545_/X _13418_/A _13419_/Y vssd1 vssd1 vccd1 vccd1 _13547_/X
+ sky130_fd_sc_hd__o211a_1
X_10759_ _11726_/A _10759_/B vssd1 vssd1 vccd1 vccd1 _10760_/C sky130_fd_sc_hd__and2_1
XFILLER_71_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16266_ _16266_/A _16266_/B vssd1 vssd1 vccd1 vccd1 _16268_/B sky130_fd_sc_hd__xor2_1
X_13478_ _13479_/A _13479_/B vssd1 vssd1 vccd1 vccd1 _13595_/A sky130_fd_sc_hd__or2_1
XFILLER_69_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15217_ _15218_/A _15218_/B vssd1 vssd1 vccd1 vccd1 _15283_/A sky130_fd_sc_hd__or2_1
XFILLER_127_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12429_ _12429_/A _12429_/B _12429_/C vssd1 vssd1 vccd1 vccd1 _12430_/B sky130_fd_sc_hd__nor3_1
X_16197_ _16197_/A _16197_/B _16195_/Y vssd1 vssd1 vccd1 vccd1 _16198_/B sky130_fd_sc_hd__or3b_1
XFILLER_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15148_ _15262_/C _15270_/B vssd1 vssd1 vccd1 vccd1 _15148_/Y sky130_fd_sc_hd__nand2_1
XFILLER_153_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_966 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15079_ _14898_/Y _15077_/Y _15110_/A vssd1 vssd1 vccd1 vccd1 _15734_/B sky130_fd_sc_hd__o21ai_2
XFILLER_87_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_1001 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09640_ _09640_/A _09795_/A vssd1 vssd1 vccd1 vccd1 _09642_/B sky130_fd_sc_hd__nor2_1
XFILLER_83_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09571_ _10255_/A _10016_/D _09570_/B _09567_/Y vssd1 vssd1 vccd1 vccd1 _09573_/B
+ sky130_fd_sc_hd__a31oi_4
XFILLER_48_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_418 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09005_ _08946_/A _08946_/B _08944_/X vssd1 vssd1 vccd1 vccd1 _09007_/B sky130_fd_sc_hd__a21oi_1
XFILLER_145_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout510 _10638_/A vssd1 vssd1 vccd1 vccd1 _14786_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_59_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout521 _17517_/Q vssd1 vssd1 vccd1 vccd1 _10638_/B sky130_fd_sc_hd__clkbuf_4
Xfanout532 _14842_/A1 vssd1 vssd1 vccd1 vccd1 _14734_/A sky130_fd_sc_hd__clkbuf_4
X_09907_ _09784_/A _09784_/B _09784_/C vssd1 vssd1 vccd1 vccd1 _09908_/B sky130_fd_sc_hd__o21ai_1
Xfanout543 _11122_/A vssd1 vssd1 vccd1 vccd1 _10933_/A sky130_fd_sc_hd__buf_2
Xfanout554 _09899_/B vssd1 vssd1 vccd1 vccd1 _14889_/C sky130_fd_sc_hd__buf_2
Xfanout565 _17164_/A vssd1 vssd1 vccd1 vccd1 _13627_/S sky130_fd_sc_hd__buf_2
XFILLER_101_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout576 fanout578/X vssd1 vssd1 vccd1 vccd1 _11124_/C sky130_fd_sc_hd__buf_2
XFILLER_19_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout587 _11629_/A vssd1 vssd1 vccd1 vccd1 _11561_/A sky130_fd_sc_hd__clkbuf_2
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09838_ _09979_/A _10109_/B _09838_/C _09981_/D vssd1 vssd1 vccd1 vccd1 _09841_/A
+ sky130_fd_sc_hd__and4_1
Xfanout598 _14794_/A vssd1 vssd1 vccd1 vccd1 _10993_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_58_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09769_ _09769_/A _09769_/B _09776_/B _09769_/D vssd1 vssd1 vccd1 vccd1 _09812_/C
+ sky130_fd_sc_hd__and4_1
XTAP_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11800_ _14888_/A _14876_/C _11800_/C _11800_/D vssd1 vssd1 vccd1 vccd1 wire209/A
+ sky130_fd_sc_hd__nor4_1
XTAP_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12780_ _12780_/A _12780_/B vssd1 vssd1 vccd1 vccd1 _12782_/C sky130_fd_sc_hd__xnor2_1
XTAP_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_791 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11731_ _11731_/A _11731_/B _11736_/A vssd1 vssd1 vccd1 vccd1 _11732_/C sky130_fd_sc_hd__nor3_1
XFILLER_26_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_942 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14450_ _16913_/C _14450_/B _14509_/A vssd1 vssd1 vccd1 vccd1 _14567_/A sky130_fd_sc_hd__and3_1
X_11662_ _11662_/A _11662_/B vssd1 vssd1 vccd1 vccd1 _11673_/A sky130_fd_sc_hd__xnor2_1
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13401_ _13526_/B _13401_/B _13401_/C vssd1 vssd1 vccd1 vccd1 _13403_/A sky130_fd_sc_hd__nand3_1
X_10613_ _10613_/A _10613_/B vssd1 vssd1 vccd1 vccd1 _10615_/C sky130_fd_sc_hd__xnor2_1
X_11593_ _11595_/A _14796_/A vssd1 vssd1 vccd1 vccd1 _11593_/Y sky130_fd_sc_hd__nor2_1
X_14381_ _14381_/A _14381_/B vssd1 vssd1 vccd1 vccd1 _14382_/B sky130_fd_sc_hd__nor2_1
XFILLER_128_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16120_ _16108_/C _16114_/A _17075_/A2 _16119_/X vssd1 vssd1 vccd1 vccd1 _16120_/X
+ sky130_fd_sc_hd__a31o_1
X_13332_ _13332_/A _13332_/B _13332_/C vssd1 vssd1 vccd1 vccd1 _13373_/B sky130_fd_sc_hd__and3_1
X_10544_ _10753_/A _12054_/B _10309_/C vssd1 vssd1 vccd1 vccd1 _10544_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_128_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_73 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16051_ _16051_/A _16051_/B vssd1 vssd1 vccd1 vccd1 _16077_/A sky130_fd_sc_hd__xnor2_1
X_10475_ _10385_/A _10385_/C _10385_/B vssd1 vssd1 vccd1 vccd1 _10475_/Y sky130_fd_sc_hd__a21oi_2
X_13263_ _13263_/A _13263_/B vssd1 vssd1 vccd1 vccd1 _13266_/A sky130_fd_sc_hd__nand2_1
XFILLER_157_73 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15002_ _14794_/A _15373_/B _11675_/B vssd1 vssd1 vccd1 vccd1 _15002_/X sky130_fd_sc_hd__a21o_1
X_12214_ _12700_/B _12546_/C vssd1 vssd1 vccd1 vccd1 _12214_/Y sky130_fd_sc_hd__nor2_1
XFILLER_155_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13194_ _13434_/A _13434_/B _13321_/D _13194_/D vssd1 vssd1 vccd1 vccd1 _13195_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_135_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12145_ _12145_/A _12145_/B vssd1 vssd1 vccd1 vccd1 _12146_/B sky130_fd_sc_hd__or2_1
XFILLER_155_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16953_ _16953_/A _16953_/B vssd1 vssd1 vccd1 vccd1 _16955_/A sky130_fd_sc_hd__nor2_1
X_12076_ _12077_/B _12077_/C _12077_/D _12077_/A vssd1 vssd1 vccd1 vccd1 _12078_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_110_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11027_ _11027_/A _11027_/B _11027_/C _11027_/D vssd1 vssd1 vccd1 vccd1 _11032_/A
+ sky130_fd_sc_hd__and4_1
X_15904_ _14924_/A _15457_/B _13516_/X _15900_/Y _15903_/X vssd1 vssd1 vccd1 vccd1
+ _15904_/X sky130_fd_sc_hd__o311a_1
XFILLER_49_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16884_ _16939_/B _16884_/B vssd1 vssd1 vccd1 vccd1 _16886_/B sky130_fd_sc_hd__xnor2_1
XFILLER_49_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15835_ _15836_/B _15836_/A vssd1 vssd1 vccd1 vccd1 _15966_/B sky130_fd_sc_hd__nand2b_1
XFILLER_92_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15766_ _15868_/B _15765_/C _15765_/A vssd1 vssd1 vccd1 vccd1 _15767_/B sky130_fd_sc_hd__o21a_1
X_12978_ _12978_/A _12978_/B vssd1 vssd1 vccd1 vccd1 _12979_/B sky130_fd_sc_hd__and2_1
XTAP_3481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17505_ fanout946/X _17505_/D vssd1 vssd1 vccd1 vccd1 _17505_/Q sky130_fd_sc_hd__dfxtp_4
X_14717_ _14717_/A _14717_/B vssd1 vssd1 vccd1 vccd1 _14718_/B sky130_fd_sc_hd__nand2_1
X_11929_ _11930_/B _12592_/D _12439_/D _17373_/A vssd1 vssd1 vccd1 vccd1 _11931_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_75_1046 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15697_ _15786_/B _15695_/X _15603_/Y _15606_/Y vssd1 vssd1 vccd1 vccd1 _15698_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_162_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17436_ fanout938/X _17436_/D vssd1 vssd1 vccd1 vccd1 _17436_/Q sky130_fd_sc_hd__dfxtp_2
X_14648_ _14765_/A _14738_/B _14679_/B vssd1 vssd1 vccd1 vccd1 _14649_/B sky130_fd_sc_hd__and3_1
XFILLER_162_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_17 _16872_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_28 _17541_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17367_ _17367_/A _17377_/B vssd1 vssd1 vccd1 vccd1 _17367_/Y sky130_fd_sc_hd__nand2_1
XANTENNA_39 _14766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14579_ _14579_/A _14579_/B vssd1 vssd1 vccd1 vccd1 _14580_/B sky130_fd_sc_hd__and2_1
XFILLER_174_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16318_ _16318_/A _16504_/B vssd1 vssd1 vccd1 vccd1 _16321_/A sky130_fd_sc_hd__xnor2_1
XFILLER_146_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17298_ _10062_/B _17308_/A2 _17297_/X _17378_/C1 vssd1 vssd1 vccd1 vccd1 _17478_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_146_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16249_ _16250_/A _16250_/B _16250_/C vssd1 vssd1 vccd1 vccd1 _16251_/A sky130_fd_sc_hd__o21a_1
XFILLER_161_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput102 _17460_/Q vssd1 vssd1 vccd1 vccd1 o_wb_data[26] sky130_fd_sc_hd__clkbuf_1
XFILLER_127_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput113 _17441_/Q vssd1 vssd1 vccd1 vccd1 o_wb_data[7] sky130_fd_sc_hd__clkbuf_1
XFILLER_99_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_1006 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_443 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09623_ _09616_/Y _09621_/X _09629_/A _09601_/Y vssd1 vssd1 vccd1 vccd1 _09629_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_95_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09554_ _17395_/A _09555_/C _09555_/D _09414_/A vssd1 vssd1 vccd1 vccd1 _09556_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_52_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09485_ _09458_/X _09628_/A _09391_/C _09399_/Y vssd1 vssd1 vccd1 vccd1 _09485_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_24_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10260_ _10260_/A _10260_/B vssd1 vssd1 vccd1 vccd1 _10262_/B sky130_fd_sc_hd__xnor2_1
XFILLER_152_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_955 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10191_ _10028_/B _10104_/X _10157_/C _10157_/Y vssd1 vssd1 vccd1 vccd1 _10192_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_160_560 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_20 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout340 _13069_/A vssd1 vssd1 vccd1 vccd1 _11922_/A sky130_fd_sc_hd__buf_2
XFILLER_120_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout351 _17537_/Q vssd1 vssd1 vccd1 vccd1 _14153_/B sky130_fd_sc_hd__clkbuf_4
Xfanout362 _17536_/Q vssd1 vssd1 vccd1 vccd1 _09502_/A sky130_fd_sc_hd__clkbuf_4
X_13950_ _13950_/A _14181_/B vssd1 vssd1 vccd1 vccd1 _13951_/B sky130_fd_sc_hd__nand2_1
XFILLER_47_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout373 _14383_/A vssd1 vssd1 vccd1 vccd1 _13893_/A sky130_fd_sc_hd__buf_2
Xfanout384 _17409_/A vssd1 vssd1 vccd1 vccd1 _09639_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_59_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout395 _17532_/Q vssd1 vssd1 vccd1 vccd1 _14772_/A sky130_fd_sc_hd__buf_6
X_12901_ _12902_/A _12902_/B _12902_/C vssd1 vssd1 vccd1 vccd1 _13065_/A sky130_fd_sc_hd__a21o_1
XFILLER_74_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13881_ _13882_/A _13882_/B vssd1 vssd1 vccd1 vccd1 _13986_/A sky130_fd_sc_hd__and2b_1
XFILLER_19_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_1046 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15620_ _15620_/A _15620_/B vssd1 vssd1 vccd1 vccd1 _15621_/B sky130_fd_sc_hd__and2_1
XFILLER_34_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12832_ _12685_/A _12685_/B _12681_/Y vssd1 vssd1 vccd1 vccd1 _12834_/C sky130_fd_sc_hd__o21ba_1
XTAP_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15551_ _16315_/D _15552_/B vssd1 vssd1 vccd1 vccd1 _15551_/Y sky130_fd_sc_hd__nor2_1
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12763_ _12764_/A _12764_/B _12764_/C vssd1 vssd1 vccd1 vccd1 _12928_/B sky130_fd_sc_hd__a21oi_2
XFILLER_43_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14502_ _14502_/A _14562_/B vssd1 vssd1 vccd1 vccd1 _14505_/A sky130_fd_sc_hd__nand2_1
XTAP_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11714_ _16206_/A _16206_/B vssd1 vssd1 vccd1 vccd1 _16294_/B sky130_fd_sc_hd__and2_1
XTAP_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15482_ _14898_/Y _15077_/Y _16533_/A _15110_/A vssd1 vssd1 vccd1 vccd1 _15567_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_43_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12694_ _12694_/A _12694_/B vssd1 vssd1 vccd1 vccd1 _13003_/A sky130_fd_sc_hd__xnor2_1
XTAP_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17221_ _17441_/Q _17245_/A2 _17219_/X _17220_/X _17275_/C1 vssd1 vssd1 vccd1 vccd1
+ _17441_/D sky130_fd_sc_hd__o221a_1
X_14433_ _14680_/A _14433_/B vssd1 vssd1 vccd1 vccd1 _14492_/A sky130_fd_sc_hd__nand2_4
X_11645_ _11641_/A _11664_/A _11644_/X vssd1 vssd1 vccd1 vccd1 _11646_/C sky130_fd_sc_hd__a21o_1
XFILLER_156_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17152_ _17153_/B _17167_/C vssd1 vssd1 vccd1 vccd1 _17152_/Y sky130_fd_sc_hd__nor2_1
XFILLER_155_310 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput15 i_wb_addr[20] vssd1 vssd1 vccd1 vccd1 input15/X sky130_fd_sc_hd__clkbuf_1
X_14364_ _14364_/A _14364_/B vssd1 vssd1 vccd1 vccd1 _14365_/B sky130_fd_sc_hd__and2_1
XFILLER_168_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11576_ _11576_/A _11576_/B vssd1 vssd1 vccd1 vccd1 _11577_/B sky130_fd_sc_hd__and2_1
Xinput26 i_wb_addr[30] vssd1 vssd1 vccd1 vccd1 input26/X sky130_fd_sc_hd__clkbuf_1
XFILLER_128_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput37 i_wb_data[10] vssd1 vssd1 vccd1 vccd1 input37/X sky130_fd_sc_hd__clkbuf_1
Xinput48 i_wb_data[20] vssd1 vssd1 vccd1 vccd1 input48/X sky130_fd_sc_hd__clkbuf_1
X_16103_ _16100_/B _16101_/Y _16102_/X vssd1 vssd1 vccd1 vccd1 _16103_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_155_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13315_ _13442_/A _13315_/B vssd1 vssd1 vccd1 vccd1 _13317_/C sky130_fd_sc_hd__and2_1
Xinput59 i_wb_data[30] vssd1 vssd1 vccd1 vccd1 input59/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_143_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10527_ _10528_/A _10526_/Y _10970_/A _10786_/B vssd1 vssd1 vccd1 vccd1 _10626_/A
+ sky130_fd_sc_hd__and4bb_1
X_17083_ _17083_/A _17083_/B _17083_/C vssd1 vssd1 vccd1 vccd1 _17085_/C sky130_fd_sc_hd__and3_1
X_14295_ _14372_/B _14295_/B vssd1 vssd1 vccd1 vccd1 _14297_/B sky130_fd_sc_hd__nor2_1
XFILLER_155_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16034_ _16034_/A _16034_/B vssd1 vssd1 vccd1 vccd1 _16035_/B sky130_fd_sc_hd__xnor2_1
XFILLER_109_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13246_ _13246_/A _13246_/B vssd1 vssd1 vccd1 vccd1 _13248_/C sky130_fd_sc_hd__and2_1
XFILLER_108_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10458_ _10459_/A _10459_/B _10459_/C vssd1 vssd1 vccd1 vccd1 _10458_/X sky130_fd_sc_hd__and3_1
XFILLER_124_730 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13177_ _13178_/A _13178_/B _13178_/C vssd1 vssd1 vccd1 vccd1 _13177_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_97_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10389_ _10390_/A _10390_/B _10390_/C vssd1 vssd1 vccd1 vccd1 _10402_/A sky130_fd_sc_hd__a21o_1
XFILLER_112_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12128_ _12128_/A _12343_/A vssd1 vssd1 vccd1 vccd1 _12131_/A sky130_fd_sc_hd__or2_1
XFILLER_69_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16936_ _16935_/A _16935_/B _16935_/C vssd1 vssd1 vccd1 vccd1 _16937_/B sky130_fd_sc_hd__a21oi_1
X_12059_ _14942_/A _15553_/A _12046_/A vssd1 vssd1 vccd1 vccd1 _12397_/B sky130_fd_sc_hd__or3b_1
XFILLER_77_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16867_ _14864_/A _14864_/B _15248_/C vssd1 vssd1 vccd1 vccd1 _16868_/B sky130_fd_sc_hd__o21ai_1
XFILLER_93_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15818_ _16809_/A _16021_/B vssd1 vssd1 vccd1 vccd1 _16497_/D sky130_fd_sc_hd__nand2_1
XFILLER_37_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_577 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16798_ _14863_/B _16652_/B _14863_/A vssd1 vssd1 vccd1 vccd1 _16798_/Y sky130_fd_sc_hd__a21oi_1
X_15749_ _15750_/A _16259_/B vssd1 vssd1 vccd1 vccd1 _15751_/B sky130_fd_sc_hd__nand2_1
XFILLER_80_558 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09270_ _17393_/A _12166_/B vssd1 vssd1 vccd1 vccd1 _16982_/A sky130_fd_sc_hd__nand2_8
XFILLER_61_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17419_ _17419_/A _17421_/B vssd1 vssd1 vccd1 vccd1 _17419_/X sky130_fd_sc_hd__or2_1
XFILLER_20_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_847 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_763 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08985_ _08985_/A _08985_/B _08985_/C vssd1 vssd1 vccd1 vccd1 _09074_/A sky130_fd_sc_hd__or3_1
XFILLER_56_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_544 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_875 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09606_ _09607_/A _09605_/Y _09894_/C _10543_/B vssd1 vssd1 vccd1 vccd1 _09735_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_71_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09537_ _17405_/A _09557_/B _09213_/B _09212_/A vssd1 vssd1 vccd1 vccd1 _09538_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_25_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09468_ _09468_/A _09468_/B vssd1 vssd1 vccd1 vccd1 _09473_/C sky130_fd_sc_hd__nor2_1
XFILLER_12_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_468 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09399_ _09339_/A _09344_/B _09339_/C vssd1 vssd1 vccd1 vccd1 _09399_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_22_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11430_ _11430_/A _11430_/B _11430_/C vssd1 vssd1 vccd1 vccd1 _11475_/A sky130_fd_sc_hd__or3_1
XFILLER_137_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11361_ _11361_/A _11361_/B vssd1 vssd1 vccd1 vccd1 _11411_/A sky130_fd_sc_hd__nand2_1
XFILLER_125_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13100_ _16965_/C _13664_/D vssd1 vssd1 vccd1 vccd1 _13101_/B sky130_fd_sc_hd__nand2_1
X_10312_ _10312_/A _10429_/A vssd1 vssd1 vccd1 vccd1 _10314_/B sky130_fd_sc_hd__nor2_1
XFILLER_152_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11292_ _11293_/A _11293_/B vssd1 vssd1 vccd1 vccd1 _11299_/A sky130_fd_sc_hd__or2_1
X_14080_ _14318_/B _14301_/C _14080_/C vssd1 vssd1 vccd1 vccd1 _14173_/A sky130_fd_sc_hd__and3_1
X_13031_ _13031_/A _13031_/B vssd1 vssd1 vccd1 vccd1 _13033_/C sky130_fd_sc_hd__xnor2_1
X_10243_ _10243_/A _10243_/B vssd1 vssd1 vccd1 vccd1 _10245_/A sky130_fd_sc_hd__nor2_1
XFILLER_65_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10174_ _10174_/A _10174_/B vssd1 vssd1 vccd1 vccd1 _10288_/C sky130_fd_sc_hd__xnor2_1
XFILLER_120_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14982_ _14982_/A _14982_/B _14982_/C vssd1 vssd1 vccd1 vccd1 _14982_/Y sky130_fd_sc_hd__nor3_1
Xfanout170 _16497_/C vssd1 vssd1 vccd1 vccd1 _16662_/C sky130_fd_sc_hd__buf_2
Xfanout181 _16061_/B vssd1 vssd1 vccd1 vccd1 _16589_/B sky130_fd_sc_hd__clkbuf_4
Xfanout192 _15151_/X vssd1 vssd1 vccd1 vccd1 _16136_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_59_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16721_ _16791_/A vssd1 vssd1 vccd1 vccd1 _16721_/Y sky130_fd_sc_hd__inv_2
X_13933_ _13936_/A _13936_/B vssd1 vssd1 vccd1 vccd1 _13935_/B sky130_fd_sc_hd__or2_1
XFILLER_59_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_83 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16652_ _17140_/A _16652_/B _16652_/C vssd1 vssd1 vccd1 vccd1 _16652_/X sky130_fd_sc_hd__or3_1
X_13864_ _13862_/X _13864_/B vssd1 vssd1 vccd1 vccd1 _13870_/A sky130_fd_sc_hd__nand2b_1
XFILLER_34_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_931 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15603_ _15604_/B _15604_/A vssd1 vssd1 vccd1 vccd1 _15603_/Y sky130_fd_sc_hd__nand2b_1
X_12815_ _12816_/A _12816_/B vssd1 vssd1 vccd1 vccd1 _12815_/Y sky130_fd_sc_hd__nand2b_1
X_16583_ _17143_/A1 _14209_/X _16581_/Y _16582_/X vssd1 vssd1 vccd1 vccd1 _16583_/X
+ sky130_fd_sc_hd__o211a_1
X_13795_ _13795_/A _13906_/A vssd1 vssd1 vccd1 vccd1 _13796_/C sky130_fd_sc_hd__and2_1
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15534_ _10716_/A _14785_/X _14806_/X vssd1 vssd1 vccd1 vccd1 _15535_/B sky130_fd_sc_hd__a21o_1
XFILLER_16_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12746_ _12747_/A _12747_/B vssd1 vssd1 vccd1 vccd1 _12920_/A sky130_fd_sc_hd__nand2_1
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15465_ _14806_/A _15804_/A2 _15464_/X vssd1 vssd1 vccd1 vccd1 _15465_/Y sky130_fd_sc_hd__a21oi_1
X_12677_ _12679_/A vssd1 vssd1 vccd1 vccd1 _12677_/Y sky130_fd_sc_hd__inv_2
X_17204_ _17577_/Q _17225_/A2 _17225_/B1 vssd1 vssd1 vccd1 vccd1 _17204_/X sky130_fd_sc_hd__a21o_1
XFILLER_30_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14416_ _14283_/B _14416_/B vssd1 vssd1 vccd1 vccd1 _14534_/A sky130_fd_sc_hd__and2b_1
X_11628_ _11628_/A _11628_/B vssd1 vssd1 vccd1 vccd1 _11635_/A sky130_fd_sc_hd__xnor2_1
X_15396_ _15396_/A _15396_/B _15472_/B vssd1 vssd1 vccd1 vccd1 _16041_/B sky130_fd_sc_hd__nand3_4
XFILLER_156_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17135_ _17133_/Y _17134_/X _17099_/Y _17102_/X vssd1 vssd1 vccd1 vccd1 _17135_/Y
+ sky130_fd_sc_hd__o211ai_1
X_14347_ _14348_/B _14348_/A vssd1 vssd1 vccd1 vccd1 _14413_/B sky130_fd_sc_hd__and2b_1
XFILLER_156_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11559_ _11520_/C _11561_/C _11521_/A _11519_/Y vssd1 vssd1 vccd1 vccd1 _11565_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_128_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17066_ _17066_/A _17066_/B vssd1 vssd1 vccd1 vccd1 _17066_/X sky130_fd_sc_hd__and2_1
XFILLER_170_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14278_ _14278_/A _14278_/B vssd1 vssd1 vccd1 vccd1 _14281_/B sky130_fd_sc_hd__nor2_1
XFILLER_143_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16017_ _16017_/A _16017_/B _16017_/C vssd1 vssd1 vccd1 vccd1 _16017_/X sky130_fd_sc_hd__and3_1
X_13229_ _14155_/A _13764_/D vssd1 vssd1 vccd1 vccd1 _13230_/B sky130_fd_sc_hd__nand2_1
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08770_ _08773_/A vssd1 vssd1 vccd1 vccd1 _08772_/C sky130_fd_sc_hd__inv_2
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_511 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_831 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16919_ _16918_/A _16918_/B _16918_/C vssd1 vssd1 vccd1 vccd1 _16919_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_92_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09322_ _09327_/C _11895_/D _09317_/A _09086_/Y vssd1 vssd1 vccd1 vccd1 _09323_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_09253_ _09250_/Y _09251_/X _09182_/Y _09342_/A vssd1 vssd1 vccd1 vccd1 _09255_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_22_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09184_ _12171_/A _09272_/D vssd1 vssd1 vccd1 vccd1 _09213_/A sky130_fd_sc_hd__nand2_1
XFILLER_147_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08968_ _11839_/S _11815_/B vssd1 vssd1 vccd1 vccd1 _08969_/C sky130_fd_sc_hd__and2_1
XFILLER_112_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08899_ _17389_/A _09042_/B _10297_/D _17391_/A vssd1 vssd1 vccd1 vccd1 _08900_/B
+ sky130_fd_sc_hd__a22oi_1
XFILLER_91_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10930_ _11124_/C _10933_/C _10842_/B _10841_/A vssd1 vssd1 vccd1 vccd1 _10940_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_95_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10861_ _10861_/A _10861_/B _10861_/C vssd1 vssd1 vccd1 vccd1 _10863_/B sky130_fd_sc_hd__and3_1
XFILLER_16_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12600_ _12600_/A _12755_/B vssd1 vssd1 vccd1 vccd1 _12603_/A sky130_fd_sc_hd__nor2_1
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13580_ _13352_/B _13966_/D _13866_/D _14153_/A vssd1 vssd1 vccd1 vccd1 _13582_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_12_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10792_ _10792_/A _10932_/B vssd1 vssd1 vccd1 vccd1 _10884_/A sky130_fd_sc_hd__nand2_1
XPHY_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12531_ _12526_/B _12361_/B _12361_/C _12366_/A vssd1 vssd1 vccd1 vccd1 _12534_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_40_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15250_ _15244_/A _15804_/A2 _15249_/X _14944_/A vssd1 vssd1 vccd1 vccd1 _15250_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_12_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12462_ _12770_/B _12618_/D _12463_/D _12770_/A vssd1 vssd1 vccd1 vccd1 _12464_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_33_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14201_ _14276_/B _14201_/B vssd1 vssd1 vccd1 vccd1 _14202_/C sky130_fd_sc_hd__nand2b_1
X_11413_ _11416_/B _11413_/B _11413_/C vssd1 vssd1 vccd1 vccd1 _11708_/A sky130_fd_sc_hd__nor3_2
XFILLER_138_663 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15181_ _12858_/Y _15180_/B _15179_/X _16011_/A vssd1 vssd1 vccd1 vccd1 _16582_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_165_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12393_ _12865_/S _12393_/B vssd1 vssd1 vccd1 vccd1 _12394_/A sky130_fd_sc_hd__nor2_2
XFILLER_165_471 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14132_ _13951_/B _14042_/Y _13947_/Y vssd1 vssd1 vccd1 vccd1 _14218_/A sky130_fd_sc_hd__a21oi_1
X_11344_ _11352_/A _11352_/B vssd1 vssd1 vccd1 vccd1 _11359_/A sky130_fd_sc_hd__or2_1
XFILLER_126_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14063_ _14153_/A _14153_/B _14063_/C _14213_/C vssd1 vssd1 vccd1 vccd1 _14064_/B
+ sky130_fd_sc_hd__and4_1
X_11275_ _11520_/C _14893_/B _11135_/C vssd1 vssd1 vccd1 vccd1 _11276_/B sky130_fd_sc_hd__a21o_1
XFILLER_4_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13014_ _11805_/X _11810_/X _11838_/X _11843_/X _17367_/A _13516_/S vssd1 vssd1 vccd1
+ vccd1 _13015_/B sky130_fd_sc_hd__mux4_1
XFILLER_140_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10226_ _10226_/A _10226_/B vssd1 vssd1 vccd1 vccd1 _10349_/A sky130_fd_sc_hd__xnor2_1
XFILLER_67_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10157_ _10155_/Y _10157_/B _10157_/C vssd1 vssd1 vccd1 vccd1 _10157_/Y sky130_fd_sc_hd__nand3b_2
XFILLER_58_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10088_ _09959_/X _09972_/Y _10060_/Y _10216_/A vssd1 vssd1 vccd1 vccd1 _10088_/X
+ sky130_fd_sc_hd__o211a_1
X_14965_ _15553_/A _16977_/A _14910_/X _14964_/Y vssd1 vssd1 vccd1 vccd1 _17543_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_75_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16704_ _16705_/A _16705_/B vssd1 vssd1 vccd1 vccd1 _16784_/A sky130_fd_sc_hd__or2_1
X_13916_ _14021_/A _13916_/B vssd1 vssd1 vccd1 vccd1 _13918_/B sky130_fd_sc_hd__nor2_1
XFILLER_63_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14896_ _15208_/A _15381_/A _08731_/A vssd1 vssd1 vccd1 vccd1 _14897_/D sky130_fd_sc_hd__or3b_1
XFILLER_75_694 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16635_ _16636_/A _16636_/B _16636_/C vssd1 vssd1 vccd1 vccd1 _16714_/A sky130_fd_sc_hd__a21oi_1
XFILLER_90_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13847_ _13950_/A _14094_/B _13848_/A vssd1 vssd1 vccd1 vccd1 _13954_/B sky130_fd_sc_hd__and3_1
XFILLER_74_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16566_ _16566_/A _16566_/B vssd1 vssd1 vccd1 vccd1 _16566_/Y sky130_fd_sc_hd__nor2_2
X_13778_ _13778_/A _13778_/B _13778_/C vssd1 vssd1 vccd1 vccd1 _13779_/B sky130_fd_sc_hd__nor3_1
XFILLER_15_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15517_ _15518_/B _15518_/A vssd1 vssd1 vccd1 vccd1 _15609_/B sky130_fd_sc_hd__and2b_1
X_12729_ _12730_/A _12730_/B _12730_/C vssd1 vssd1 vccd1 vccd1 _12902_/A sky130_fd_sc_hd__a21o_1
X_16497_ _16497_/A _16814_/A _16497_/C _16497_/D vssd1 vssd1 vccd1 vccd1 _16609_/A
+ sky130_fd_sc_hd__or4_1
XFILLER_88_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15448_ _15396_/A _15373_/B _15463_/A vssd1 vssd1 vccd1 vccd1 _15532_/A sky130_fd_sc_hd__a21bo_1
XFILLER_30_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_814 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15379_ _10799_/Y _14803_/Y _15456_/B _15378_/X vssd1 vssd1 vccd1 vccd1 _15379_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_129_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17118_ _17118_/A _17118_/B vssd1 vssd1 vccd1 vccd1 _17127_/A sky130_fd_sc_hd__nand2_1
XFILLER_143_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_858 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17049_ _17049_/A _17049_/B vssd1 vssd1 vccd1 vccd1 _17050_/B sky130_fd_sc_hd__nor2_1
X_09940_ _10321_/A _10067_/B _09801_/B _09798_/Y vssd1 vssd1 vccd1 vccd1 _09941_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_171_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout906 _17478_/Q vssd1 vssd1 vccd1 vccd1 _10062_/B sky130_fd_sc_hd__buf_4
XFILLER_135_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout917 _17245_/A2 vssd1 vssd1 vccd1 vccd1 _17275_/A2 sky130_fd_sc_hd__clkbuf_4
X_09871_ _09730_/C _10534_/D _09731_/A _09729_/Y vssd1 vssd1 vccd1 vccd1 _09872_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_112_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout928 _17422_/C1 vssd1 vssd1 vccd1 vccd1 _17406_/C1 sky130_fd_sc_hd__buf_2
XFILLER_98_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout939 fanout940/X vssd1 vssd1 vccd1 vccd1 fanout939/X sky130_fd_sc_hd__buf_2
XFILLER_97_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08822_ _08822_/A _08822_/B vssd1 vssd1 vccd1 vccd1 _08829_/B sky130_fd_sc_hd__xnor2_1
XFILLER_58_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08753_ _17399_/A _11859_/D _09229_/B _17403_/A vssd1 vssd1 vccd1 vccd1 _08754_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_38_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_558 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09305_ _17375_/A _11900_/D _09081_/A _09079_/Y vssd1 vssd1 vccd1 vccd1 _09306_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_139_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09236_ _09236_/A _09236_/B vssd1 vssd1 vccd1 vccd1 _09238_/C sky130_fd_sc_hd__xnor2_1
XFILLER_103_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09167_ _09167_/A _09167_/B vssd1 vssd1 vccd1 vccd1 _09333_/A sky130_fd_sc_hd__or2_1
XFILLER_107_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09098_ _09493_/A _17139_/A _14981_/A vssd1 vssd1 vccd1 vccd1 _09101_/A sky130_fd_sc_hd__and3_1
XFILLER_108_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11060_ _11051_/A _11051_/C _11051_/B vssd1 vssd1 vccd1 vccd1 _11061_/C sky130_fd_sc_hd__a21o_1
XFILLER_89_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10011_ _10271_/A _10036_/D _09876_/A _09874_/Y vssd1 vssd1 vccd1 vccd1 _10018_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_89_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14750_ _14750_/A _14750_/B vssd1 vssd1 vccd1 vccd1 _14751_/B sky130_fd_sc_hd__nand2_1
XFILLER_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11962_ _17407_/A _11961_/B _11961_/C vssd1 vssd1 vccd1 vccd1 _11963_/B sky130_fd_sc_hd__a21o_1
X_13701_ _13702_/A _13702_/B _13702_/C vssd1 vssd1 vccd1 vccd1 _13703_/A sky130_fd_sc_hd__a21oi_1
X_10913_ _10963_/B _11117_/D _11115_/C _10963_/A vssd1 vssd1 vccd1 vccd1 _10914_/B
+ sky130_fd_sc_hd__a22oi_1
XFILLER_17_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14681_ _14682_/A _14682_/B vssd1 vssd1 vccd1 vccd1 _14736_/A sky130_fd_sc_hd__nor2_1
X_11893_ _11890_/X _11891_/Y _08801_/A _08801_/Y vssd1 vssd1 vccd1 vccd1 _11915_/B
+ sky130_fd_sc_hd__o211a_1
X_16420_ _16420_/A vssd1 vssd1 vccd1 vccd1 _16422_/B sky130_fd_sc_hd__inv_2
XFILLER_71_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13632_ _13632_/A _13632_/B _13738_/B _13632_/D vssd1 vssd1 vccd1 vccd1 _13741_/A
+ sky130_fd_sc_hd__and4_1
X_10844_ _10844_/A _10844_/B vssd1 vssd1 vccd1 vccd1 _10846_/B sky130_fd_sc_hd__xnor2_1
XFILLER_71_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16351_ _16619_/A _16681_/C vssd1 vssd1 vccd1 vccd1 _16352_/C sky130_fd_sc_hd__nor2_1
XFILLER_158_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13563_ _13893_/A _13564_/C _13450_/C _14167_/A vssd1 vssd1 vccd1 vccd1 _13565_/A
+ sky130_fd_sc_hd__a22oi_1
X_10775_ _10774_/A _11722_/A _10678_/B _10691_/X vssd1 vssd1 vccd1 vccd1 _10778_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_158_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15302_ _15302_/A _15302_/B vssd1 vssd1 vccd1 vccd1 _15303_/B sky130_fd_sc_hd__or2_1
X_12514_ _12514_/A _12514_/B vssd1 vssd1 vccd1 vccd1 _12515_/B sky130_fd_sc_hd__and2_1
X_16282_ _16282_/A _16282_/B vssd1 vssd1 vccd1 vccd1 _16283_/B sky130_fd_sc_hd__xor2_1
XFILLER_40_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13494_ _13494_/A _13494_/B _13494_/C vssd1 vssd1 vccd1 vccd1 _13495_/B sky130_fd_sc_hd__nor3_1
XFILLER_74_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15233_ _15233_/A _15233_/B vssd1 vssd1 vccd1 vccd1 _15233_/X sky130_fd_sc_hd__or2_1
XFILLER_138_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12445_ _13182_/A _13051_/B _12445_/C _12445_/D vssd1 vssd1 vccd1 vccd1 _12446_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_60_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_622 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15164_ _16086_/A _15164_/B vssd1 vssd1 vccd1 vccd1 _15230_/A sky130_fd_sc_hd__nand2_1
X_12376_ _12015_/Y _12377_/B _12375_/Y _12208_/B vssd1 vssd1 vccd1 vccd1 _13005_/A
+ sky130_fd_sc_hd__o22ai_1
X_14115_ _14115_/A _14115_/B vssd1 vssd1 vccd1 vccd1 _14117_/B sky130_fd_sc_hd__nand2_1
X_11327_ _11331_/B _11327_/B vssd1 vssd1 vccd1 vccd1 _11369_/B sky130_fd_sc_hd__and2_1
XFILLER_126_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15095_ _15097_/A _15095_/B _14979_/B vssd1 vssd1 vccd1 vccd1 _17164_/D sky130_fd_sc_hd__or3b_4
XFILLER_119_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14046_ _14047_/A _14047_/B vssd1 vssd1 vccd1 vccd1 _14150_/A sky130_fd_sc_hd__nor2_1
X_11258_ _15396_/A _15373_/C _11561_/D _11592_/B vssd1 vssd1 vccd1 vccd1 _11261_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_140_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10209_ _10209_/A _10209_/B vssd1 vssd1 vccd1 vccd1 _10210_/B sky130_fd_sc_hd__nor2_1
X_11189_ _11218_/B _11187_/X _11053_/Y _11055_/X vssd1 vssd1 vccd1 vccd1 _11190_/C
+ sky130_fd_sc_hd__a211oi_1
XFILLER_121_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15997_ _15997_/A _15997_/B vssd1 vssd1 vccd1 vccd1 _15998_/B sky130_fd_sc_hd__nor2_1
XFILLER_55_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14948_ _14948_/A _14948_/B _14948_/C vssd1 vssd1 vccd1 vccd1 _14948_/Y sky130_fd_sc_hd__nor3_1
XFILLER_47_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14879_ _15147_/C _17614_/Q vssd1 vssd1 vccd1 vccd1 _14879_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_39_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_804 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16618_ _16695_/A _16533_/B _16695_/B _16533_/A vssd1 vssd1 vccd1 vccd1 _16620_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_126_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17598_ fanout933/X _17598_/D vssd1 vssd1 vccd1 vccd1 _17598_/Q sky130_fd_sc_hd__dfxtp_1
X_16549_ _16550_/A _16550_/B _16550_/C vssd1 vssd1 vccd1 vccd1 _16636_/A sky130_fd_sc_hd__a21o_1
XFILLER_31_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09021_ _17401_/A _12340_/B _08882_/A _08880_/Y vssd1 vssd1 vccd1 vccd1 _09027_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_163_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1020 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09923_ _09923_/A _09923_/B vssd1 vssd1 vccd1 vccd1 _09956_/A sky130_fd_sc_hd__and2_1
Xfanout703 _16654_/B2 vssd1 vssd1 vccd1 vccd1 _16651_/A sky130_fd_sc_hd__clkbuf_4
Xfanout714 _17498_/Q vssd1 vssd1 vccd1 vccd1 _12079_/B sky130_fd_sc_hd__clkbuf_4
Xfanout725 _13866_/C vssd1 vssd1 vccd1 vccd1 _13966_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_86_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout736 _10171_/D vssd1 vssd1 vccd1 vccd1 _16298_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_131_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout747 _10297_/D vssd1 vssd1 vccd1 vccd1 _10993_/D sky130_fd_sc_hd__buf_4
X_09854_ _09854_/A _09854_/B vssd1 vssd1 vccd1 vccd1 _09862_/A sky130_fd_sc_hd__xnor2_1
Xfanout758 _10899_/D vssd1 vssd1 vccd1 vccd1 _10647_/D sky130_fd_sc_hd__clkbuf_4
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout769 _10532_/D vssd1 vssd1 vccd1 vccd1 _10745_/D sky130_fd_sc_hd__buf_2
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08805_ _17403_/A _17399_/A _11961_/B _12340_/B vssd1 vssd1 vccd1 vccd1 _08808_/A
+ sky130_fd_sc_hd__and4_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09785_ _09502_/A _09172_/B _09502_/B _09172_/A vssd1 vssd1 vccd1 vccd1 _09786_/B
+ sky130_fd_sc_hd__a22oi_1
XTAP_3107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_801 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08736_ _17607_/Q _17608_/Q vssd1 vssd1 vccd1 vccd1 _14929_/A sky130_fd_sc_hd__nand2_2
XFILLER_67_992 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_299 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10560_ _10560_/A _10560_/B _11027_/C _11027_/D vssd1 vssd1 vccd1 vccd1 _11749_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_155_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09219_ _09219_/A _11958_/A _09219_/C vssd1 vssd1 vccd1 vccd1 _11958_/B sky130_fd_sc_hd__nor3_1
XFILLER_10_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10491_ _15393_/A _10962_/B vssd1 vssd1 vccd1 vccd1 _10601_/A sky130_fd_sc_hd__nand2_1
XFILLER_108_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12230_ _12710_/A _12230_/B vssd1 vssd1 vccd1 vccd1 _12230_/X sky130_fd_sc_hd__or2_1
XFILLER_107_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12161_ _12161_/A _12325_/A _12161_/C vssd1 vssd1 vccd1 vccd1 _12325_/B sky130_fd_sc_hd__nor3_1
XFILLER_146_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11112_ _11112_/A _11112_/B _11112_/C vssd1 vssd1 vccd1 vccd1 _11146_/A sky130_fd_sc_hd__or3_1
XFILLER_122_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12092_ _12093_/A _12093_/B _12093_/C vssd1 vssd1 vccd1 vccd1 _12286_/A sky130_fd_sc_hd__o21ai_1
XFILLER_151_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11043_ _11043_/A _11043_/B vssd1 vssd1 vccd1 vccd1 _11058_/B sky130_fd_sc_hd__xnor2_1
X_15920_ _16315_/C _16499_/B vssd1 vssd1 vccd1 vccd1 _15921_/B sky130_fd_sc_hd__nor2_1
XFILLER_39_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_756 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15851_ _16446_/A _16667_/A vssd1 vssd1 vccd1 vccd1 _15853_/B sky130_fd_sc_hd__nor2_2
XFILLER_162_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14802_ _14801_/B _14801_/C _11100_/A vssd1 vssd1 vccd1 vccd1 _14803_/B sky130_fd_sc_hd__o21a_1
XFILLER_64_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15782_ _15782_/A _15782_/B vssd1 vssd1 vccd1 vccd1 _15784_/B sky130_fd_sc_hd__nand2_1
XFILLER_149_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12994_ _12993_/A _12993_/B _12991_/X vssd1 vssd1 vccd1 vccd1 _12997_/B sky130_fd_sc_hd__o21ba_1
XFILLER_91_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17521_ fanout943/X _17521_/D vssd1 vssd1 vccd1 vccd1 _17521_/Q sky130_fd_sc_hd__dfxtp_4
X_14733_ _13624_/B _13627_/X _14733_/S vssd1 vssd1 vccd1 vccd1 _14734_/B sky130_fd_sc_hd__mux2_1
X_11945_ _09006_/X _09010_/A _11943_/Y _11944_/X vssd1 vssd1 vccd1 vccd1 _12156_/B
+ sky130_fd_sc_hd__a211o_1
XTAP_2940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17452_ fanout951/X _17452_/D vssd1 vssd1 vccd1 vccd1 _17452_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14664_ _14664_/A _14669_/B vssd1 vssd1 vccd1 vccd1 _14664_/X sky130_fd_sc_hd__or2_1
XTAP_2984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11876_ _11877_/A _11877_/B _11877_/C vssd1 vssd1 vccd1 vccd1 _11891_/A sky130_fd_sc_hd__a21oi_4
XFILLER_33_848 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16403_ _17143_/A1 _14036_/X _16582_/A _15040_/X vssd1 vssd1 vccd1 vccd1 _16404_/C
+ sky130_fd_sc_hd__o22a_1
X_13615_ _13501_/B _13503_/B _13501_/A vssd1 vssd1 vccd1 vccd1 _13618_/B sky130_fd_sc_hd__o21ba_1
X_10827_ _10827_/A _10827_/B vssd1 vssd1 vccd1 vccd1 _10828_/B sky130_fd_sc_hd__nor2_1
X_17383_ _17383_/A _17389_/B vssd1 vssd1 vccd1 vccd1 _17383_/X sky130_fd_sc_hd__or2_1
XFILLER_60_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14595_ _14676_/A _14641_/C vssd1 vssd1 vccd1 vccd1 _14597_/B sky130_fd_sc_hd__and2_2
XFILLER_158_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16334_ _16334_/A _16827_/A _16334_/C _16827_/B vssd1 vssd1 vccd1 vccd1 _16335_/B
+ sky130_fd_sc_hd__or4_1
X_13546_ _13418_/A _13419_/Y _13662_/A _13545_/X vssd1 vssd1 vccd1 vccd1 _13662_/B
+ sky130_fd_sc_hd__a211oi_2
X_10758_ _10757_/A _10757_/B _10757_/C vssd1 vssd1 vccd1 vccd1 _10759_/B sky130_fd_sc_hd__o21ai_1
XFILLER_13_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16265_ _16172_/A _16172_/B _16170_/A vssd1 vssd1 vccd1 vccd1 _16266_/B sky130_fd_sc_hd__o21ai_1
XFILLER_145_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13477_ _13477_/A _13477_/B vssd1 vssd1 vccd1 vccd1 _13479_/B sky130_fd_sc_hd__nor2_1
X_10689_ _10690_/A _10690_/B vssd1 vssd1 vccd1 vccd1 _10689_/X sky130_fd_sc_hd__and2_1
XFILLER_139_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15216_ _15216_/A _15216_/B vssd1 vssd1 vccd1 vccd1 _15218_/B sky130_fd_sc_hd__xor2_1
XFILLER_127_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12428_ _12429_/A _12429_/B _12429_/C vssd1 vssd1 vccd1 vccd1 _12607_/A sky130_fd_sc_hd__o21a_1
X_16196_ _16197_/A _16197_/B _16195_/Y vssd1 vssd1 vccd1 vccd1 _16290_/B sky130_fd_sc_hd__o21ba_1
XFILLER_126_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15147_ _15147_/A _17614_/Q _15147_/C _15147_/D vssd1 vssd1 vccd1 vccd1 _15147_/Y
+ sky130_fd_sc_hd__nor4_1
XFILLER_114_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12359_ _12526_/A _12358_/B _12358_/C vssd1 vssd1 vccd1 vccd1 _12361_/B sky130_fd_sc_hd__a21o_1
XFILLER_5_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15078_ _14898_/Y _15077_/Y _15110_/A vssd1 vssd1 vccd1 vccd1 _15647_/A sky130_fd_sc_hd__o21a_4
XFILLER_45_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14029_ _14030_/A _14030_/B _14030_/C vssd1 vssd1 vccd1 vccd1 _14029_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_68_723 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_1046 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_767 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09570_ _09567_/Y _09570_/B vssd1 vssd1 vccd1 vccd1 _09707_/B sky130_fd_sc_hd__and2b_1
XFILLER_82_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_566 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09004_ _09004_/A _09004_/B vssd1 vssd1 vccd1 vccd1 _09007_/A sky130_fd_sc_hd__xnor2_1
XFILLER_129_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_444 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout500 _17519_/Q vssd1 vssd1 vccd1 vccd1 _12907_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_104_157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout511 _10638_/A vssd1 vssd1 vccd1 vccd1 _11115_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_132_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout522 _09894_/C vssd1 vssd1 vccd1 vccd1 _17375_/A sky130_fd_sc_hd__clkbuf_4
X_09906_ _09906_/A _09906_/B _10035_/A vssd1 vssd1 vccd1 vccd1 _09909_/B sky130_fd_sc_hd__nand3_1
Xfanout533 _14842_/A1 vssd1 vssd1 vccd1 vccd1 _15457_/A sky130_fd_sc_hd__buf_4
XFILLER_116_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout544 _09899_/A vssd1 vssd1 vccd1 vccd1 _11122_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_76_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout555 _09899_/B vssd1 vssd1 vccd1 vccd1 _11553_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_59_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout566 _17112_/A1 vssd1 vssd1 vccd1 vccd1 _17164_/A sky130_fd_sc_hd__clkbuf_2
Xfanout577 fanout578/X vssd1 vssd1 vccd1 vccd1 _10745_/C sky130_fd_sc_hd__clkbuf_2
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09837_ _09842_/A _09842_/B vssd1 vssd1 vccd1 vccd1 _09848_/A sky130_fd_sc_hd__nor2_1
XFILLER_112_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout588 _10991_/A vssd1 vssd1 vccd1 vccd1 _11629_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_100_341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout599 _10792_/A vssd1 vssd1 vccd1 vccd1 _14794_/A sky130_fd_sc_hd__buf_2
XFILLER_101_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09768_ _09768_/A _09768_/B _09832_/A vssd1 vssd1 vccd1 vccd1 _09769_/D sky130_fd_sc_hd__or3_1
XFILLER_73_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08719_ _14421_/S vssd1 vssd1 vccd1 vccd1 _14962_/A sky130_fd_sc_hd__clkinv_2
XFILLER_92_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09699_ _09699_/A _09706_/A vssd1 vssd1 vccd1 vccd1 _09701_/C sky130_fd_sc_hd__nor2_1
XTAP_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_59 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11730_ _11731_/B _11736_/A _11731_/A vssd1 vssd1 vccd1 vccd1 _11732_/B sky130_fd_sc_hd__o21a_1
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11661_ _11662_/A _11662_/B vssd1 vssd1 vccd1 vccd1 _11666_/A sky130_fd_sc_hd__and2b_1
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13400_ _13846_/A _14065_/B _13282_/A _13280_/B vssd1 vssd1 vccd1 vccd1 _13401_/C
+ sky130_fd_sc_hd__a31o_1
X_10612_ _10598_/X _10611_/Y _10499_/Y _10589_/X vssd1 vssd1 vccd1 vccd1 _10632_/A
+ sky130_fd_sc_hd__a211o_2
X_14380_ _14381_/A _14381_/B vssd1 vssd1 vccd1 vccd1 _14382_/A sky130_fd_sc_hd__and2_1
X_11592_ _11629_/A _11592_/B vssd1 vssd1 vccd1 vccd1 _14796_/A sky130_fd_sc_hd__nand2_1
XFILLER_41_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13331_ _13332_/A _13332_/B _13332_/C vssd1 vssd1 vccd1 vccd1 _13494_/A sky130_fd_sc_hd__a21oi_2
X_10543_ _10753_/A _10543_/B _10543_/C vssd1 vssd1 vccd1 vccd1 _10546_/A sky130_fd_sc_hd__and3_1
X_16050_ _16051_/B _16051_/A vssd1 vssd1 vccd1 vccd1 _16183_/A sky130_fd_sc_hd__and2b_1
XFILLER_127_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13262_ _13261_/A _13261_/B _13261_/C vssd1 vssd1 vccd1 vccd1 _13263_/B sky130_fd_sc_hd__a21o_1
XFILLER_109_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10474_ _10405_/B _10405_/C _10405_/D _10405_/A vssd1 vssd1 vccd1 vccd1 _10474_/Y
+ sky130_fd_sc_hd__o22ai_1
X_15001_ _14995_/X _15538_/B _15538_/A vssd1 vssd1 vccd1 vccd1 _15001_/X sky130_fd_sc_hd__mux2_1
XFILLER_157_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_912 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12213_ _12211_/X _12212_/X _12848_/S vssd1 vssd1 vccd1 vccd1 _12213_/X sky130_fd_sc_hd__mux2_1
XFILLER_108_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13193_ _13434_/B _13321_/D _13194_/D _13434_/A vssd1 vssd1 vccd1 vccd1 _13195_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_163_580 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12144_ _12145_/A _12145_/B vssd1 vssd1 vccd1 vccd1 _12146_/A sky130_fd_sc_hd__nand2_1
XFILLER_123_455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16952_ _16952_/A _16952_/B _16952_/C vssd1 vssd1 vccd1 vccd1 _16953_/B sky130_fd_sc_hd__and3_1
X_12075_ _12075_/A _12075_/B vssd1 vssd1 vccd1 vccd1 _12082_/A sky130_fd_sc_hd__xnor2_1
XFILLER_96_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11026_ _11027_/B _11027_/D vssd1 vssd1 vccd1 vccd1 _11058_/A sky130_fd_sc_hd__nand2_1
X_15903_ _17371_/A _15901_/X _15902_/X _15808_/A vssd1 vssd1 vccd1 vccd1 _15903_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_110_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16883_ _16883_/A _16938_/D _16883_/C vssd1 vssd1 vccd1 vccd1 _16884_/B sky130_fd_sc_hd__or3_1
XFILLER_65_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15834_ _15834_/A _15834_/B vssd1 vssd1 vccd1 vccd1 _15836_/B sky130_fd_sc_hd__xnor2_1
XFILLER_37_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15765_ _15765_/A _15868_/B _15765_/C vssd1 vssd1 vccd1 vccd1 _15866_/B sky130_fd_sc_hd__nor3_1
X_12977_ _12976_/A _12976_/B _12975_/X vssd1 vssd1 vccd1 vccd1 _12978_/B sky130_fd_sc_hd__o21bai_1
XTAP_3471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17504_ fanout946/X _17504_/D vssd1 vssd1 vccd1 vccd1 _17504_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_61_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11928_ _11930_/B _12592_/D vssd1 vssd1 vccd1 vccd1 _12470_/B sky130_fd_sc_hd__nand2_1
XFILLER_61_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14716_ _14717_/A _14717_/B vssd1 vssd1 vccd1 vccd1 _14747_/A sky130_fd_sc_hd__or2_1
X_15696_ _15603_/Y _15606_/Y _15786_/B _15695_/X vssd1 vssd1 vccd1 vccd1 _15698_/A
+ sky130_fd_sc_hd__a211oi_1
XTAP_2770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_807 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17435_ fanout940/X _17435_/D vssd1 vssd1 vccd1 vccd1 _17435_/Q sky130_fd_sc_hd__dfxtp_2
X_14647_ _14594_/A _14596_/Y _14594_/B vssd1 vssd1 vccd1 vccd1 _14649_/A sky130_fd_sc_hd__o21bai_2
X_11859_ _12068_/A _12068_/B _12500_/B _11859_/D vssd1 vssd1 vccd1 vccd1 _11860_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_20_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_18 _16873_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_29 _17543_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17366_ input47/X _17377_/B _17365_/Y _17378_/C1 vssd1 vssd1 vccd1 vccd1 _17511_/D
+ sky130_fd_sc_hd__o211a_1
X_14578_ _14579_/A _14579_/B vssd1 vssd1 vccd1 vccd1 _14627_/B sky130_fd_sc_hd__nor2_1
XFILLER_119_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16317_ _16317_/A _16317_/B vssd1 vssd1 vccd1 vccd1 _16504_/B sky130_fd_sc_hd__nand2_1
X_13529_ _13527_/X _13529_/B vssd1 vssd1 vccd1 vccd1 _13535_/A sky130_fd_sc_hd__and2b_1
X_17297_ input36/X _17362_/C _17429_/C vssd1 vssd1 vccd1 vccd1 _17297_/X sky130_fd_sc_hd__or3_1
XFILLER_70_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16248_ _16248_/A _16248_/B vssd1 vssd1 vccd1 vccd1 _16250_/C sky130_fd_sc_hd__nor2_1
XFILLER_146_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput103 _17461_/Q vssd1 vssd1 vccd1 vccd1 o_wb_data[27] sky130_fd_sc_hd__clkbuf_1
X_16179_ _16179_/A _16179_/B vssd1 vssd1 vccd1 vccd1 _16180_/B sky130_fd_sc_hd__nor2_1
Xoutput114 _17442_/Q vssd1 vssd1 vccd1 vccd1 o_wb_data[8] sky130_fd_sc_hd__clkbuf_1
XFILLER_115_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1018 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_907 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09622_ _09629_/A _09601_/Y _09616_/Y _09621_/X vssd1 vssd1 vccd1 vccd1 _09626_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_55_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09553_ _09559_/B _09559_/A vssd1 vssd1 vccd1 vccd1 _09574_/B sky130_fd_sc_hd__and2b_1
XFILLER_71_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09484_ _09484_/A _09484_/B _09484_/C vssd1 vssd1 vccd1 vccd1 _09628_/A sky130_fd_sc_hd__and3_1
XFILLER_24_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_967 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10190_ _10188_/A _10188_/Y _10207_/A _10161_/X vssd1 vssd1 vccd1 vccd1 _10207_/B
+ sky130_fd_sc_hd__a211oi_2
XFILLER_127_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_328 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout330 _14708_/B vssd1 vssd1 vccd1 vccd1 _14641_/B sky130_fd_sc_hd__buf_2
Xfanout341 _17539_/Q vssd1 vssd1 vccd1 vccd1 _13069_/A sky130_fd_sc_hd__buf_4
Xfanout352 _17537_/Q vssd1 vssd1 vccd1 vccd1 _13352_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_143_32 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout363 _14167_/A vssd1 vssd1 vccd1 vccd1 _14318_/A sky130_fd_sc_hd__buf_2
Xfanout374 fanout380/X vssd1 vssd1 vccd1 vccd1 _14383_/A sky130_fd_sc_hd__buf_2
XFILLER_87_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout385 _17409_/A vssd1 vssd1 vccd1 vccd1 _10321_/A sky130_fd_sc_hd__clkbuf_2
X_12900_ _12900_/A _13049_/B vssd1 vssd1 vccd1 vccd1 _12902_/C sky130_fd_sc_hd__nand2_1
XFILLER_4_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout396 _13908_/A vssd1 vssd1 vccd1 vccd1 _14254_/A sky130_fd_sc_hd__buf_2
XFILLER_59_586 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13880_ _13880_/A _13880_/B vssd1 vssd1 vccd1 vccd1 _13882_/B sky130_fd_sc_hd__xnor2_1
XFILLER_47_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12831_ _12991_/A _12829_/Y _12672_/X _12674_/Y vssd1 vssd1 vccd1 vccd1 _12834_/B
+ sky130_fd_sc_hd__o211a_1
XTAP_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15550_ _08731_/A _14888_/B _15262_/B vssd1 vssd1 vccd1 vccd1 _15552_/B sky130_fd_sc_hd__a21bo_1
XFILLER_15_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12762_ _12928_/A _12762_/B vssd1 vssd1 vccd1 vccd1 _12764_/C sky130_fd_sc_hd__or2_1
XFILLER_36_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_634 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14501_ _14500_/B _14501_/B vssd1 vssd1 vccd1 vccd1 _14562_/B sky130_fd_sc_hd__nand2b_1
XTAP_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11713_ _11713_/A _11713_/B vssd1 vssd1 vccd1 vccd1 _16206_/B sky130_fd_sc_hd__xor2_1
XTAP_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15481_ _15481_/A _15481_/B vssd1 vssd1 vccd1 vccd1 _15504_/A sky130_fd_sc_hd__xnor2_1
X_12693_ _12694_/A _12694_/B vssd1 vssd1 vccd1 vccd1 _12693_/X sky130_fd_sc_hd__or2_1
XTAP_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17220_ _17550_/Q _17244_/B vssd1 vssd1 vccd1 vccd1 _17220_/X sky130_fd_sc_hd__and2_1
X_14432_ _14766_/A _14433_/B _14593_/D _14765_/A vssd1 vssd1 vccd1 vccd1 _14432_/X
+ sky130_fd_sc_hd__a22o_1
X_11644_ _11607_/B _11648_/A _11644_/C vssd1 vssd1 vccd1 vccd1 _11644_/X sky130_fd_sc_hd__and3b_1
XFILLER_42_497 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17151_ _17151_/A _17151_/B vssd1 vssd1 vccd1 vccd1 _17167_/C sky130_fd_sc_hd__nand2_1
X_14363_ _14364_/A _14364_/B vssd1 vssd1 vccd1 vccd1 _14440_/B sky130_fd_sc_hd__nor2_1
XFILLER_156_834 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11575_ _11576_/A _11576_/B vssd1 vssd1 vccd1 vccd1 _11582_/A sky130_fd_sc_hd__nor2_1
Xinput16 i_wb_addr[21] vssd1 vssd1 vccd1 vccd1 input16/X sky130_fd_sc_hd__clkbuf_1
XFILLER_155_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput27 i_wb_addr[31] vssd1 vssd1 vccd1 vccd1 input27/X sky130_fd_sc_hd__clkbuf_1
XFILLER_11_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16102_ _15991_/X _15994_/X _16100_/Y _16911_/A vssd1 vssd1 vccd1 vccd1 _16102_/X
+ sky130_fd_sc_hd__o31a_1
X_13314_ _13314_/A _13314_/B _13314_/C vssd1 vssd1 vccd1 vccd1 _13315_/B sky130_fd_sc_hd__or3_1
Xinput38 i_wb_data[11] vssd1 vssd1 vccd1 vccd1 input38/X sky130_fd_sc_hd__clkbuf_1
X_10526_ _10638_/B _10743_/D _10933_/D _10638_/A vssd1 vssd1 vccd1 vccd1 _10526_/Y
+ sky130_fd_sc_hd__a22oi_1
X_17082_ _09412_/A _10897_/B _17038_/B _11006_/A _10899_/D vssd1 vssd1 vccd1 vccd1
+ _17083_/C sky130_fd_sc_hd__a32o_1
Xinput49 i_wb_data[21] vssd1 vssd1 vccd1 vccd1 input49/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14294_ _14294_/A _14294_/B vssd1 vssd1 vccd1 vccd1 _14295_/B sky130_fd_sc_hd__and2_1
XFILLER_143_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16033_ _16136_/B _16591_/B vssd1 vssd1 vccd1 vccd1 _16034_/B sky130_fd_sc_hd__nand2_1
XFILLER_6_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13245_ _13244_/B _13244_/C _13244_/A vssd1 vssd1 vccd1 vccd1 _13246_/B sky130_fd_sc_hd__a21o_1
XFILLER_143_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10457_ _10319_/Y _10354_/X _10407_/Y _10442_/Y vssd1 vssd1 vccd1 vccd1 _10459_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_124_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13176_ _13176_/A _13176_/B vssd1 vssd1 vccd1 vccd1 _13178_/C sky130_fd_sc_hd__xnor2_1
X_10388_ _10388_/A _10388_/B vssd1 vssd1 vccd1 vccd1 _10390_/C sky130_fd_sc_hd__or2_1
XFILLER_151_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12127_ _17425_/A _17423_/A _12127_/C _12127_/D vssd1 vssd1 vccd1 vccd1 _12343_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_97_637 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1002 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16935_ _16935_/A _16935_/B _16935_/C vssd1 vssd1 vccd1 vccd1 _16937_/A sky130_fd_sc_hd__and3_1
X_12058_ _12038_/X _12057_/X _14356_/S vssd1 vssd1 vccd1 vccd1 _12058_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11009_ _11009_/A _11009_/B vssd1 vssd1 vccd1 vccd1 _11025_/A sky130_fd_sc_hd__xor2_1
XFILLER_42_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16866_ _16866_/A _16866_/B vssd1 vssd1 vccd1 vccd1 _16866_/Y sky130_fd_sc_hd__nand2_1
X_15817_ _16809_/A _17083_/A vssd1 vssd1 vccd1 vccd1 _16987_/B sky130_fd_sc_hd__and2_1
XFILLER_65_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16797_ _16797_/A _16797_/B vssd1 vssd1 vccd1 vccd1 _16797_/X sky130_fd_sc_hd__xor2_1
XFILLER_19_995 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15748_ _15414_/B _15746_/X _15747_/X vssd1 vssd1 vccd1 vccd1 _15751_/A sky130_fd_sc_hd__o21a_1
XFILLER_34_954 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15679_ _15679_/A _15772_/B _15679_/C vssd1 vssd1 vccd1 vccd1 _15769_/B sky130_fd_sc_hd__and3_1
X_17418_ input55/X _17424_/A2 _17417_/X _17420_/C1 vssd1 vssd1 vccd1 vccd1 _17537_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_20_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17349_ input54/X _17353_/B _17353_/C vssd1 vssd1 vccd1 vccd1 _17349_/X sky130_fd_sc_hd__or3_1
XFILLER_174_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_506 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08984_ _09242_/B _08984_/B vssd1 vssd1 vccd1 vccd1 _08985_/C sky130_fd_sc_hd__nand2_1
XFILLER_102_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09605_ _09892_/B _10545_/D _10299_/D _09892_/A vssd1 vssd1 vccd1 vccd1 _09605_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_56_567 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_28 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09536_ _09536_/A _09536_/B vssd1 vssd1 vccd1 vccd1 _09538_/A sky130_fd_sc_hd__nor2_1
XFILLER_83_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09467_ _09327_/C _11808_/B _09462_/A _09326_/Y vssd1 vssd1 vccd1 vccd1 _09468_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_25_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09398_ _09393_/B _09393_/C _09393_/D _09395_/B vssd1 vssd1 vccd1 vccd1 _09398_/Y
+ sky130_fd_sc_hd__o22ai_1
XFILLER_40_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11360_ _11354_/A _11354_/C _11354_/B vssd1 vssd1 vccd1 vccd1 _11361_/B sky130_fd_sc_hd__o21ai_1
XFILLER_164_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10311_ _10312_/A _10310_/Y _14954_/A _10311_/D vssd1 vssd1 vccd1 vccd1 _10429_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_138_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11291_ _11291_/A _11291_/B vssd1 vssd1 vccd1 vccd1 _11293_/B sky130_fd_sc_hd__and2_1
XFILLER_152_336 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13030_ _13031_/A _13031_/B vssd1 vssd1 vccd1 vccd1 _13165_/B sky130_fd_sc_hd__nand2_1
X_10242_ _10242_/A1 _10359_/B _10479_/B _10591_/A vssd1 vssd1 vccd1 vccd1 _10243_/B
+ sky130_fd_sc_hd__a22oi_1
XFILLER_133_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10173_ _10288_/A _10172_/Y _15805_/A _10545_/D vssd1 vssd1 vccd1 vccd1 _10296_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_121_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_767 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout160 _17425_/B vssd1 vssd1 vccd1 vccd1 _17421_/B sky130_fd_sc_hd__clkbuf_2
X_14981_ _14981_/A _14981_/B vssd1 vssd1 vccd1 vccd1 _14981_/Y sky130_fd_sc_hd__nor2_1
Xfanout171 _15724_/X vssd1 vssd1 vccd1 vccd1 _16743_/C sky130_fd_sc_hd__buf_2
XFILLER_59_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout182 _15472_/Y vssd1 vssd1 vccd1 vccd1 _16827_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_120_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16720_ _16723_/A _16965_/B _16722_/A vssd1 vssd1 vccd1 vccd1 _16791_/A sky130_fd_sc_hd__a21bo_1
Xfanout193 _15145_/X vssd1 vssd1 vccd1 vccd1 _15493_/A sky130_fd_sc_hd__buf_2
X_13932_ _13932_/A _13932_/B vssd1 vssd1 vccd1 vccd1 _14122_/A sky130_fd_sc_hd__xnor2_1
XFILLER_19_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13863_ _13964_/A _13862_/C _13862_/A vssd1 vssd1 vccd1 vccd1 _13864_/B sky130_fd_sc_hd__a21o_1
XFILLER_47_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16651_ _16651_/A _16651_/B vssd1 vssd1 vccd1 vccd1 _16652_/C sky130_fd_sc_hd__nor2_1
XFILLER_35_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12814_ _12976_/A _12976_/B vssd1 vssd1 vccd1 vccd1 _12816_/B sky130_fd_sc_hd__xor2_1
XFILLER_62_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15602_ _15505_/A _15505_/B _15511_/X vssd1 vssd1 vccd1 vccd1 _15604_/B sky130_fd_sc_hd__a21oi_1
XFILLER_16_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13794_ _13793_/A _13793_/B _13793_/C vssd1 vssd1 vccd1 vccd1 _13906_/A sky130_fd_sc_hd__o21ai_1
X_16582_ _16582_/A _16582_/B vssd1 vssd1 vccd1 vccd1 _16582_/X sky130_fd_sc_hd__or2_1
XFILLER_103_90 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12745_ _12585_/B _12585_/C _12585_/A vssd1 vssd1 vccd1 vccd1 _12747_/B sky130_fd_sc_hd__a21bo_1
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15533_ _15533_/A _15533_/B vssd1 vssd1 vccd1 vccd1 _15533_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_42_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_609 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15464_ _14805_/B _14928_/Y _15713_/B1 _15463_/A _16869_/C1 vssd1 vssd1 vccd1 vccd1
+ _15464_/X sky130_fd_sc_hd__a221o_1
X_12676_ _12676_/A _12676_/B _12676_/C vssd1 vssd1 vccd1 vccd1 _12679_/A sky130_fd_sc_hd__or3_1
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14415_ _14352_/A _14349_/X _14351_/B vssd1 vssd1 vccd1 vccd1 _14415_/X sky130_fd_sc_hd__o21a_1
X_17203_ _17435_/Q _17245_/A2 _17201_/X _17202_/X _17364_/C1 vssd1 vssd1 vccd1 vccd1
+ _17435_/D sky130_fd_sc_hd__o221a_1
X_11627_ _11613_/A _11612_/B _11612_/C vssd1 vssd1 vccd1 vccd1 _11646_/B sky130_fd_sc_hd__a21o_1
XFILLER_30_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15395_ _15396_/A _15396_/B _15472_/B vssd1 vssd1 vccd1 vccd1 _16606_/B sky130_fd_sc_hd__and3_1
X_14346_ _14254_/A _14450_/B _14255_/A _14253_/A vssd1 vssd1 vccd1 vccd1 _14348_/B
+ sky130_fd_sc_hd__a31oi_1
X_17134_ _17134_/A _17134_/B _17134_/C vssd1 vssd1 vccd1 vccd1 _17134_/X sky130_fd_sc_hd__and3_1
X_11558_ _11558_/A _11558_/B _11558_/C vssd1 vssd1 vccd1 vccd1 _11568_/A sky130_fd_sc_hd__nand3_1
XFILLER_10_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10509_ _10509_/A _10617_/A vssd1 vssd1 vccd1 vccd1 _10511_/B sky130_fd_sc_hd__nor2_1
X_17065_ _17065_/A _17153_/B _14765_/A vssd1 vssd1 vccd1 vccd1 _17065_/X sky130_fd_sc_hd__or3b_1
X_14277_ _14352_/A _14277_/B vssd1 vssd1 vccd1 vccd1 _14283_/B sky130_fd_sc_hd__nand2b_1
X_11489_ _11496_/A _11496_/B vssd1 vssd1 vccd1 vccd1 _11502_/A sky130_fd_sc_hd__or2_1
XFILLER_6_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16016_ _16111_/A _16004_/Y _16007_/X _16015_/X vssd1 vssd1 vccd1 vccd1 _16017_/C
+ sky130_fd_sc_hd__o211a_1
X_13228_ _13228_/A _13228_/B vssd1 vssd1 vccd1 vccd1 _13230_/A sky130_fd_sc_hd__nor2_1
XFILLER_143_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13159_ _13159_/A _13159_/B vssd1 vssd1 vccd1 vccd1 _13161_/B sky130_fd_sc_hd__xnor2_1
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16918_ _16918_/A _16918_/B _16918_/C vssd1 vssd1 vccd1 vccd1 _16918_/X sky130_fd_sc_hd__and3_1
XFILLER_66_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16849_ _16850_/A _16850_/B vssd1 vssd1 vccd1 vccd1 _16851_/A sky130_fd_sc_hd__nand2_1
XFILLER_93_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09321_ _09328_/A _09320_/Y _09321_/C _09321_/D vssd1 vssd1 vccd1 vccd1 _09451_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_22_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09252_ _09182_/Y _09342_/A _09250_/Y _09251_/X vssd1 vssd1 vccd1 vccd1 _09255_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_21_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09183_ _09155_/Y _09156_/X _09179_/A _09346_/A vssd1 vssd1 vccd1 vccd1 _09214_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_146_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_391 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08967_ _11839_/S _08967_/B vssd1 vssd1 vccd1 vccd1 _12700_/C sky130_fd_sc_hd__and2_2
XFILLER_130_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_1041 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08898_ _17387_/A _09446_/D vssd1 vssd1 vccd1 vccd1 _09037_/A sky130_fd_sc_hd__nand2_1
XFILLER_56_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_707 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10860_ _10860_/A _10860_/B vssd1 vssd1 vccd1 vccd1 _10861_/C sky130_fd_sc_hd__xnor2_1
XFILLER_17_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09519_ _09519_/A _09519_/B vssd1 vssd1 vccd1 vccd1 _09520_/C sky130_fd_sc_hd__xnor2_1
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10791_ _11629_/A _11132_/B _10897_/B _10933_/C vssd1 vssd1 vccd1 vccd1 _10794_/A
+ sky130_fd_sc_hd__and4_1
XPHY_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12530_ _12530_/A _12530_/B vssd1 vssd1 vccd1 vccd1 _12534_/A sky130_fd_sc_hd__or2_1
XFILLER_24_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12461_ _12307_/A _12307_/B _12306_/A vssd1 vssd1 vccd1 vccd1 _12478_/A sky130_fd_sc_hd__a21o_1
XFILLER_138_620 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14200_ _14200_/A _14200_/B _14198_/X vssd1 vssd1 vccd1 vccd1 _14201_/B sky130_fd_sc_hd__or3b_1
X_11412_ _11419_/A _11419_/B _11410_/Y vssd1 vssd1 vccd1 vccd1 _11413_/C sky130_fd_sc_hd__a21oi_1
XFILLER_149_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15180_ _16011_/B _15180_/B vssd1 vssd1 vccd1 vccd1 _15180_/X sky130_fd_sc_hd__or2_1
XFILLER_166_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12392_ _12035_/C _12033_/Y _12700_/B vssd1 vssd1 vccd1 vccd1 _12393_/B sky130_fd_sc_hd__mux2_1
XFILLER_138_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14131_ _14131_/A vssd1 vssd1 vccd1 vccd1 _14138_/A sky130_fd_sc_hd__inv_2
X_11343_ _11343_/A _11349_/A vssd1 vssd1 vccd1 vccd1 _11352_/B sky130_fd_sc_hd__and2_1
XFILLER_165_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14062_ _14153_/B _14063_/C _14213_/C _14153_/A vssd1 vssd1 vccd1 vccd1 _14064_/A
+ sky130_fd_sc_hd__a22oi_1
X_11274_ _11274_/A _11274_/B _11274_/C vssd1 vssd1 vccd1 vccd1 _11285_/B sky130_fd_sc_hd__nand3_1
XFILLER_98_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_166 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13013_ _12710_/A _13012_/X _16653_/A vssd1 vssd1 vccd1 vccd1 _13013_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_79_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10225_ _10348_/A _10348_/B _10348_/C vssd1 vssd1 vccd1 vccd1 _11775_/A sky130_fd_sc_hd__o21ai_1
XFILLER_133_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_916 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10156_ _10005_/X _10105_/Y _10134_/A _10134_/Y vssd1 vssd1 vccd1 vccd1 _10157_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_121_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_8 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10087_ _10060_/Y _10216_/A _09959_/X _09972_/Y vssd1 vssd1 vccd1 vccd1 _10090_/A
+ sky130_fd_sc_hd__a211oi_2
X_14964_ _14961_/X _14963_/X _14927_/X _14945_/X vssd1 vssd1 vccd1 vccd1 _14964_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_75_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16703_ _16628_/A _16628_/B _16617_/A vssd1 vssd1 vccd1 vccd1 _16705_/B sky130_fd_sc_hd__a21oi_1
X_13915_ _13915_/A _13915_/B _13915_/C vssd1 vssd1 vccd1 vccd1 _13916_/B sky130_fd_sc_hd__nor3_1
XFILLER_75_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14895_ _15208_/A _14895_/B vssd1 vssd1 vccd1 vccd1 _14905_/C sky130_fd_sc_hd__or2_1
XFILLER_63_846 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16634_ _16634_/A _16634_/B vssd1 vssd1 vccd1 vccd1 _16636_/C sky130_fd_sc_hd__xnor2_1
XFILLER_90_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13846_ _13846_/A _13846_/B vssd1 vssd1 vccd1 vccd1 _13848_/B sky130_fd_sc_hd__nand2_1
XFILLER_74_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16565_ _16203_/X _16293_/A _16561_/X _16562_/Y _16564_/Y vssd1 vssd1 vccd1 vccd1
+ _16566_/B sky130_fd_sc_hd__o311a_2
X_13777_ _13778_/A _13778_/B _13778_/C vssd1 vssd1 vccd1 vccd1 _13779_/A sky130_fd_sc_hd__o21a_1
X_10989_ _10990_/A _10990_/B _10990_/C vssd1 vssd1 vccd1 vccd1 _10999_/A sky130_fd_sc_hd__a21o_1
XFILLER_43_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15516_ _16281_/A _16505_/A _15431_/A _15428_/X vssd1 vssd1 vccd1 vccd1 _15518_/B
+ sky130_fd_sc_hd__a31oi_2
X_12728_ _12886_/B _12728_/B vssd1 vssd1 vccd1 vccd1 _12730_/C sky130_fd_sc_hd__or2_1
XFILLER_31_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16496_ _16334_/A _16497_/C _16497_/D _16497_/A vssd1 vssd1 vccd1 vccd1 _16498_/A
+ sky130_fd_sc_hd__o22ai_1
XFILLER_148_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15447_ _15447_/A _16207_/B vssd1 vssd1 vccd1 vccd1 _15447_/X sky130_fd_sc_hd__or2_1
X_12659_ _17415_/A _13321_/D vssd1 vssd1 vccd1 vccd1 _12660_/B sky130_fd_sc_hd__nand2_1
XFILLER_157_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15378_ _10800_/C _14803_/A _14803_/B vssd1 vssd1 vccd1 vccd1 _15378_/X sky130_fd_sc_hd__o21a_1
XFILLER_117_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17117_ _17096_/A _17096_/B _17093_/Y _17095_/B vssd1 vssd1 vccd1 vccd1 _17130_/A
+ sky130_fd_sc_hd__o31a_1
X_14329_ _14330_/A _14330_/B _14330_/C vssd1 vssd1 vccd1 vccd1 _14409_/A sky130_fd_sc_hd__a21oi_1
XFILLER_144_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17048_ _17049_/A _17049_/B vssd1 vssd1 vccd1 vccd1 _17088_/B sky130_fd_sc_hd__and2_1
XFILLER_98_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09870_ _09870_/A _09870_/B _09870_/C vssd1 vssd1 vccd1 vccd1 _09870_/Y sky130_fd_sc_hd__nand3_1
Xfanout907 _11095_/D vssd1 vssd1 vccd1 vccd1 _15008_/B sky130_fd_sc_hd__clkbuf_4
Xfanout918 _17293_/A2 vssd1 vssd1 vccd1 vccd1 _17290_/A2 sky130_fd_sc_hd__buf_2
XFILLER_97_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout929 _17420_/C1 vssd1 vssd1 vccd1 vccd1 _17422_/C1 sky130_fd_sc_hd__buf_2
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08821_ _08821_/A _08822_/A _08821_/C vssd1 vssd1 vccd1 vccd1 _08869_/A sky130_fd_sc_hd__or3_1
XFILLER_98_776 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_553 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08752_ _08755_/A vssd1 vssd1 vccd1 vccd1 _08754_/C sky130_fd_sc_hd__inv_2
XFILLER_39_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09304_ _09304_/A _09304_/B vssd1 vssd1 vccd1 vccd1 _09438_/A sky130_fd_sc_hd__xnor2_1
XFILLER_62_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09235_ _17415_/A _12174_/D vssd1 vssd1 vccd1 vccd1 _09236_/B sky130_fd_sc_hd__nand2_1
XFILLER_21_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09166_ _11922_/A _09172_/B _09502_/B _08988_/B vssd1 vssd1 vccd1 vccd1 _09167_/B
+ sky130_fd_sc_hd__a22oi_1
XFILLER_119_34 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09097_ _11839_/S _17139_/A vssd1 vssd1 vccd1 vccd1 _14978_/A sky130_fd_sc_hd__and2_1
XFILLER_119_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10010_ _10010_/A _10010_/B vssd1 vssd1 vccd1 vccd1 _10023_/A sky130_fd_sc_hd__nand2_1
XFILLER_88_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09999_ _10126_/B _10270_/B _10255_/B _10254_/A vssd1 vssd1 vccd1 vccd1 _10000_/B
+ sky130_fd_sc_hd__a22oi_1
XFILLER_92_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11961_ _17407_/A _11961_/B _11961_/C vssd1 vssd1 vccd1 vccd1 _12169_/B sky130_fd_sc_hd__nand3_1
XFILLER_57_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_418 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10912_ _10963_/A _10963_/B _11117_/D _11115_/C vssd1 vssd1 vccd1 vccd1 _10914_/A
+ sky130_fd_sc_hd__and4_1
X_13700_ _13800_/B _13700_/B vssd1 vssd1 vccd1 vccd1 _13702_/C sky130_fd_sc_hd__nand2_1
XFILLER_72_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14680_ _14680_/A _14738_/B _14680_/C vssd1 vssd1 vccd1 vccd1 _14682_/B sky130_fd_sc_hd__nand3_1
X_11892_ _08801_/A _08801_/Y _11890_/X _11891_/Y vssd1 vssd1 vccd1 vccd1 _11915_/A
+ sky130_fd_sc_hd__a211oi_4
XFILLER_56_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13631_ _13632_/B _13738_/B _13632_/D _13735_/A vssd1 vssd1 vccd1 vccd1 _13635_/A
+ sky130_fd_sc_hd__a22oi_2
X_10843_ _10844_/A _10844_/B vssd1 vssd1 vccd1 vccd1 _10943_/A sky130_fd_sc_hd__nand2b_1
XFILLER_44_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16350_ _16252_/A _16252_/B _16251_/A vssd1 vssd1 vccd1 vccd1 _16362_/A sky130_fd_sc_hd__a21o_1
X_13562_ _13562_/A _13562_/B vssd1 vssd1 vccd1 vccd1 _13605_/A sky130_fd_sc_hd__nor2_1
XFILLER_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10774_ _10774_/A _10774_/B _10774_/C vssd1 vssd1 vccd1 vccd1 _11722_/A sky130_fd_sc_hd__nor3_1
XFILLER_12_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12513_ _12514_/A _12514_/B vssd1 vssd1 vccd1 vccd1 _12670_/A sky130_fd_sc_hd__nor2_1
X_15301_ _15233_/X _15299_/Y _15300_/Y vssd1 vssd1 vccd1 vccd1 _15301_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_157_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16281_ _16281_/A _16695_/B vssd1 vssd1 vccd1 vccd1 _16282_/B sky130_fd_sc_hd__nand2_1
X_13493_ _13494_/A _13494_/B _13494_/C vssd1 vssd1 vccd1 vccd1 _13495_/A sky130_fd_sc_hd__o21a_1
XFILLER_13_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12444_ _12275_/B _12445_/C _12445_/D _12275_/A vssd1 vssd1 vccd1 vccd1 _12446_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_60_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15232_ _15171_/A _15171_/B _15168_/Y vssd1 vssd1 vccd1 vccd1 _15233_/B sky130_fd_sc_hd__a21boi_1
XFILLER_173_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15163_ _16226_/B _16086_/A _15164_/B vssd1 vssd1 vccd1 vccd1 _15165_/A sky130_fd_sc_hd__a21o_1
XFILLER_126_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12375_ _12375_/A _12375_/B vssd1 vssd1 vccd1 vccd1 _12375_/Y sky130_fd_sc_hd__nor2_1
XFILLER_126_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14114_ _14202_/A _14114_/B vssd1 vssd1 vccd1 vccd1 _14117_/A sky130_fd_sc_hd__nand2_1
XFILLER_114_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11326_ _11320_/A _11320_/C _11320_/B vssd1 vssd1 vccd1 vccd1 _11327_/B sky130_fd_sc_hd__o21ai_1
XFILLER_153_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15094_ _15094_/A _15170_/C vssd1 vssd1 vccd1 vccd1 _15094_/X sky130_fd_sc_hd__xor2_1
XFILLER_141_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14045_ _14134_/B _14045_/B vssd1 vssd1 vccd1 vccd1 _14047_/B sky130_fd_sc_hd__xnor2_1
X_11257_ _11257_/A _11257_/B vssd1 vssd1 vccd1 vccd1 _11274_/A sky130_fd_sc_hd__xnor2_1
XFILLER_140_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10208_ _10208_/A _10208_/B vssd1 vssd1 vccd1 vccd1 _10209_/B sky130_fd_sc_hd__and2_1
XFILLER_95_702 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11188_ _11053_/Y _11055_/X _11218_/B _11187_/X vssd1 vssd1 vccd1 vccd1 _11222_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_122_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10139_ _10271_/A _10016_/D _10017_/A _10015_/Y vssd1 vssd1 vccd1 vccd1 _10140_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_48_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15996_ _15994_/A _15993_/X _15995_/Y vssd1 vssd1 vccd1 vccd1 _15996_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_48_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14947_ _15131_/A _14947_/B vssd1 vssd1 vccd1 vccd1 _15180_/B sky130_fd_sc_hd__nand2_1
XFILLER_76_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14878_ _15147_/C _14888_/B _14877_/Y vssd1 vssd1 vccd1 vccd1 _14878_/X sky130_fd_sc_hd__a21o_1
XFILLER_63_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_816 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16617_ _16617_/A _16617_/B vssd1 vssd1 vccd1 vccd1 _16628_/A sky130_fd_sc_hd__nor2_1
XFILLER_63_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13829_ _13936_/B _13830_/B vssd1 vssd1 vccd1 vccd1 _13829_/Y sky130_fd_sc_hd__nand2_1
XFILLER_23_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17597_ fanout936/X _17597_/D vssd1 vssd1 vccd1 vccd1 _17597_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16548_ _16630_/B _16548_/B vssd1 vssd1 vccd1 vccd1 _16550_/C sky130_fd_sc_hd__nand2_1
XFILLER_148_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_759 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16479_ _14775_/A _16644_/B _16480_/A vssd1 vssd1 vccd1 vccd1 _16481_/A sky130_fd_sc_hd__a21bo_1
X_09020_ _09020_/A _09020_/B vssd1 vssd1 vccd1 vccd1 _09048_/A sky130_fd_sc_hd__xnor2_1
XFILLER_117_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1043 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09922_ _09922_/A _09922_/B vssd1 vssd1 vccd1 vccd1 _09923_/B sky130_fd_sc_hd__or2_1
XFILLER_160_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout704 _17499_/Q vssd1 vssd1 vccd1 vccd1 _16654_/B2 sky130_fd_sc_hd__buf_4
Xfanout715 _10308_/B vssd1 vssd1 vccd1 vccd1 _10543_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_131_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout726 _13866_/C vssd1 vssd1 vccd1 vccd1 _13208_/C sky130_fd_sc_hd__buf_4
XFILLER_131_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout737 _11867_/D vssd1 vssd1 vccd1 vccd1 _09042_/B sky130_fd_sc_hd__clkbuf_4
X_09853_ _09854_/A _09854_/B vssd1 vssd1 vccd1 vccd1 _09870_/A sky130_fd_sc_hd__nand2b_1
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout748 _14859_/B vssd1 vssd1 vccd1 vccd1 _10297_/D sky130_fd_sc_hd__clkbuf_8
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout759 _10036_/D vssd1 vssd1 vccd1 vccd1 _10899_/D sky130_fd_sc_hd__buf_6
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08804_ _08804_/A _08804_/B vssd1 vssd1 vccd1 vccd1 _08815_/A sky130_fd_sc_hd__nor2_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09784_ _09784_/A _09784_/B _09784_/C vssd1 vssd1 vccd1 vccd1 _09932_/A sky130_fd_sc_hd__or3_1
XFILLER_100_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08735_ _17613_/Q _14836_/B _17131_/A vssd1 vssd1 vccd1 vccd1 _17613_/D sky130_fd_sc_hd__mux2_1
XFILLER_22_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_952 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_8 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_28 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_567 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09218_ _09219_/A _11958_/A _09219_/C vssd1 vssd1 vccd1 vccd1 _09220_/A sky130_fd_sc_hd__o21a_1
XFILLER_10_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10490_ _10954_/A _11006_/B _14849_/A _10703_/B vssd1 vssd1 vccd1 vccd1 _10493_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_5_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09149_ _09150_/A _09150_/B vssd1 vssd1 vccd1 vccd1 _09245_/B sky130_fd_sc_hd__nand2b_1
XFILLER_108_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12160_ _12161_/A _12325_/A _12161_/C vssd1 vssd1 vccd1 vccd1 _12162_/A sky130_fd_sc_hd__o21a_1
XFILLER_162_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11111_ _10893_/A _10893_/B _10893_/C vssd1 vssd1 vccd1 vccd1 _11112_/C sky130_fd_sc_hd__a21oi_1
XFILLER_1_411 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12091_ _12091_/A _12091_/B vssd1 vssd1 vccd1 vccd1 _12093_/C sky130_fd_sc_hd__xnor2_1
XFILLER_89_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11042_ _11041_/A _11041_/B _11041_/C vssd1 vssd1 vccd1 vccd1 _11042_/X sky130_fd_sc_hd__a21o_1
XFILLER_39_30 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15850_ _15850_/A _15850_/B vssd1 vssd1 vccd1 vccd1 _15859_/A sky130_fd_sc_hd__xor2_1
XFILLER_76_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14801_ _14801_/A _14801_/B _14801_/C vssd1 vssd1 vccd1 vccd1 _14801_/X sky130_fd_sc_hd__or3_1
XFILLER_18_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15781_ _15781_/A _15781_/B vssd1 vssd1 vccd1 vccd1 _15784_/A sky130_fd_sc_hd__xnor2_1
X_12993_ _12993_/A _12993_/B _12991_/X vssd1 vssd1 vccd1 vccd1 _12993_/X sky130_fd_sc_hd__or3b_1
XFILLER_57_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17520_ fanout942/X _17520_/D vssd1 vssd1 vccd1 vccd1 _17520_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14732_ _14756_/A1 _14730_/Y _14731_/X _14705_/Y _14706_/X vssd1 vssd1 vccd1 vccd1
+ _17604_/D sky130_fd_sc_hd__a32o_1
X_11944_ _11940_/X _11941_/Y _08868_/X _08873_/C vssd1 vssd1 vccd1 vccd1 _11944_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_55_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_62 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17451_ fanout951/X _17451_/D vssd1 vssd1 vccd1 vccd1 _17451_/Q sky130_fd_sc_hd__dfxtp_1
X_11875_ _12085_/B _11875_/B vssd1 vssd1 vccd1 vccd1 _11877_/C sky130_fd_sc_hd__nand2_1
X_14663_ _14664_/A _14669_/B vssd1 vssd1 vccd1 vccd1 _14663_/Y sky130_fd_sc_hd__nand2_1
XTAP_2974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16402_ _12235_/C _17075_/A2 _16401_/X vssd1 vssd1 vccd1 vccd1 _16404_/B sky130_fd_sc_hd__a21oi_1
X_10826_ _11115_/B _10963_/C _11117_/D _11115_/A vssd1 vssd1 vccd1 vccd1 _10827_/B
+ sky130_fd_sc_hd__a22oi_1
X_13614_ _13614_/A _13614_/B vssd1 vssd1 vccd1 vccd1 _13618_/A sky130_fd_sc_hd__xor2_2
X_17382_ input67/X _17424_/A2 _17381_/X _17388_/C1 vssd1 vssd1 vccd1 vccd1 _17519_/D
+ sky130_fd_sc_hd__o211a_1
X_14594_ _14594_/A _14594_/B vssd1 vssd1 vccd1 vccd1 _14597_/A sky130_fd_sc_hd__or2_1
XFILLER_60_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_90 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16333_ _16827_/A _16334_/C _16827_/B _16334_/A vssd1 vssd1 vccd1 vccd1 _16333_/X
+ sky130_fd_sc_hd__o22a_1
X_10757_ _10757_/A _10757_/B _10757_/C vssd1 vssd1 vccd1 vccd1 _11726_/A sky130_fd_sc_hd__or3_1
X_13545_ _13545_/A _13545_/B _13545_/C vssd1 vssd1 vccd1 vccd1 _13545_/X sky130_fd_sc_hd__and3_1
XFILLER_9_522 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16264_ _16358_/B _16264_/B vssd1 vssd1 vccd1 vccd1 _16266_/A sky130_fd_sc_hd__nor2_1
XFILLER_158_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13476_ _13476_/A _13476_/B vssd1 vssd1 vccd1 vccd1 _13479_/A sky130_fd_sc_hd__xor2_1
X_10688_ _10688_/A _10688_/B vssd1 vssd1 vccd1 vccd1 _10784_/A sky130_fd_sc_hd__nand2_2
XFILLER_145_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12427_ _12427_/A _12427_/B vssd1 vssd1 vccd1 vccd1 _12429_/C sky130_fd_sc_hd__xnor2_1
X_15215_ _15278_/A _16317_/B vssd1 vssd1 vccd1 vccd1 _15216_/B sky130_fd_sc_hd__nand2_1
XFILLER_173_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16195_ _16195_/A _16195_/B vssd1 vssd1 vccd1 vccd1 _16195_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_127_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15146_ _15553_/A _15553_/B _15493_/A vssd1 vssd1 vccd1 vccd1 _15155_/A sky130_fd_sc_hd__or3_1
X_12358_ _12526_/A _12358_/B _12358_/C vssd1 vssd1 vccd1 vccd1 _12526_/B sky130_fd_sc_hd__nand3_2
XFILLER_114_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11309_ _11399_/A _11399_/B vssd1 vssd1 vccd1 vccd1 _11311_/B sky130_fd_sc_hd__nand2b_1
XFILLER_99_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15077_ _15147_/D _15077_/B vssd1 vssd1 vccd1 vccd1 _15077_/Y sky130_fd_sc_hd__nor2_1
X_12289_ _12267_/Y _12268_/X _12476_/B _12290_/D vssd1 vssd1 vccd1 vccd1 _12289_/Y
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_141_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14028_ _14119_/B _14028_/B vssd1 vssd1 vccd1 vccd1 _14030_/C sky130_fd_sc_hd__nand2b_1
XFILLER_45_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_854 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_779 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15979_ _15980_/A _15980_/B _15980_/C vssd1 vssd1 vccd1 vccd1 _15979_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_49_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_578 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09003_ _09003_/A _09003_/B vssd1 vssd1 vccd1 vccd1 _09004_/B sky130_fd_sc_hd__xnor2_1
XFILLER_118_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout501 _10271_/A vssd1 vssd1 vccd1 vccd1 _11097_/C sky130_fd_sc_hd__buf_2
XFILLER_99_860 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09905_ _09909_/A vssd1 vssd1 vccd1 vccd1 _09910_/A sky130_fd_sc_hd__inv_2
XFILLER_104_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout512 _11370_/A vssd1 vssd1 vccd1 vccd1 _10638_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_160_798 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout523 _09894_/C vssd1 vssd1 vccd1 vccd1 _09321_/C sky130_fd_sc_hd__clkbuf_2
Xfanout534 _12471_/A vssd1 vssd1 vccd1 vccd1 _14842_/A1 sky130_fd_sc_hd__clkbuf_2
Xfanout545 _17515_/Q vssd1 vssd1 vccd1 vccd1 _09899_/A sky130_fd_sc_hd__buf_4
XFILLER_58_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout556 _09899_/B vssd1 vssd1 vccd1 vccd1 _11506_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout567 _17513_/Q vssd1 vssd1 vccd1 vccd1 _17112_/A1 sky130_fd_sc_hd__clkbuf_2
X_09836_ _10366_/A _09838_/C _09695_/A _09693_/Y vssd1 vssd1 vccd1 vccd1 _09842_/B
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout578 _17513_/Q vssd1 vssd1 vccd1 vccd1 fanout578/X sky130_fd_sc_hd__clkbuf_4
Xfanout589 _17512_/Q vssd1 vssd1 vccd1 vccd1 _10991_/A sky130_fd_sc_hd__clkbuf_2
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_470 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09767_ _09761_/A _09765_/X _09776_/A _09745_/Y vssd1 vssd1 vccd1 vccd1 _09776_/B
+ sky130_fd_sc_hd__o211ai_2
XTAP_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08718_ _15457_/A vssd1 vssd1 vccd1 vccd1 _11849_/A sky130_fd_sc_hd__clkinv_2
XTAP_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09698_ _10694_/A _10241_/B _12338_/C _09843_/C vssd1 vssd1 vccd1 vccd1 _09706_/A
+ sky130_fd_sc_hd__and4_1
XTAP_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_440 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11660_ _11678_/A _11681_/B vssd1 vssd1 vccd1 vccd1 _11662_/B sky130_fd_sc_hd__nor2_1
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10611_ _10711_/A _10711_/B vssd1 vssd1 vccd1 vccd1 _10611_/Y sky130_fd_sc_hd__nand2_1
XFILLER_41_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11591_ _11629_/A _11592_/B vssd1 vssd1 vccd1 vccd1 _11595_/B sky130_fd_sc_hd__and2_1
XFILLER_41_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13330_ _13330_/A _13330_/B vssd1 vssd1 vccd1 vccd1 _13332_/C sky130_fd_sc_hd__nand2_1
X_10542_ _11651_/A _12054_/B vssd1 vssd1 vccd1 vccd1 _10543_/C sky130_fd_sc_hd__and2_2
XFILLER_155_515 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13261_ _13261_/A _13261_/B _13261_/C vssd1 vssd1 vccd1 vccd1 _13263_/A sky130_fd_sc_hd__nand3_1
X_10473_ _10473_/A _10473_/B vssd1 vssd1 vccd1 vccd1 _10571_/A sky130_fd_sc_hd__xnor2_1
XFILLER_41_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12212_ _11809_/Y _11814_/Y _12212_/S vssd1 vssd1 vccd1 vccd1 _12212_/X sky130_fd_sc_hd__mux2_1
X_15000_ _14998_/Y _14999_/Y _15254_/S vssd1 vssd1 vccd1 vccd1 _15538_/B sky130_fd_sc_hd__mux2_1
XFILLER_142_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13192_ _13188_/X _13190_/Y _13061_/A _13063_/A vssd1 vssd1 vccd1 vccd1 _13202_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_123_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_592 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12143_ _12143_/A _12143_/B vssd1 vssd1 vccd1 vccd1 _12145_/B sky130_fd_sc_hd__xor2_1
XFILLER_2_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16951_ _16952_/A _16952_/B _16952_/C vssd1 vssd1 vccd1 vccd1 _16953_/A sky130_fd_sc_hd__a21oi_1
X_12074_ _12075_/B _12075_/A vssd1 vssd1 vccd1 vccd1 _12252_/A sky130_fd_sc_hd__and2b_1
XFILLER_96_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11025_ _11025_/A _11025_/B vssd1 vssd1 vccd1 vccd1 _11025_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_49_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15902_ _16011_/A _15252_/X _16012_/S vssd1 vssd1 vccd1 vccd1 _15902_/X sky130_fd_sc_hd__o21a_1
X_16882_ _16882_/A _16882_/B vssd1 vssd1 vccd1 vccd1 _16886_/A sky130_fd_sc_hd__or2_1
XFILLER_77_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15833_ _15834_/A _15834_/B vssd1 vssd1 vccd1 vccd1 _15966_/A sky130_fd_sc_hd__nand2_1
XFILLER_66_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15764_ _15764_/A _15764_/B _15764_/C vssd1 vssd1 vccd1 vccd1 _15765_/C sky130_fd_sc_hd__and3_1
XFILLER_80_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12976_ _12976_/A _12976_/B _12975_/X vssd1 vssd1 vccd1 vccd1 _12978_/A sky130_fd_sc_hd__or3b_1
XFILLER_18_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17503_ fanout946/X _17503_/D vssd1 vssd1 vccd1 vccd1 _17503_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14715_ _14742_/A _14715_/B vssd1 vssd1 vccd1 vccd1 _14717_/B sky130_fd_sc_hd__nand2_1
XTAP_3494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11927_ _17375_/A _11895_/C _08856_/A _08854_/B vssd1 vssd1 vccd1 vccd1 _11935_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_18_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15695_ _15786_/A _15693_/Y _15595_/A _15599_/A vssd1 vssd1 vccd1 vccd1 _15695_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17434_ fanout941/X _17434_/D vssd1 vssd1 vccd1 vccd1 _17434_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14646_ _14646_/A _14646_/B vssd1 vssd1 vccd1 vccd1 _14710_/C sky130_fd_sc_hd__nand2_1
XFILLER_162_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_819 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11858_ _12068_/B _12500_/B _11859_/D _12068_/A vssd1 vssd1 vccd1 vccd1 _11860_/A
+ sky130_fd_sc_hd__a22oi_1
X_10809_ _11095_/A _11095_/B _17469_/D _17468_/D vssd1 vssd1 vccd1 vccd1 _10812_/A
+ sky130_fd_sc_hd__and4_1
X_17365_ _17365_/A _17377_/B vssd1 vssd1 vccd1 vccd1 _17365_/Y sky130_fd_sc_hd__nand2_1
XANTENNA_19 _17063_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11789_ _16108_/C _14873_/B _11790_/A vssd1 vssd1 vccd1 vccd1 _11789_/X sky130_fd_sc_hd__or3_1
XFILLER_60_498 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14577_ _14577_/A _14577_/B vssd1 vssd1 vccd1 vccd1 _14579_/B sky130_fd_sc_hd__xnor2_1
XFILLER_159_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16316_ _16316_/A _16316_/B vssd1 vssd1 vccd1 vccd1 _16318_/A sky130_fd_sc_hd__nand2_1
X_13528_ _13637_/B _13527_/B _13527_/C vssd1 vssd1 vccd1 vccd1 _13529_/B sky130_fd_sc_hd__a21o_1
XFILLER_119_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17296_ _17353_/B _17353_/C vssd1 vssd1 vccd1 vccd1 _17296_/Y sky130_fd_sc_hd__nor2_1
XFILLER_118_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16247_ _16760_/B _16589_/B _16246_/C vssd1 vssd1 vccd1 vccd1 _16248_/B sky130_fd_sc_hd__a21oi_1
X_13459_ _13459_/A _13459_/B vssd1 vssd1 vccd1 vccd1 _13460_/B sky130_fd_sc_hd__or2_1
XFILLER_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_879 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput104 _17462_/Q vssd1 vssd1 vccd1 vccd1 o_wb_data[28] sky130_fd_sc_hd__clkbuf_1
X_16178_ _16179_/A _16179_/B vssd1 vssd1 vccd1 vccd1 _16279_/C sky130_fd_sc_hd__and2_1
Xoutput115 _17443_/Q vssd1 vssd1 vccd1 vccd1 o_wb_data[9] sky130_fd_sc_hd__clkbuf_1
XFILLER_114_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15129_ _10594_/B _10479_/B _10359_/B _14788_/B _10430_/A _10545_/C vssd1 vssd1 vccd1
+ vccd1 _15129_/X sky130_fd_sc_hd__mux4_1
XFILLER_99_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_307 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09621_ _09621_/A _09621_/B _09621_/C vssd1 vssd1 vccd1 vccd1 _09621_/X sky130_fd_sc_hd__and3_1
XFILLER_55_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09552_ _09552_/A _09696_/A vssd1 vssd1 vccd1 vccd1 _09559_/B sky130_fd_sc_hd__nor2_1
XFILLER_83_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09483_ _09483_/A _09483_/B vssd1 vssd1 vccd1 vccd1 _09484_/C sky130_fd_sc_hd__xnor2_1
XFILLER_64_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_988 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_802 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwire209 wire209/A vssd1 vssd1 vccd1 vccd1 wire209/X sky130_fd_sc_hd__clkbuf_2
XFILLER_127_8 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_34 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout320 _14832_/A vssd1 vssd1 vccd1 vccd1 _13434_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_59_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout331 _17134_/A vssd1 vssd1 vccd1 vccd1 _14708_/B sky130_fd_sc_hd__buf_2
Xfanout342 _14153_/A vssd1 vssd1 vccd1 vccd1 _13977_/A sky130_fd_sc_hd__buf_2
XFILLER_87_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout353 _14766_/A vssd1 vssd1 vccd1 vccd1 _14599_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_143_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout364 _16913_/C vssd1 vssd1 vccd1 vccd1 _14167_/A sky130_fd_sc_hd__buf_2
Xfanout375 fanout380/X vssd1 vssd1 vccd1 vccd1 _13450_/B sky130_fd_sc_hd__buf_2
XFILLER_19_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout386 _12788_/A vssd1 vssd1 vccd1 vccd1 _17409_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_86_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout397 _13578_/A vssd1 vssd1 vccd1 vccd1 _13908_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_09819_ _09819_/A _09819_/B _09819_/C vssd1 vssd1 vccd1 vccd1 _09822_/A sky130_fd_sc_hd__nor3_1
XFILLER_59_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12830_ _12672_/X _12674_/Y _12991_/A _12829_/Y vssd1 vssd1 vccd1 vccd1 _12991_/B
+ sky130_fd_sc_hd__a211oi_2
XFILLER_46_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12761_ _12761_/A _12761_/B _12761_/C vssd1 vssd1 vccd1 vccd1 _12762_/B sky130_fd_sc_hd__nor3_1
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14500_ _14501_/B _14500_/B vssd1 vssd1 vccd1 vccd1 _14502_/A sky130_fd_sc_hd__nand2b_1
XTAP_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11712_ _11713_/A _11713_/B vssd1 vssd1 vccd1 vccd1 _16294_/A sky130_fd_sc_hd__and2_1
XFILLER_14_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12692_ _12533_/X _12536_/B _12532_/Y vssd1 vssd1 vccd1 vccd1 _12694_/B sky130_fd_sc_hd__o21a_1
XTAP_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15480_ _15913_/A _15832_/A _15481_/B vssd1 vssd1 vccd1 vccd1 _15590_/A sky130_fd_sc_hd__or3_1
XTAP_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11643_ _11607_/B _11644_/C vssd1 vssd1 vccd1 vccd1 _11648_/B sky130_fd_sc_hd__nand2b_1
XFILLER_14_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14431_ _14497_/B _14431_/B vssd1 vssd1 vccd1 vccd1 _14463_/A sky130_fd_sc_hd__nor2_1
XFILLER_30_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17150_ _17125_/A _17128_/A _17131_/B _17149_/X _17063_/A vssd1 vssd1 vccd1 vccd1
+ _17150_/X sky130_fd_sc_hd__a41o_1
XFILLER_52_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11574_ _11574_/A _11607_/A _11574_/C vssd1 vssd1 vccd1 vccd1 _11579_/A sky130_fd_sc_hd__or3_1
XFILLER_128_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14362_ _17100_/C _14865_/B vssd1 vssd1 vccd1 vccd1 _14364_/B sky130_fd_sc_hd__nand2_1
XFILLER_10_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput17 i_wb_addr[22] vssd1 vssd1 vccd1 vccd1 input17/X sky130_fd_sc_hd__clkbuf_1
XFILLER_168_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput28 i_wb_addr[3] vssd1 vssd1 vccd1 vccd1 input28/X sky130_fd_sc_hd__clkbuf_2
X_16101_ _15991_/X _15994_/X _16203_/A vssd1 vssd1 vccd1 vccd1 _16101_/Y sky130_fd_sc_hd__o21bai_2
XFILLER_155_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10525_ _10638_/A _10638_/B _10743_/D _10525_/D vssd1 vssd1 vccd1 vccd1 _10528_/A
+ sky130_fd_sc_hd__and4_1
X_13313_ _13314_/B _13314_/C _13314_/A vssd1 vssd1 vccd1 vccd1 _13442_/A sky130_fd_sc_hd__o21ai_1
Xinput39 i_wb_data[12] vssd1 vssd1 vccd1 vccd1 input39/X sky130_fd_sc_hd__clkbuf_1
X_14293_ _14294_/A _14294_/B vssd1 vssd1 vccd1 vccd1 _14372_/B sky130_fd_sc_hd__nor2_1
X_17081_ _17081_/A _17081_/B _17038_/B vssd1 vssd1 vccd1 vccd1 _17083_/B sky130_fd_sc_hd__or3b_1
XFILLER_6_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16032_ _16032_/A _16032_/B vssd1 vssd1 vccd1 vccd1 _16034_/A sky130_fd_sc_hd__or2_1
X_13244_ _13244_/A _13244_/B _13244_/C vssd1 vssd1 vccd1 vccd1 _13246_/A sky130_fd_sc_hd__nand3_1
XFILLER_171_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10456_ _10564_/A _10456_/B vssd1 vssd1 vccd1 vccd1 _10459_/B sky130_fd_sc_hd__xor2_1
XFILLER_170_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13175_ _13176_/A _13176_/B vssd1 vssd1 vccd1 vccd1 _13314_/C sky130_fd_sc_hd__and2b_1
XFILLER_124_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10387_ _10387_/A _10387_/B vssd1 vssd1 vccd1 vccd1 _10388_/B sky130_fd_sc_hd__nor2_1
XFILLER_124_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12126_ _17423_/A _12127_/C _12127_/D _17425_/A vssd1 vssd1 vccd1 vccd1 _12128_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_151_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_649 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12057_ _12047_/X _12056_/X _13833_/S vssd1 vssd1 vccd1 vccd1 _12057_/X sky130_fd_sc_hd__mux2_1
X_16934_ _16990_/A _09852_/A _17083_/A _16933_/Y vssd1 vssd1 vccd1 vccd1 _16935_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_42_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11008_ _10805_/D _11006_/X _11007_/X vssd1 vssd1 vccd1 vccd1 _11009_/B sky130_fd_sc_hd__a21bo_1
XFILLER_65_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16865_ _16865_/A _16865_/B vssd1 vssd1 vccd1 vccd1 _16865_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_92_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15816_ _16315_/B _16938_/B vssd1 vssd1 vccd1 vccd1 _15825_/A sky130_fd_sc_hd__nor2_1
XFILLER_53_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16796_ _16796_/A _16796_/B vssd1 vssd1 vccd1 vccd1 _16797_/B sky130_fd_sc_hd__nand2_1
XFILLER_93_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_782 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15747_ _15493_/A _16814_/A _16165_/B _16056_/A vssd1 vssd1 vccd1 vccd1 _15747_/X
+ sky130_fd_sc_hd__a2bb2o_1
XTAP_3291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12959_ _12959_/A _12959_/B vssd1 vssd1 vccd1 vccd1 _12960_/B sky130_fd_sc_hd__nand2_1
XFILLER_34_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15678_ _15674_/X _15676_/A _15572_/Y _15583_/Y vssd1 vssd1 vccd1 vccd1 _15679_/C
+ sky130_fd_sc_hd__o211ai_1
XFILLER_61_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17417_ _17417_/A _17421_/B vssd1 vssd1 vccd1 vccd1 _17417_/X sky130_fd_sc_hd__or2_1
XFILLER_60_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14629_ _14629_/A _14629_/B _14629_/C vssd1 vssd1 vccd1 vccd1 _14631_/A sky130_fd_sc_hd__and3_1
XFILLER_159_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17348_ _11902_/B _17356_/A2 _17347_/X _17420_/C1 vssd1 vssd1 vccd1 vccd1 _17503_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_119_526 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17279_ _17602_/Q _17282_/A2 _17282_/B1 vssd1 vssd1 vccd1 vccd1 _17279_/X sky130_fd_sc_hd__a21o_1
XFILLER_146_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1042 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08983_ _08983_/A _08983_/B vssd1 vssd1 vccd1 vccd1 _08984_/B sky130_fd_sc_hd__or2_1
XFILLER_69_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09604_ _09892_/A _09892_/B _10545_/D _10299_/D vssd1 vssd1 vccd1 vccd1 _09607_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_113_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09535_ _12005_/B _09397_/X _09531_/X _09540_/A vssd1 vssd1 vccd1 vccd1 _09536_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_37_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09466_ _09473_/A _09465_/Y _09894_/C _10311_/D vssd1 vssd1 vccd1 vccd1 _09591_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_169_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09397_ _12005_/A _09395_/X _09343_/X _09393_/B vssd1 vssd1 vccd1 vccd1 _09397_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_138_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10310_ _10753_/A _10308_/B _09926_/C vssd1 vssd1 vccd1 vccd1 _10310_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_98_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11290_ _11295_/A _11295_/B vssd1 vssd1 vccd1 vccd1 _11290_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_98_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10241_ _10591_/A _10241_/B _10359_/B _10479_/B vssd1 vssd1 vccd1 vccd1 _10243_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_133_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10172_ _10419_/B _10299_/D _10171_/D _14789_/A vssd1 vssd1 vccd1 vccd1 _10172_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_152_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14980_ _15096_/S _14978_/Y _14979_/Y _15097_/A vssd1 vssd1 vccd1 vccd1 _15252_/B
+ sky130_fd_sc_hd__a211o_1
Xfanout150 _15100_/A vssd1 vssd1 vccd1 vccd1 _15131_/A sky130_fd_sc_hd__clkbuf_4
Xfanout161 _17389_/B vssd1 vssd1 vccd1 vccd1 _17425_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_47_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_811 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout172 _16743_/B vssd1 vssd1 vccd1 vccd1 _16809_/C sky130_fd_sc_hd__clkbuf_4
Xfanout183 _15472_/Y vssd1 vssd1 vccd1 vccd1 _16681_/A sky130_fd_sc_hd__clkbuf_2
X_13931_ _13932_/A _13932_/B vssd1 vssd1 vccd1 vccd1 _14032_/A sky130_fd_sc_hd__nor2_1
Xfanout194 _15145_/X vssd1 vssd1 vccd1 vccd1 _16055_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_87_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16650_ _16649_/A _16649_/B _16649_/C vssd1 vssd1 vccd1 vccd1 _16650_/Y sky130_fd_sc_hd__a21oi_1
X_13862_ _13862_/A _13964_/A _13862_/C vssd1 vssd1 vccd1 vccd1 _13862_/X sky130_fd_sc_hd__and3_1
XFILLER_47_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15601_ _15601_/A _15601_/B vssd1 vssd1 vccd1 vccd1 _15604_/A sky130_fd_sc_hd__xor2_1
XFILLER_170_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12813_ _12663_/B _12665_/B _12663_/A vssd1 vssd1 vccd1 vccd1 _12976_/B sky130_fd_sc_hd__o21ba_1
X_16581_ _12869_/C _17075_/A2 _16580_/X vssd1 vssd1 vccd1 vccd1 _16581_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_27_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13793_ _13793_/A _13793_/B _13793_/C vssd1 vssd1 vccd1 vccd1 _13795_/A sky130_fd_sc_hd__or3_1
XFILLER_90_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15532_ _15532_/A _15532_/B vssd1 vssd1 vccd1 vccd1 _15533_/B sky130_fd_sc_hd__nand2_1
X_12744_ _12744_/A _12902_/B vssd1 vssd1 vccd1 vccd1 _12747_/A sky130_fd_sc_hd__and2_1
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15463_ _15463_/A _15463_/B vssd1 vssd1 vccd1 vccd1 _15463_/Y sky130_fd_sc_hd__nor2_1
X_12675_ _12675_/A _12675_/B vssd1 vssd1 vccd1 vccd1 _12676_/C sky130_fd_sc_hd__xor2_1
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17202_ _17544_/Q _17274_/B vssd1 vssd1 vccd1 vccd1 _17202_/X sky130_fd_sc_hd__and2_1
X_14414_ _14414_/A _14414_/B vssd1 vssd1 vccd1 vccd1 _14533_/A sky130_fd_sc_hd__nor2_1
X_11626_ _11672_/A _11672_/B vssd1 vssd1 vccd1 vccd1 _15524_/B sky130_fd_sc_hd__and2_1
X_15394_ _15071_/A _11789_/X _16315_/D vssd1 vssd1 vccd1 vccd1 _15472_/B sky130_fd_sc_hd__a21oi_2
XFILLER_168_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17133_ _17133_/A vssd1 vssd1 vccd1 vccd1 _17133_/Y sky130_fd_sc_hd__inv_2
X_14345_ _14413_/A _14345_/B vssd1 vssd1 vccd1 vccd1 _14348_/A sky130_fd_sc_hd__nor2_1
X_11557_ _11558_/A _11558_/B _11558_/C vssd1 vssd1 vccd1 vccd1 _11557_/X sky130_fd_sc_hd__and3_1
XFILLER_11_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10508_ _10509_/A _10507_/Y _10719_/C _10508_/D vssd1 vssd1 vccd1 vccd1 _10617_/A
+ sky130_fd_sc_hd__and4bb_1
X_17064_ _14765_/A _16965_/B _17065_/A vssd1 vssd1 vccd1 vccd1 _17064_/X sky130_fd_sc_hd__a21bo_1
X_11488_ _11487_/A _11527_/A _11444_/Y _11466_/X vssd1 vssd1 vccd1 vccd1 _11496_/B
+ sky130_fd_sc_hd__o211ai_2
X_14276_ _14276_/A _14276_/B _14274_/X vssd1 vssd1 vccd1 vccd1 _14277_/B sky130_fd_sc_hd__or3b_1
XFILLER_143_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16015_ _16015_/A _16114_/B _16015_/C vssd1 vssd1 vccd1 vccd1 _16015_/X sky130_fd_sc_hd__or3_1
X_13227_ _13227_/A _14153_/B _13664_/D _13551_/D vssd1 vssd1 vccd1 vccd1 _13228_/B
+ sky130_fd_sc_hd__and4_1
X_10439_ _10425_/Y _10437_/X _10453_/A _10410_/Y vssd1 vssd1 vccd1 vccd1 _10453_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_98_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13158_ _13643_/A _13908_/B vssd1 vssd1 vccd1 vccd1 _13159_/B sky130_fd_sc_hd__nand2_1
XFILLER_151_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12109_ _12907_/A _12445_/D vssd1 vssd1 vccd1 vccd1 _12110_/B sky130_fd_sc_hd__nand2_1
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13089_ _13903_/A _13966_/C _13088_/C vssd1 vssd1 vccd1 vccd1 _13090_/B sky130_fd_sc_hd__a21o_1
XFILLER_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16917_ _16917_/A _16917_/B vssd1 vssd1 vccd1 vccd1 _16917_/Y sky130_fd_sc_hd__nand2_1
XFILLER_38_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16848_ _16848_/A vssd1 vssd1 vccd1 vccd1 _16850_/B sky130_fd_sc_hd__inv_2
XFILLER_53_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16779_ _16699_/A _16698_/B _16698_/A vssd1 vssd1 vccd1 vccd1 _16781_/B sky130_fd_sc_hd__a21boi_1
X_09320_ _11895_/B _09319_/C _09319_/D _17379_/A vssd1 vssd1 vccd1 vccd1 _09320_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_81_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09251_ _09248_/Y _09249_/X _09115_/A _09114_/Y vssd1 vssd1 vccd1 vccd1 _09251_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_61_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09182_ _09214_/A vssd1 vssd1 vccd1 vccd1 _09182_/Y sky130_fd_sc_hd__inv_2
XFILLER_105_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_356 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_36 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08966_ _08993_/C _08965_/Y _08963_/X vssd1 vssd1 vccd1 vccd1 _08973_/A sky130_fd_sc_hd__o21a_1
XFILLER_124_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08897_ _17391_/A _17389_/A _09042_/B _10297_/D vssd1 vssd1 vccd1 vccd1 _08900_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_112_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_77 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09518_ _09519_/B _09519_/A vssd1 vssd1 vccd1 vccd1 _09522_/B sky130_fd_sc_hd__and2b_1
XFILLER_169_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10790_ _10901_/B _10796_/B vssd1 vssd1 vccd1 vccd1 _10860_/A sky130_fd_sc_hd__nor2_1
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09449_ _09449_/A _09449_/B vssd1 vssd1 vccd1 vccd1 _09578_/A sky130_fd_sc_hd__xnor2_1
XPHY_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12460_ _12457_/X _12458_/Y _12267_/Y _12290_/X vssd1 vssd1 vccd1 vccd1 _12481_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_130_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11411_ _11411_/A _11411_/B vssd1 vssd1 vccd1 vccd1 _11419_/B sky130_fd_sc_hd__xor2_2
XFILLER_32_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12391_ _12389_/X _12390_/X _12865_/S vssd1 vssd1 vccd1 vccd1 _12391_/X sky130_fd_sc_hd__mux2_1
X_11342_ _11329_/Y _11367_/A _11343_/A _11312_/Y vssd1 vssd1 vccd1 vccd1 _11349_/A
+ sky130_fd_sc_hd__o211ai_1
XFILLER_4_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14130_ _14130_/A _14134_/B _13958_/C vssd1 vssd1 vccd1 vccd1 _14131_/A sky130_fd_sc_hd__nor3b_1
XFILLER_138_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_646 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11273_ _11274_/B _11274_/C _11274_/A vssd1 vssd1 vccd1 vccd1 _11285_/A sky130_fd_sc_hd__a21o_1
XFILLER_152_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14061_ _13967_/A _13969_/B _13967_/B vssd1 vssd1 vccd1 vccd1 _14068_/A sky130_fd_sc_hd__o21ba_1
XFILLER_4_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13012_ _13516_/S _11833_/X _11854_/C _12858_/Y vssd1 vssd1 vccd1 vccd1 _13012_/X
+ sky130_fd_sc_hd__o22a_2
X_10224_ _10226_/A _10226_/B _10221_/X vssd1 vssd1 vccd1 vccd1 _10348_/C sky130_fd_sc_hd__a21oi_1
XFILLER_134_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10155_ _10155_/A _10155_/B vssd1 vssd1 vccd1 vccd1 _10155_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_928 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10086_ _10086_/A _10086_/B _10086_/C vssd1 vssd1 vccd1 vccd1 _10216_/A sky130_fd_sc_hd__or3_1
X_14963_ _15175_/A _15808_/A vssd1 vssd1 vccd1 vccd1 _14963_/X sky130_fd_sc_hd__or2_2
XFILLER_59_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16702_ _16777_/B _16702_/B vssd1 vssd1 vccd1 vccd1 _16705_/A sky130_fd_sc_hd__nand2_1
X_13914_ _13915_/A _13915_/B _13915_/C vssd1 vssd1 vccd1 vccd1 _14021_/A sky130_fd_sc_hd__o21a_1
XFILLER_47_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14894_ _16938_/A _15709_/A _15617_/A vssd1 vssd1 vccd1 vccd1 _15208_/D sky130_fd_sc_hd__or3_1
XFILLER_35_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16633_ _16634_/A _16634_/B vssd1 vssd1 vccd1 vccd1 _16711_/B sky130_fd_sc_hd__nor2_1
XFILLER_74_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13845_ _13845_/A _13954_/A vssd1 vssd1 vccd1 vccd1 _13848_/A sky130_fd_sc_hd__nor2_1
XFILLER_74_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_858 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16564_ _16564_/A _16564_/B vssd1 vssd1 vccd1 vccd1 _16564_/Y sky130_fd_sc_hd__nor2_1
XFILLER_90_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13776_ _13776_/A _13776_/B vssd1 vssd1 vccd1 vccd1 _13778_/C sky130_fd_sc_hd__xnor2_1
XFILLER_90_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10988_ _10990_/A _10990_/B _10990_/C vssd1 vssd1 vccd1 vccd1 _10988_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_128_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15515_ _15609_/A _15515_/B vssd1 vssd1 vccd1 vccd1 _15518_/A sky130_fd_sc_hd__nor2_1
XFILLER_149_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12727_ _12727_/A _12727_/B vssd1 vssd1 vccd1 vccd1 _12728_/B sky130_fd_sc_hd__nor2_1
X_16495_ _16495_/A vssd1 vssd1 vccd1 vccd1 _17562_/D sky130_fd_sc_hd__inv_2
XFILLER_148_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15446_ _11672_/Y _11694_/X _11693_/Y _11691_/Y vssd1 vssd1 vccd1 vccd1 _15446_/Y
+ sky130_fd_sc_hd__a211oi_1
X_12658_ _12658_/A _12658_/B vssd1 vssd1 vccd1 vccd1 _12660_/A sky130_fd_sc_hd__nor2_1
XFILLER_90_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11609_ _11610_/A _11610_/B vssd1 vssd1 vccd1 vccd1 _11617_/A sky130_fd_sc_hd__or2_1
X_15377_ _15374_/X _15375_/X _15376_/Y vssd1 vssd1 vccd1 vccd1 _15377_/Y sky130_fd_sc_hd__o21ai_1
X_12589_ _12452_/A _12452_/B _12450_/X vssd1 vssd1 vccd1 vccd1 _12610_/A sky130_fd_sc_hd__a21oi_2
XFILLER_128_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17116_ _14867_/A _17170_/B1 _17103_/X _17115_/X vssd1 vssd1 vccd1 vccd1 _17572_/D
+ sky130_fd_sc_hd__a22oi_1
XFILLER_7_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14328_ _14393_/B _14328_/B vssd1 vssd1 vccd1 vccd1 _14330_/C sky130_fd_sc_hd__nand2_1
XFILLER_128_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17047_ _17088_/A _17047_/B vssd1 vssd1 vccd1 vccd1 _17049_/B sky130_fd_sc_hd__nor2_1
X_14259_ _14164_/X _14186_/A _14257_/Y _14258_/X vssd1 vssd1 vccd1 vccd1 _14340_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_99_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout908 _11095_/D vssd1 vssd1 vccd1 vccd1 _11605_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout919 _17245_/A2 vssd1 vssd1 vccd1 vccd1 _17293_/A2 sky130_fd_sc_hd__buf_2
XFILLER_140_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08820_ _08821_/A _08821_/C vssd1 vssd1 vccd1 vccd1 _08822_/B sky130_fd_sc_hd__nor2_1
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_896 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08751_ _17403_/A _17399_/A _12328_/B _09229_/B vssd1 vssd1 vccd1 vccd1 _08755_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_39_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_622 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1022 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09303_ _09304_/B _09304_/A vssd1 vssd1 vccd1 vccd1 _09303_/X sky130_fd_sc_hd__and2b_1
XFILLER_110_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_1019 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09234_ _09234_/A _09234_/B vssd1 vssd1 vccd1 vccd1 _09236_/A sky130_fd_sc_hd__nor2_1
XFILLER_148_930 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09165_ _09165_/A _09165_/B _09168_/B vssd1 vssd1 vccd1 vccd1 _09178_/A sky130_fd_sc_hd__or3_1
XFILLER_119_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_13 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09096_ _11839_/S _14765_/B vssd1 vssd1 vccd1 vccd1 _14981_/A sky130_fd_sc_hd__and2_1
XFILLER_119_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_635 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_167 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_906 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09998_ _10255_/A _10142_/B vssd1 vssd1 vccd1 vccd1 _10123_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08949_ _08950_/A _08948_/Y _17375_/A _12258_/B vssd1 vssd1 vccd1 vccd1 _09065_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_69_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11960_ _11960_/A _12169_/A vssd1 vssd1 vccd1 vccd1 _11961_/C sky130_fd_sc_hd__and2_1
XFILLER_17_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10911_ _11097_/C _10963_/C vssd1 vssd1 vccd1 vccd1 _10915_/A sky130_fd_sc_hd__nand2_1
XFILLER_56_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11891_ _11891_/A _11891_/B _11891_/C vssd1 vssd1 vccd1 vccd1 _11891_/Y sky130_fd_sc_hd__nor3_4
XFILLER_44_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13630_ _14734_/A _13624_/X _13629_/X vssd1 vssd1 vccd1 vccd1 _13630_/Y sky130_fd_sc_hd__a21oi_1
X_10842_ _10842_/A _10842_/B vssd1 vssd1 vccd1 vccd1 _10844_/B sky130_fd_sc_hd__xnor2_1
XFILLER_44_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13561_ _13557_/Y _13559_/A _13443_/B _13444_/Y vssd1 vssd1 vccd1 vccd1 _13562_/B
+ sky130_fd_sc_hd__o211a_1
X_10773_ _10667_/Y _10692_/X _10766_/C _11725_/A vssd1 vssd1 vccd1 vccd1 _10774_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_12_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15300_ _15233_/X _15299_/Y _08743_/A vssd1 vssd1 vccd1 vccd1 _15300_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_157_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12512_ _12344_/B _12346_/B _12344_/A vssd1 vssd1 vccd1 vccd1 _12514_/B sky130_fd_sc_hd__o21ba_1
XFILLER_157_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16280_ _16280_/A _16280_/B vssd1 vssd1 vccd1 vccd1 _16282_/A sky130_fd_sc_hd__nor2_1
XFILLER_9_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13492_ _13492_/A _13492_/B vssd1 vssd1 vccd1 vccd1 _13494_/C sky130_fd_sc_hd__nor2_1
XFILLER_157_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15231_ _15231_/A _15231_/B vssd1 vssd1 vccd1 vccd1 _15233_/A sky130_fd_sc_hd__nand2_1
X_12443_ _12443_/A _12616_/B vssd1 vssd1 vccd1 vccd1 _12452_/A sky130_fd_sc_hd__nor2_1
XFILLER_60_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15162_ _15162_/A _15162_/B vssd1 vssd1 vccd1 vccd1 _15166_/A sky130_fd_sc_hd__nand2_1
X_12374_ _12374_/A _12374_/B vssd1 vssd1 vccd1 vccd1 _12377_/B sky130_fd_sc_hd__nand2_1
XFILLER_165_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14113_ _14113_/A _14113_/B _14113_/C vssd1 vssd1 vccd1 vccd1 _14114_/B sky130_fd_sc_hd__nand3_1
X_11325_ _11325_/A _11376_/A vssd1 vssd1 vccd1 vccd1 _11369_/A sky130_fd_sc_hd__nand2_1
XFILLER_5_976 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15093_ _15093_/A _15093_/B vssd1 vssd1 vccd1 vccd1 _15170_/C sky130_fd_sc_hd__nand2_1
XFILLER_119_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11256_ _11255_/A _11255_/C _11255_/B vssd1 vssd1 vccd1 vccd1 _11256_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_125_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14044_ _14044_/A _14044_/B vssd1 vssd1 vccd1 vccd1 _14045_/B sky130_fd_sc_hd__nor2_1
XFILLER_69_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10207_ _10207_/A _10207_/B vssd1 vssd1 vccd1 vccd1 _10210_/A sky130_fd_sc_hd__nor2_1
X_11187_ _11202_/B _11186_/B _11218_/A _11186_/D vssd1 vssd1 vccd1 vccd1 _11187_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_121_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10138_ _10138_/A _10138_/B _10138_/C vssd1 vssd1 vccd1 vccd1 _10138_/Y sky130_fd_sc_hd__nand3_1
XFILLER_67_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15995_ _15994_/A _15993_/X _15523_/A vssd1 vssd1 vccd1 vccd1 _15995_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_95_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14946_ _14765_/B _15033_/A3 _17139_/A _11932_/B _09925_/A _15095_/B vssd1 vssd1
+ vccd1 vccd1 _14947_/B sky130_fd_sc_hd__mux4_1
X_10069_ _10069_/A _10069_/B _10200_/A vssd1 vssd1 vccd1 vccd1 _10070_/B sky130_fd_sc_hd__or3_1
XFILLER_78_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14877_ _17614_/Q _15147_/C _17613_/Q vssd1 vssd1 vccd1 vccd1 _14877_/Y sky130_fd_sc_hd__o21bai_4
XFILLER_35_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16616_ _16616_/A _16616_/B _16616_/C vssd1 vssd1 vccd1 vccd1 _16617_/B sky130_fd_sc_hd__nor3_1
XFILLER_35_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13828_ _13727_/A _13828_/B vssd1 vssd1 vccd1 vccd1 _13830_/B sky130_fd_sc_hd__and2b_1
XFILLER_50_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17596_ fanout936/X _17596_/D vssd1 vssd1 vccd1 vccd1 _17596_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16547_ _16547_/A _16547_/B vssd1 vssd1 vccd1 vccd1 _16548_/B sky130_fd_sc_hd__or2_1
X_13759_ _13656_/B _13659_/B _13654_/X vssd1 vssd1 vccd1 vccd1 _13761_/B sky130_fd_sc_hd__a21oi_1
XFILLER_93_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16478_ _16478_/A _16478_/B vssd1 vssd1 vccd1 vccd1 _16478_/X sky130_fd_sc_hd__or2_2
X_15429_ _15429_/A _15429_/B vssd1 vssd1 vccd1 vccd1 _15431_/A sky130_fd_sc_hd__xnor2_1
XFILLER_102_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09921_ _09922_/A _09922_/B vssd1 vssd1 vccd1 vccd1 _09923_/A sky130_fd_sc_hd__nand2_1
Xfanout705 _12088_/D vssd1 vssd1 vccd1 vccd1 _09319_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_113_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout716 _17498_/Q vssd1 vssd1 vccd1 vccd1 _10308_/B sky130_fd_sc_hd__buf_4
Xfanout727 _16399_/A vssd1 vssd1 vccd1 vccd1 _13866_/C sky130_fd_sc_hd__clkbuf_4
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09852_ _09852_/A _09852_/B vssd1 vssd1 vccd1 vccd1 _09854_/B sky130_fd_sc_hd__xnor2_4
Xfanout738 _10171_/D vssd1 vssd1 vccd1 vccd1 _11867_/D sky130_fd_sc_hd__clkbuf_4
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout749 _17494_/Q vssd1 vssd1 vccd1 vccd1 _14859_/B sky130_fd_sc_hd__buf_4
XFILLER_59_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08803_ _17401_/A _11961_/B _08772_/C _08772_/D vssd1 vssd1 vccd1 vccd1 _08804_/B
+ sky130_fd_sc_hd__a22oi_1
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09783_ _09783_/A _09930_/A vssd1 vssd1 vccd1 vccd1 _09784_/C sky130_fd_sc_hd__nor2_1
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08734_ _17608_/Q _17607_/Q vssd1 vssd1 vccd1 vccd1 _14836_/B sky130_fd_sc_hd__and2b_1
XFILLER_27_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_535 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09217_ _17409_/A _09555_/C vssd1 vssd1 vccd1 vccd1 _09219_/C sky130_fd_sc_hd__nand2_1
XFILLER_167_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09148_ _09148_/A _09148_/B vssd1 vssd1 vccd1 vccd1 _09150_/B sky130_fd_sc_hd__xnor2_1
XFILLER_147_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09079_ _11895_/B _09321_/D _09319_/C _17379_/A vssd1 vssd1 vccd1 vccd1 _09079_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_30_66 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11110_ _11110_/A _11110_/B _11110_/C vssd1 vssd1 vccd1 vccd1 _11144_/A sky130_fd_sc_hd__nand3_1
X_12090_ _17387_/A _12256_/C vssd1 vssd1 vccd1 vccd1 _12091_/B sky130_fd_sc_hd__nand2_1
XFILLER_1_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11041_ _11041_/A _11041_/B _11041_/C vssd1 vssd1 vccd1 vccd1 _11041_/Y sky130_fd_sc_hd__nand3_2
XFILLER_89_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14800_ _15244_/B _15244_/C _15244_/A vssd1 vssd1 vccd1 vccd1 _14801_/C sky130_fd_sc_hd__o21ba_1
XTAP_3610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15780_ _15781_/A _15781_/B vssd1 vssd1 vccd1 vccd1 _15883_/A sky130_fd_sc_hd__and2b_1
X_12992_ _12993_/A _12993_/B _12991_/X vssd1 vssd1 vccd1 vccd1 _12997_/A sky130_fd_sc_hd__nor3b_1
XFILLER_57_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14731_ _14731_/A _14731_/B vssd1 vssd1 vccd1 vccd1 _14731_/X sky130_fd_sc_hd__or2_1
X_11943_ _12156_/A vssd1 vssd1 vccd1 vccd1 _11943_/Y sky130_fd_sc_hd__inv_2
XTAP_2920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17450_ fanout951/X _17450_/D vssd1 vssd1 vccd1 vccd1 _17450_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14662_ _14662_/A _14662_/B vssd1 vssd1 vccd1 vccd1 _14669_/B sky130_fd_sc_hd__xnor2_2
XTAP_2964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11874_ _11874_/A _11874_/B vssd1 vssd1 vccd1 vccd1 _11875_/B sky130_fd_sc_hd__or2_1
XFILLER_45_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16401_ _16397_/B _16799_/A2 _16580_/B1 _16399_/A _16401_/C1 vssd1 vssd1 vccd1 vccd1
+ _16401_/X sky130_fd_sc_hd__a221o_1
X_13613_ _13578_/A _13464_/B _13465_/A _13463_/A vssd1 vssd1 vccd1 vccd1 _13614_/B
+ sky130_fd_sc_hd__a31o_1
X_10825_ _11115_/A _11115_/B _10963_/C _11117_/D vssd1 vssd1 vccd1 vccd1 _10827_/A
+ sky130_fd_sc_hd__and4_1
XTAP_2997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17381_ _17381_/A _17389_/B vssd1 vssd1 vccd1 vccd1 _17381_/X sky130_fd_sc_hd__or2_1
X_14593_ _14738_/A _14708_/B _14641_/D _14593_/D vssd1 vssd1 vccd1 vccd1 _14594_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_25_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16332_ _16245_/A _16245_/B _16248_/A vssd1 vssd1 vccd1 vccd1 _16342_/A sky130_fd_sc_hd__a21oi_1
X_13544_ _13545_/A _13545_/B _13545_/C vssd1 vssd1 vccd1 vccd1 _13662_/A sky130_fd_sc_hd__a21oi_2
X_10756_ _10756_/A _11165_/A vssd1 vssd1 vccd1 vccd1 _10757_/C sky130_fd_sc_hd__nor2_1
XFILLER_146_708 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16263_ _16262_/A _16681_/C _16262_/C vssd1 vssd1 vccd1 vccd1 _16264_/B sky130_fd_sc_hd__o21a_1
XFILLER_173_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13475_ _13476_/B _13476_/A vssd1 vssd1 vccd1 vccd1 _13590_/B sky130_fd_sc_hd__and2b_1
X_10687_ _10685_/B _10685_/C _10685_/A vssd1 vssd1 vccd1 vccd1 _10688_/B sky130_fd_sc_hd__a21o_1
X_15214_ _15214_/A _15494_/A vssd1 vssd1 vccd1 vccd1 _15216_/A sky130_fd_sc_hd__xnor2_1
X_12426_ _13302_/A _13704_/B vssd1 vssd1 vccd1 vccd1 _12427_/B sky130_fd_sc_hd__nand2_1
X_16194_ _16195_/A _16195_/B vssd1 vssd1 vccd1 vccd1 _16290_/A sky130_fd_sc_hd__nor2_1
XFILLER_126_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15145_ _14886_/D _15144_/X _15175_/A vssd1 vssd1 vccd1 vccd1 _15145_/X sky130_fd_sc_hd__a21o_1
X_12357_ _12357_/A _12357_/B vssd1 vssd1 vccd1 vccd1 _12358_/C sky130_fd_sc_hd__xnor2_1
XFILLER_153_251 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11308_ _11308_/A _11308_/B vssd1 vssd1 vccd1 vccd1 _11399_/B sky130_fd_sc_hd__xnor2_1
XFILLER_5_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15076_ _14967_/C _14967_/D _15075_/X _14877_/Y vssd1 vssd1 vccd1 vccd1 _15077_/B
+ sky130_fd_sc_hd__o22a_1
X_12288_ _12476_/A _12286_/Y _12112_/X _12116_/A vssd1 vssd1 vccd1 vccd1 _12290_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_141_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14027_ _14027_/A _14027_/B _14025_/Y vssd1 vssd1 vccd1 vccd1 _14028_/B sky130_fd_sc_hd__or3b_1
X_11239_ _15472_/A _17466_/D vssd1 vssd1 vccd1 vccd1 _11492_/A sky130_fd_sc_hd__nand2_1
XFILLER_95_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_888 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15978_ _15980_/A _15980_/B _15980_/C vssd1 vssd1 vccd1 vccd1 _15981_/A sky130_fd_sc_hd__o21a_1
XFILLER_48_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14929_ _14929_/A _14933_/B vssd1 vssd1 vccd1 vccd1 _14929_/X sky130_fd_sc_hd__or2_4
XFILLER_64_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17579_ fanout939/X _17579_/D vssd1 vssd1 vccd1 vccd1 _17579_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_524 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09002_ _09003_/A _09003_/B vssd1 vssd1 vccd1 vccd1 _09002_/X sky130_fd_sc_hd__and2b_1
XFILLER_129_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout502 _10271_/A vssd1 vssd1 vccd1 vccd1 _10719_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_132_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09904_ _09906_/B _10035_/A _09906_/A vssd1 vssd1 vccd1 vccd1 _09909_/A sky130_fd_sc_hd__a21o_1
XFILLER_99_872 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout513 _17518_/Q vssd1 vssd1 vccd1 vccd1 _11370_/A sky130_fd_sc_hd__clkbuf_4
Xfanout524 _12442_/A vssd1 vssd1 vccd1 vccd1 _09894_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_113_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout535 _09755_/A vssd1 vssd1 vccd1 vccd1 _17373_/A sky130_fd_sc_hd__clkbuf_4
Xfanout546 _16012_/S vssd1 vssd1 vccd1 vccd1 _14356_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_76_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09835_ _09835_/A _09835_/B vssd1 vssd1 vccd1 vccd1 _09863_/A sky130_fd_sc_hd__xnor2_1
XFILLER_86_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout557 _09899_/B vssd1 vssd1 vccd1 vccd1 _10419_/B sky130_fd_sc_hd__clkbuf_4
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout568 _11932_/A vssd1 vssd1 vccd1 vccd1 _09327_/C sky130_fd_sc_hd__buf_2
Xfanout579 _12845_/S vssd1 vssd1 vccd1 vccd1 _09493_/A sky130_fd_sc_hd__clkbuf_2
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09766_ _09776_/A _09745_/Y _09761_/A _09765_/X vssd1 vssd1 vccd1 vccd1 _09769_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_100_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08717_ _12592_/B vssd1 vssd1 vccd1 vccd1 _17377_/A sky130_fd_sc_hd__clkinv_4
XTAP_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09697_ _10241_/B _09555_/D _09843_/C _10694_/A vssd1 vssd1 vccd1 vccd1 _09699_/A
+ sky130_fd_sc_hd__a22oi_1
XTAP_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_452 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10610_ _10610_/A _10610_/B vssd1 vssd1 vccd1 vccd1 _10711_/B sky130_fd_sc_hd__xnor2_2
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11590_ _11590_/A _11590_/B vssd1 vssd1 vccd1 vccd1 _11598_/A sky130_fd_sc_hd__nor2_1
XFILLER_23_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10541_ _10545_/C _10543_/B _10434_/A _10432_/Y vssd1 vssd1 vccd1 vccd1 _10547_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_155_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13260_ _13260_/A vssd1 vssd1 vccd1 vccd1 _13261_/C sky130_fd_sc_hd__inv_2
XFILLER_157_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10472_ _10459_/A _10459_/C _10459_/B vssd1 vssd1 vccd1 vccd1 _10472_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_68_1001 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12211_ _11804_/Y _11807_/Y _17365_/A vssd1 vssd1 vccd1 vccd1 _12211_/X sky130_fd_sc_hd__mux2_1
XFILLER_136_774 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13191_ _13061_/A _13063_/A _13188_/X _13190_/Y vssd1 vssd1 vccd1 vccd1 _13332_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_68_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12142_ _11937_/A _11937_/B _11936_/A vssd1 vssd1 vccd1 vccd1 _12143_/B sky130_fd_sc_hd__a21oi_1
XFILLER_135_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16950_ _16950_/A _16950_/B vssd1 vssd1 vccd1 vccd1 _16952_/C sky130_fd_sc_hd__xor2_1
X_12073_ _11860_/A _11862_/B _11860_/B vssd1 vssd1 vccd1 vccd1 _12075_/B sky130_fd_sc_hd__o21ba_1
XFILLER_2_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11024_ _11024_/A _11024_/B _11024_/C vssd1 vssd1 vccd1 vccd1 _11041_/B sky130_fd_sc_hd__or3_1
X_15901_ _15245_/X _15253_/X _15901_/S vssd1 vssd1 vccd1 vccd1 _15901_/X sky130_fd_sc_hd__mux2_1
X_16881_ _16880_/A _16935_/B _16880_/C vssd1 vssd1 vccd1 vccd1 _16882_/B sky130_fd_sc_hd__a21oi_1
XFILLER_89_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15832_ _15832_/A _15832_/B vssd1 vssd1 vccd1 vccd1 _15834_/B sky130_fd_sc_hd__xnor2_1
XFILLER_65_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_611 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15763_ _15764_/A _15764_/B _15764_/C vssd1 vssd1 vccd1 vccd1 _15868_/B sky130_fd_sc_hd__a21oi_1
X_12975_ _13112_/A _12975_/B vssd1 vssd1 vccd1 vccd1 _12975_/X sky130_fd_sc_hd__and2_1
XFILLER_45_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17502_ fanout946/X _17502_/D vssd1 vssd1 vccd1 vccd1 _17502_/Q sky130_fd_sc_hd__dfxtp_4
X_14714_ _14713_/A _14713_/B _14713_/C vssd1 vssd1 vccd1 vccd1 _14715_/B sky130_fd_sc_hd__a21o_1
XTAP_3484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11926_ _09327_/C _17139_/A _09001_/A _08999_/B vssd1 vssd1 vccd1 vccd1 _11937_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_33_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15694_ _15595_/A _15599_/A _15786_/A _15693_/Y vssd1 vssd1 vccd1 vccd1 _15786_/B
+ sky130_fd_sc_hd__a211oi_1
XTAP_3495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17433_ input61/X _17477_/D _17433_/S vssd1 vssd1 vccd1 vccd1 _17610_/D sky130_fd_sc_hd__mux2_1
XTAP_2783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14645_ _14645_/A _14678_/B vssd1 vssd1 vccd1 vccd1 _14655_/A sky130_fd_sc_hd__nor2_1
XTAP_2794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_444 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11857_ _11785_/X _11786_/Y _11856_/X vssd1 vssd1 vccd1 vccd1 _17576_/D sky130_fd_sc_hd__o21ai_1
XFILLER_159_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10808_ _10808_/A _10808_/B vssd1 vssd1 vccd1 vccd1 _10814_/A sky130_fd_sc_hd__xnor2_1
X_17364_ input36/X _17377_/B _17363_/Y _17364_/C1 vssd1 vssd1 vccd1 vccd1 _17510_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_60_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14576_ _14577_/A _14577_/B vssd1 vssd1 vccd1 vccd1 _14627_/A sky130_fd_sc_hd__nor2_1
XFILLER_14_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11788_ _16108_/C _16317_/A vssd1 vssd1 vccd1 vccd1 _14888_/B sky130_fd_sc_hd__or2_2
X_16315_ _16315_/A _16315_/B _16315_/C _16315_/D vssd1 vssd1 vccd1 vccd1 _16316_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_159_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13527_ _13637_/B _13527_/B _13527_/C vssd1 vssd1 vccd1 vccd1 _13527_/X sky130_fd_sc_hd__and3_1
XFILLER_158_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10739_ _10739_/A _11018_/A vssd1 vssd1 vccd1 vccd1 _10747_/A sky130_fd_sc_hd__nor2_1
X_17295_ input25/X _17362_/D input28/X _17428_/C vssd1 vssd1 vccd1 vccd1 _17295_/X
+ sky130_fd_sc_hd__or4b_1
XFILLER_174_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16246_ _16760_/B _16589_/B _16246_/C vssd1 vssd1 vccd1 vccd1 _16248_/A sky130_fd_sc_hd__and3_1
XFILLER_146_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13458_ _13459_/A _13459_/B vssd1 vssd1 vccd1 vccd1 _13576_/B sky130_fd_sc_hd__nand2_1
XFILLER_174_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12409_ _12409_/A _12561_/B vssd1 vssd1 vccd1 vccd1 _12412_/A sky130_fd_sc_hd__nor2_1
X_16177_ _16177_/A _16177_/B vssd1 vssd1 vccd1 vccd1 _16179_/B sky130_fd_sc_hd__xnor2_1
Xoutput105 _17463_/Q vssd1 vssd1 vccd1 vccd1 o_wb_data[29] sky130_fd_sc_hd__clkbuf_1
XFILLER_127_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13389_ _14756_/A1 _13387_/Y _13388_/X _13274_/Y _13277_/X vssd1 vssd1 vccd1 vccd1
+ _17586_/D sky130_fd_sc_hd__a32o_1
XFILLER_126_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15128_ _15381_/A _15463_/A _10255_/B _10270_/B _10430_/A _10545_/C vssd1 vssd1 vccd1
+ vccd1 _15131_/B sky130_fd_sc_hd__mux4_1
XFILLER_99_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15059_ _15131_/A _15059_/B vssd1 vssd1 vccd1 vccd1 _15059_/Y sky130_fd_sc_hd__nand2_1
XFILLER_87_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09620_ _09620_/A _09620_/B vssd1 vssd1 vccd1 vccd1 _09621_/C sky130_fd_sc_hd__and2_1
XFILLER_28_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09551_ _09552_/A _09550_/Y _10366_/A _09985_/D vssd1 vssd1 vccd1 vccd1 _09696_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_37_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09482_ _09476_/Y _09480_/X _09460_/X _09461_/Y vssd1 vssd1 vccd1 vccd1 _09484_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_102_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_814 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout310 _17613_/Q vssd1 vssd1 vccd1 vccd1 _15147_/A sky130_fd_sc_hd__buf_2
XFILLER_120_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout321 _14290_/A vssd1 vssd1 vccd1 vccd1 _14641_/A sky130_fd_sc_hd__buf_2
Xfanout332 _08988_/B vssd1 vssd1 vccd1 vccd1 _17134_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_99_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout343 _17538_/Q vssd1 vssd1 vccd1 vccd1 _14153_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_115_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout354 _17537_/Q vssd1 vssd1 vccd1 vccd1 _14766_/A sky130_fd_sc_hd__buf_2
XFILLER_101_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout365 _14769_/A vssd1 vssd1 vccd1 vccd1 _16913_/C sky130_fd_sc_hd__buf_2
Xfanout376 fanout380/X vssd1 vssd1 vccd1 vccd1 _12787_/B sky130_fd_sc_hd__buf_2
Xfanout387 _17533_/Q vssd1 vssd1 vccd1 vccd1 _12788_/A sky130_fd_sc_hd__buf_4
X_09818_ _09828_/A _09817_/B _09814_/X vssd1 vssd1 vccd1 vccd1 _09819_/C sky130_fd_sc_hd__a21oi_1
Xfanout398 _16644_/C vssd1 vssd1 vccd1 vccd1 _13578_/A sky130_fd_sc_hd__buf_2
XFILLER_87_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09749_ _09892_/B _10299_/D _10421_/D _09892_/A vssd1 vssd1 vccd1 vccd1 _09749_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_27_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_761 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12760_ _12761_/A _12761_/B _12761_/C vssd1 vssd1 vccd1 vccd1 _12928_/A sky130_fd_sc_hd__o21a_1
XTAP_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11711_ _11711_/A _11711_/B vssd1 vssd1 vccd1 vccd1 _11713_/B sky130_fd_sc_hd__xnor2_1
XFILLER_36_98 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12691_ _12691_/A _12691_/B vssd1 vssd1 vccd1 vccd1 _12694_/A sky130_fd_sc_hd__or2_1
XTAP_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14430_ _14430_/A _14430_/B vssd1 vssd1 vccd1 vccd1 _14431_/B sky130_fd_sc_hd__and2_1
X_11642_ _15305_/C _11605_/B _11610_/B _11605_/D vssd1 vssd1 vccd1 vccd1 _11644_/C
+ sky130_fd_sc_hd__a22o_1
XTAP_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14361_ _14361_/A _14440_/A vssd1 vssd1 vccd1 vccd1 _14364_/A sky130_fd_sc_hd__or2_1
XFILLER_168_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11573_ _11534_/B _11530_/B _11530_/C vssd1 vssd1 vccd1 vccd1 _11574_/C sky130_fd_sc_hd__a21oi_1
XFILLER_167_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput18 i_wb_addr[23] vssd1 vssd1 vccd1 vccd1 input18/X sky130_fd_sc_hd__clkbuf_1
X_16100_ _16203_/A _16100_/B vssd1 vssd1 vccd1 vccd1 _16100_/Y sky130_fd_sc_hd__nor2_1
X_13312_ _13312_/A _13312_/B _13312_/C vssd1 vssd1 vccd1 vccd1 _13317_/B sky130_fd_sc_hd__or3_1
XFILLER_167_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10524_ _10524_/A _10524_/B vssd1 vssd1 vccd1 vccd1 _10540_/A sky130_fd_sc_hd__xnor2_1
XFILLER_7_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput29 i_wb_addr[4] vssd1 vssd1 vccd1 vccd1 input29/X sky130_fd_sc_hd__dlymetal6s2s_1
X_17080_ _17065_/A _17170_/B1 _17063_/Y _17079_/X vssd1 vssd1 vccd1 vccd1 _17571_/D
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_168_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14292_ _14676_/A _16859_/A vssd1 vssd1 vccd1 vccd1 _14294_/B sky130_fd_sc_hd__nand2_1
XFILLER_156_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16031_ _16129_/A _16743_/C _16136_/C vssd1 vssd1 vccd1 vccd1 _16032_/B sky130_fd_sc_hd__and3_1
X_13243_ _13243_/A _13243_/B vssd1 vssd1 vccd1 vccd1 _13244_/C sky130_fd_sc_hd__or2_1
X_10455_ _10564_/A _10456_/B vssd1 vssd1 vccd1 vccd1 _10455_/X sky130_fd_sc_hd__or2_1
XFILLER_109_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13174_ _13174_/A _13174_/B vssd1 vssd1 vccd1 vccd1 _13176_/B sky130_fd_sc_hd__xnor2_1
X_10386_ _10385_/A _10385_/Y _10262_/X _10357_/Y vssd1 vssd1 vccd1 vccd1 _10405_/A
+ sky130_fd_sc_hd__a211oi_1
XFILLER_151_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12125_ _11939_/A _11939_/B _11940_/X vssd1 vssd1 vccd1 vccd1 _12150_/A sky130_fd_sc_hd__o21ba_1
XFILLER_97_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12056_ _12049_/Y _12051_/Y _12053_/Y _12055_/Y _14948_/A _15384_/S vssd1 vssd1 vccd1
+ vccd1 _12056_/X sky130_fd_sc_hd__mux4_1
XFILLER_111_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16933_ _16933_/A _16989_/A vssd1 vssd1 vccd1 vccd1 _16933_/Y sky130_fd_sc_hd__nand2_1
XFILLER_77_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11007_ _11006_/B _10805_/D _11006_/C _11006_/A vssd1 vssd1 vccd1 vccd1 _11007_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_42_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16864_ _16864_/A _16864_/B vssd1 vssd1 vccd1 vccd1 _16865_/B sky130_fd_sc_hd__nand2_1
XFILLER_93_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15815_ _15815_/A vssd1 vssd1 vccd1 vccd1 _17555_/D sky130_fd_sc_hd__inv_2
XFILLER_19_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16795_ _16795_/A _16795_/B vssd1 vssd1 vccd1 vccd1 _16795_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_80_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15746_ _16055_/A _16681_/C vssd1 vssd1 vccd1 vccd1 _15746_/X sky130_fd_sc_hd__or2_2
XTAP_3270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12958_ _12959_/A _12959_/B vssd1 vssd1 vccd1 vccd1 _12960_/A sky130_fd_sc_hd__or2_1
XTAP_3281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11909_ _11909_/A _11909_/B vssd1 vssd1 vccd1 vccd1 _11911_/C sky130_fd_sc_hd__or2_1
X_15677_ _15572_/Y _15583_/Y _15674_/X _15676_/A vssd1 vssd1 vccd1 vccd1 _15772_/B
+ sky130_fd_sc_hd__a211o_1
X_12889_ _13414_/B _13908_/B _13802_/B _13658_/A vssd1 vssd1 vccd1 vccd1 _12889_/Y
+ sky130_fd_sc_hd__a22oi_1
XTAP_2580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17416_ input54/X _17426_/A2 _17415_/X _17422_/C1 vssd1 vssd1 vccd1 vccd1 _17536_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_33_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14628_ _14638_/A _14628_/B vssd1 vssd1 vccd1 vccd1 _14633_/A sky130_fd_sc_hd__and2_1
XFILLER_159_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17347_ input53/X _17355_/B _17355_/C vssd1 vssd1 vccd1 vccd1 _17347_/X sky130_fd_sc_hd__or3_1
XFILLER_20_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14559_ _14492_/A _14492_/B _14495_/A vssd1 vssd1 vccd1 vccd1 _14560_/B sky130_fd_sc_hd__o21ba_1
XFILLER_119_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_622 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17278_ _17460_/Q _17293_/A2 _17276_/X _17277_/X _17284_/C1 vssd1 vssd1 vccd1 vccd1
+ _17460_/D sky130_fd_sc_hd__o221a_1
X_16229_ _16229_/A _16229_/B vssd1 vssd1 vccd1 vccd1 _16232_/A sky130_fd_sc_hd__xor2_1
XFILLER_114_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08982_ _08983_/A _08983_/B vssd1 vssd1 vccd1 vccd1 _09242_/B sky130_fd_sc_hd__nand2_1
XFILLER_115_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09603_ _09603_/A _09603_/B vssd1 vssd1 vccd1 vccd1 _09618_/A sky130_fd_sc_hd__nand2_1
XFILLER_28_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09534_ _09531_/X _09540_/A _12005_/B _09397_/X vssd1 vssd1 vccd1 vccd1 _09536_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_58_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09465_ _09892_/B _10543_/B _10545_/D _09892_/A vssd1 vssd1 vccd1 vccd1 _09465_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_24_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09396_ _09343_/X _09393_/B _12005_/A _09395_/X vssd1 vssd1 vccd1 vccd1 _12005_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_51_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10240_ _10246_/A _10246_/B vssd1 vssd1 vccd1 vccd1 _10261_/B sky130_fd_sc_hd__nand2_1
XFILLER_145_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1015 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10171_ _14789_/A _10419_/B _10299_/D _10171_/D vssd1 vssd1 vccd1 vccd1 _10288_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_160_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout140 _16086_/A vssd1 vssd1 vccd1 vccd1 _16281_/A sky130_fd_sc_hd__clkbuf_4
Xfanout151 _15100_/A vssd1 vssd1 vccd1 vccd1 _15102_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout162 _17361_/Y vssd1 vssd1 vccd1 vccd1 _17389_/B sky130_fd_sc_hd__buf_2
X_13930_ _13930_/A _13930_/B vssd1 vssd1 vccd1 vccd1 _13932_/B sky130_fd_sc_hd__nor2_1
Xfanout173 _16743_/B vssd1 vssd1 vccd1 vccd1 _16259_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_75_823 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout184 _16334_/A vssd1 vssd1 vccd1 vccd1 _16814_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_87_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout195 _16582_/A vssd1 vssd1 vccd1 vccd1 _17164_/C sky130_fd_sc_hd__buf_2
XFILLER_47_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13861_ _13861_/A _13861_/B _13861_/C vssd1 vssd1 vccd1 vccd1 _13862_/C sky130_fd_sc_hd__nand3_1
XFILLER_47_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15600_ _15601_/A _15601_/B vssd1 vssd1 vccd1 vccd1 _15600_/Y sky130_fd_sc_hd__nor2_1
X_12812_ _12812_/A _12812_/B vssd1 vssd1 vccd1 vccd1 _12976_/A sky130_fd_sc_hd__xor2_1
XFILLER_90_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16580_ _16576_/B _17162_/A2 _16580_/B1 _16571_/A _17162_/C1 vssd1 vssd1 vccd1 vccd1
+ _16580_/X sky130_fd_sc_hd__a221o_1
X_13792_ _13792_/A _13792_/B vssd1 vssd1 vccd1 vccd1 _13793_/C sky130_fd_sc_hd__xnor2_1
X_15531_ _15529_/Y _15620_/A vssd1 vssd1 vccd1 vccd1 _15533_/A sky130_fd_sc_hd__and2b_1
XFILLER_27_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12743_ _12902_/A _12743_/B _12743_/C vssd1 vssd1 vccd1 vccd1 _12902_/B sky130_fd_sc_hd__nand3_1
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15462_ _15458_/Y _15459_/Y _15461_/Y vssd1 vssd1 vccd1 vccd1 _15462_/Y sky130_fd_sc_hd__o21ai_1
X_12674_ _12675_/B _12675_/A vssd1 vssd1 vccd1 vccd1 _12674_/Y sky130_fd_sc_hd__nand2b_1
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17201_ _17576_/Q _17273_/A2 _17273_/B1 vssd1 vssd1 vccd1 vccd1 _17201_/X sky130_fd_sc_hd__a21o_1
X_14413_ _14413_/A _14413_/B _14413_/C vssd1 vssd1 vccd1 vccd1 _14414_/B sky130_fd_sc_hd__nor3_1
X_11625_ _11617_/B _11617_/C _11617_/A vssd1 vssd1 vccd1 vccd1 _11672_/B sky130_fd_sc_hd__o21ai_1
X_15393_ _15393_/A _15393_/B vssd1 vssd1 vccd1 vccd1 _15396_/B sky130_fd_sc_hd__nand2_1
XFILLER_128_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_622 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17132_ _17134_/A _16965_/B _17134_/B vssd1 vssd1 vccd1 vccd1 _17133_/A sky130_fd_sc_hd__a21o_1
X_14344_ _14344_/A _14344_/B _14344_/C vssd1 vssd1 vccd1 vccd1 _14345_/B sky130_fd_sc_hd__nor3_1
X_11556_ _11512_/A _11512_/C _11512_/B vssd1 vssd1 vccd1 vccd1 _11558_/C sky130_fd_sc_hd__a21o_1
XFILLER_155_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10507_ _10963_/B _10736_/D _10875_/C _10963_/A vssd1 vssd1 vccd1 vccd1 _10507_/Y
+ sky130_fd_sc_hd__a22oi_1
X_17063_ _17063_/A _17063_/B vssd1 vssd1 vccd1 vccd1 _17063_/Y sky130_fd_sc_hd__nor2_2
XFILLER_10_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14275_ _14276_/A _14276_/B _14274_/X vssd1 vssd1 vccd1 vccd1 _14352_/A sky130_fd_sc_hd__o21ba_1
X_11487_ _11487_/A _11487_/B _11485_/X vssd1 vssd1 vccd1 vccd1 _11527_/A sky130_fd_sc_hd__nor3b_2
XFILLER_143_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_571 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16014_ _16014_/A _16014_/B vssd1 vssd1 vccd1 vccd1 _16015_/C sky130_fd_sc_hd__nor2_1
X_13226_ _14153_/B _13664_/D _13551_/D _13227_/A vssd1 vssd1 vccd1 vccd1 _13228_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_124_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10438_ _10453_/A _10410_/Y _10425_/Y _10437_/X vssd1 vssd1 vccd1 vccd1 _10440_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_98_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13157_ _13157_/A _13157_/B vssd1 vssd1 vccd1 vccd1 _13159_/A sky130_fd_sc_hd__nor2_1
XFILLER_69_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10369_ _10484_/A _10369_/B vssd1 vssd1 vccd1 vccd1 _10383_/B sky130_fd_sc_hd__nand2_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12108_ _12108_/A _12108_/B vssd1 vssd1 vccd1 vccd1 _12110_/A sky130_fd_sc_hd__nor2_1
XFILLER_2_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13088_ _13903_/A _13966_/C _13088_/C vssd1 vssd1 vccd1 vccd1 _13220_/B sky130_fd_sc_hd__nand3_1
XFILLER_97_469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16916_ _16916_/A _16916_/B vssd1 vssd1 vccd1 vccd1 _16917_/B sky130_fd_sc_hd__xnor2_1
X_12039_ _17306_/A1 _17304_/A1 _14942_/A vssd1 vssd1 vccd1 vccd1 _12040_/B sky130_fd_sc_hd__mux2_1
XFILLER_111_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16847_ _16909_/A _16847_/B vssd1 vssd1 vccd1 vccd1 _16848_/A sky130_fd_sc_hd__nand2_1
XFILLER_92_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16778_ _16846_/A _16778_/B vssd1 vssd1 vccd1 vccd1 _16781_/A sky130_fd_sc_hd__or2_1
XFILLER_129_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15729_ _15730_/A _15730_/B vssd1 vssd1 vccd1 vccd1 _15827_/A sky130_fd_sc_hd__nand2_1
XFILLER_61_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09250_ _09115_/A _09114_/Y _09248_/Y _09249_/X vssd1 vssd1 vccd1 vccd1 _09250_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_22_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09181_ _09179_/A _09346_/A _09155_/Y _09156_/X vssd1 vssd1 vccd1 vccd1 _09214_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_21_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_614 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_48 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_511 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_447 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_224 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08965_ _09493_/A _11932_/B vssd1 vssd1 vccd1 vccd1 _08965_/Y sky130_fd_sc_hd__nand2_1
XFILLER_97_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08896_ _17389_/A _12500_/B vssd1 vssd1 vccd1 vccd1 _09043_/A sky130_fd_sc_hd__nand2_1
XFILLER_84_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_12 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09517_ _09517_/A _09636_/A vssd1 vssd1 vccd1 vccd1 _09519_/B sky130_fd_sc_hd__nor2_1
XFILLER_25_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09448_ _09449_/B _09449_/A vssd1 vssd1 vccd1 vccd1 _09448_/X sky130_fd_sc_hd__and2b_1
XPHY_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09379_ _09379_/A _09513_/A vssd1 vssd1 vccd1 vccd1 _09381_/B sky130_fd_sc_hd__nor2_1
XFILLER_8_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11410_ _11411_/A _11411_/B vssd1 vssd1 vccd1 vccd1 _11410_/Y sky130_fd_sc_hd__nor2_1
XFILLER_21_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12390_ _12026_/Y _12031_/Y _14948_/A vssd1 vssd1 vccd1 vccd1 _12390_/X sky130_fd_sc_hd__mux2_1
XFILLER_123_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11341_ _11341_/A _11341_/B _11341_/C vssd1 vssd1 vccd1 vccd1 _11367_/A sky130_fd_sc_hd__and3_1
XFILLER_138_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14060_ _14060_/A _14060_/B vssd1 vssd1 vccd1 vccd1 _14104_/A sky130_fd_sc_hd__xnor2_1
X_11272_ _11274_/B _11274_/C _11274_/A vssd1 vssd1 vccd1 vccd1 _11272_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_134_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13011_ _16922_/A _13009_/Y _13138_/B _12860_/Y _12867_/X vssd1 vssd1 vccd1 vccd1
+ _17583_/D sky130_fd_sc_hd__a32o_1
XFILLER_79_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10223_ _10223_/A _10223_/B vssd1 vssd1 vccd1 vccd1 _10226_/B sky130_fd_sc_hd__xnor2_1
XFILLER_134_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10154_ _10137_/X _10138_/Y _10149_/A _10152_/X vssd1 vssd1 vccd1 vccd1 _10155_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_121_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14962_ _14962_/A _14962_/B vssd1 vssd1 vccd1 vccd1 _15386_/A sky130_fd_sc_hd__nor2_1
XFILLER_59_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10085_ _10059_/A _10059_/B _10059_/C vssd1 vssd1 vccd1 vccd1 _10086_/C sky130_fd_sc_hd__o21a_1
XFILLER_87_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16701_ _16701_/A _16701_/B vssd1 vssd1 vccd1 vccd1 _16702_/B sky130_fd_sc_hd__nand2_1
XFILLER_59_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13913_ _14013_/B _13913_/B vssd1 vssd1 vccd1 vccd1 _13915_/C sky130_fd_sc_hd__and2_1
X_14893_ _16938_/A _14893_/B vssd1 vssd1 vccd1 vccd1 _14967_/C sky130_fd_sc_hd__or2_1
XFILLER_63_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16632_ _16543_/A _16543_/B _16544_/X vssd1 vssd1 vccd1 vccd1 _16634_/B sky130_fd_sc_hd__a21oi_1
X_13844_ _13948_/A _13948_/B _13844_/C _14008_/B vssd1 vssd1 vccd1 vccd1 _13954_/A
+ sky130_fd_sc_hd__and4_1
Xwb_buttons_leds_970 vssd1 vssd1 vccd1 vccd1 wb_buttons_leds_970/HI o_wb_stall sky130_fd_sc_hd__conb_1
XFILLER_90_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16563_ _16563_/A _16563_/B vssd1 vssd1 vccd1 vccd1 _16564_/B sky130_fd_sc_hd__nor2_1
X_13775_ _14155_/A _14213_/D vssd1 vssd1 vccd1 vccd1 _13776_/B sky130_fd_sc_hd__nand2_1
X_10987_ _10987_/A _10987_/B vssd1 vssd1 vccd1 vccd1 _10990_/C sky130_fd_sc_hd__xnor2_1
XFILLER_15_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12726_ _12727_/A _12727_/B vssd1 vssd1 vccd1 vccd1 _12886_/B sky130_fd_sc_hd__and2_1
X_15514_ _15514_/A _15514_/B _15514_/C vssd1 vssd1 vccd1 vccd1 _15515_/B sky130_fd_sc_hd__and3_1
X_16494_ _16475_/X _16478_/X _16493_/X _16494_/B1 _16480_/A vssd1 vssd1 vccd1 vccd1
+ _16495_/A sky130_fd_sc_hd__a32o_1
XFILLER_90_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15445_ _15442_/Y _15443_/X _15444_/Y vssd1 vssd1 vccd1 vccd1 _15445_/X sky130_fd_sc_hd__a21o_1
X_12657_ _12804_/A _12804_/B _13194_/D _13067_/D vssd1 vssd1 vccd1 vccd1 _12658_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_129_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11608_ _11607_/A _11607_/C _11607_/B vssd1 vssd1 vccd1 vccd1 _11612_/B sky130_fd_sc_hd__a21o_1
XFILLER_12_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15376_ _15374_/X _15375_/X _16111_/A vssd1 vssd1 vccd1 vccd1 _15376_/Y sky130_fd_sc_hd__a21oi_1
X_12588_ _12588_/A _12588_/B _12588_/C vssd1 vssd1 vccd1 vccd1 _12612_/B sky130_fd_sc_hd__and3_1
X_17115_ _17063_/A _17096_/Y _17097_/X _17114_/X vssd1 vssd1 vccd1 vccd1 _17115_/X
+ sky130_fd_sc_hd__o31a_1
X_14327_ _16723_/A _14450_/B _14326_/C vssd1 vssd1 vccd1 vccd1 _14328_/B sky130_fd_sc_hd__a21o_1
XFILLER_172_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11539_ _11539_/A _11539_/B _11538_/X vssd1 vssd1 vccd1 vccd1 _11542_/A sky130_fd_sc_hd__nor3b_1
XFILLER_7_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17046_ _17046_/A _17046_/B _17046_/C vssd1 vssd1 vccd1 vccd1 _17047_/B sky130_fd_sc_hd__nor3_1
X_14258_ _14258_/A _14258_/B vssd1 vssd1 vccd1 vccd1 _14258_/X sky130_fd_sc_hd__or2_1
XFILLER_99_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13209_ _13897_/A _13966_/C vssd1 vssd1 vccd1 vccd1 _13211_/C sky130_fd_sc_hd__nand2_1
XFILLER_48_1043 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14189_ _14268_/A _14189_/B vssd1 vssd1 vccd1 vccd1 _14190_/B sky130_fd_sc_hd__nor2_1
XFILLER_124_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout909 _11095_/D vssd1 vssd1 vccd1 vccd1 _17466_/D sky130_fd_sc_hd__clkbuf_4
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1046 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08750_ _08750_/A _08750_/B vssd1 vssd1 vccd1 vccd1 _08757_/A sky130_fd_sc_hd__xnor2_4
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_303 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09302_ _09302_/A _09443_/A vssd1 vssd1 vccd1 vccd1 _09304_/B sky130_fd_sc_hd__nor2_1
XFILLER_62_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09233_ _12804_/A _12804_/B _12129_/B _12127_/C vssd1 vssd1 vccd1 vccd1 _09234_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_148_942 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09164_ _09164_/A _09354_/A vssd1 vssd1 vccd1 vccd1 _09168_/B sky130_fd_sc_hd__nor2_1
XFILLER_119_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09095_ _09095_/A _09095_/B vssd1 vssd1 vccd1 vccd1 _09103_/A sky130_fd_sc_hd__nor2_1
XFILLER_107_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_850 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_511 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09997_ _10254_/A _11790_/A _10508_/D _10255_/B vssd1 vssd1 vccd1 vccd1 _10000_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_131_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08948_ _08947_/B _11900_/D _12256_/D _09078_/A vssd1 vssd1 vccd1 vccd1 _08948_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_76_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_34 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_66 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08879_ _12068_/A _17399_/A _09272_/D _12338_/C vssd1 vssd1 vccd1 vccd1 _08882_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_57_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10910_ _11107_/A _11073_/B vssd1 vssd1 vccd1 vccd1 _11074_/A sky130_fd_sc_hd__nand2_1
XFILLER_85_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11890_ _11891_/A _11891_/B _11891_/C vssd1 vssd1 vccd1 vccd1 _11890_/X sky130_fd_sc_hd__o21a_1
XFILLER_45_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10841_ _10841_/A _10841_/B vssd1 vssd1 vccd1 vccd1 _10842_/B sky130_fd_sc_hd__nor2_1
XFILLER_44_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13560_ _13443_/B _13444_/Y _13557_/Y _13559_/A vssd1 vssd1 vccd1 vccd1 _13562_/A
+ sky130_fd_sc_hd__a211oi_2
XFILLER_44_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10772_ _10777_/A _10772_/B vssd1 vssd1 vccd1 vccd1 _10774_/B sky130_fd_sc_hd__nand2_1
XFILLER_13_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12511_ _12511_/A _12511_/B vssd1 vssd1 vccd1 vccd1 _12514_/A sky130_fd_sc_hd__xor2_1
XFILLER_12_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13491_ _13607_/A _13490_/B _13490_/C _13490_/D vssd1 vssd1 vccd1 vccd1 _13492_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_40_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15230_ _15230_/A _15230_/B vssd1 vssd1 vccd1 vccd1 _15231_/B sky130_fd_sc_hd__nand2_1
XFILLER_139_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12442_ _12442_/A _12592_/C _12442_/C vssd1 vssd1 vccd1 vccd1 _12616_/B sky130_fd_sc_hd__and3_1
XFILLER_139_975 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15161_ _15161_/A _15161_/B vssd1 vssd1 vccd1 vccd1 _15162_/B sky130_fd_sc_hd__nand2_1
X_12373_ _12373_/A _12373_/B vssd1 vssd1 vccd1 vccd1 _12696_/A sky130_fd_sc_hd__xnor2_1
XFILLER_138_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14112_ _14113_/A _14113_/B _14113_/C vssd1 vssd1 vccd1 vccd1 _14202_/A sky130_fd_sc_hd__a21o_1
X_11324_ _11553_/B _11518_/C _11325_/A _11324_/D vssd1 vssd1 vccd1 vccd1 _11376_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_4_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15092_ _15170_/A _15170_/B vssd1 vssd1 vccd1 vccd1 _15094_/A sky130_fd_sc_hd__nand2_1
XFILLER_158_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_988 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14043_ _14043_/A _14043_/B vssd1 vssd1 vccd1 vccd1 _14134_/B sky130_fd_sc_hd__xnor2_2
X_11255_ _11255_/A _11255_/B _11255_/C vssd1 vssd1 vccd1 vccd1 _11291_/A sky130_fd_sc_hd__or3_1
XFILLER_122_820 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10206_ _10331_/A _10331_/B vssd1 vssd1 vccd1 vccd1 _10212_/A sky130_fd_sc_hd__and2b_1
X_11186_ _11202_/B _11186_/B _11218_/A _11186_/D vssd1 vssd1 vccd1 vccd1 _11218_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_122_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10137_ _10138_/A _10138_/B _10138_/C vssd1 vssd1 vccd1 vccd1 _10137_/X sky130_fd_sc_hd__a21o_1
XFILLER_121_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15994_ _15994_/A _15994_/B vssd1 vssd1 vccd1 vccd1 _15994_/X sky130_fd_sc_hd__and2_1
X_10068_ _10069_/B _10200_/A _10069_/A vssd1 vssd1 vccd1 vccd1 _10070_/A sky130_fd_sc_hd__o21ai_1
X_14945_ _15237_/A1 _15457_/B _14841_/B _14944_/Y vssd1 vssd1 vccd1 vccd1 _14945_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_35_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14876_ _15396_/A _14888_/C _14876_/C _14876_/D vssd1 vssd1 vccd1 vccd1 _14876_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_62_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16615_ _16616_/A _16616_/B _16616_/C vssd1 vssd1 vccd1 vccd1 _16617_/A sky130_fd_sc_hd__o21a_1
X_13827_ _13827_/A _13827_/B vssd1 vssd1 vccd1 vccd1 _13936_/B sky130_fd_sc_hd__xor2_1
XFILLER_90_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17595_ fanout933/X _17595_/D vssd1 vssd1 vccd1 vccd1 _17595_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16546_ _16547_/A _16547_/B vssd1 vssd1 vccd1 vccd1 _16630_/B sky130_fd_sc_hd__nand2_1
X_13758_ _13862_/A _13758_/B vssd1 vssd1 vccd1 vccd1 _13761_/A sky130_fd_sc_hd__or2_1
XFILLER_16_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12709_ _13627_/S _12709_/B vssd1 vssd1 vccd1 vccd1 _12710_/B sky130_fd_sc_hd__or2_1
X_16477_ _11200_/Y _11229_/Y _16389_/C _16207_/B vssd1 vssd1 vccd1 vccd1 _16478_/B
+ sky130_fd_sc_hd__a31o_1
X_13689_ _13689_/A _16789_/A vssd1 vssd1 vccd1 vccd1 _16796_/A sky130_fd_sc_hd__nand2_2
XFILLER_86_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15428_ _15428_/A _15428_/B _15429_/B vssd1 vssd1 vccd1 vccd1 _15428_/X sky130_fd_sc_hd__and3_1
X_15359_ _15359_/A _15359_/B vssd1 vssd1 vccd1 vccd1 _15362_/A sky130_fd_sc_hd__xor2_1
XFILLER_156_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09920_ _09920_/A _09920_/B vssd1 vssd1 vccd1 vccd1 _09922_/B sky130_fd_sc_hd__and2_1
XFILLER_160_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17029_ _17140_/A _17029_/B _17029_/C vssd1 vssd1 vccd1 vccd1 _17033_/B sky130_fd_sc_hd__or3_1
XFILLER_116_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout706 _17499_/Q vssd1 vssd1 vccd1 vccd1 _12088_/D sky130_fd_sc_hd__clkbuf_4
Xfanout717 _13966_/C vssd1 vssd1 vccd1 vccd1 _14050_/D sky130_fd_sc_hd__clkbuf_4
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09851_ _09845_/B _09847_/B _09845_/A vssd1 vssd1 vccd1 vccd1 _09854_/A sky130_fd_sc_hd__o21ba_1
Xfanout728 _17496_/Q vssd1 vssd1 vccd1 vccd1 _16399_/A sky130_fd_sc_hd__buf_4
XFILLER_59_918 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout739 _11841_/B vssd1 vssd1 vccd1 vccd1 _10421_/D sky130_fd_sc_hd__buf_2
X_08802_ _08802_/A _08802_/B vssd1 vssd1 vccd1 vccd1 _08831_/A sky130_fd_sc_hd__xnor2_1
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09782_ _09783_/A _09781_/Y _10182_/C _09926_/B vssd1 vssd1 vccd1 vccd1 _09930_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_85_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08733_ _17476_/D _17477_/D vssd1 vssd1 vccd1 vccd1 _08733_/Y sky130_fd_sc_hd__nand2_1
XFILLER_22_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_564 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09216_ _17413_/A _17411_/A _09555_/D _12338_/D vssd1 vssd1 vccd1 vccd1 _11958_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_22_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09147_ _09148_/A _09147_/B _09231_/B vssd1 vssd1 vccd1 vccd1 _09245_/A sky130_fd_sc_hd__or3_1
XFILLER_107_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09078_ _09078_/A _11895_/B _12256_/D _12088_/D vssd1 vssd1 vccd1 vccd1 _09081_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_146_34 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11040_ _11046_/A _11040_/B vssd1 vssd1 vccd1 vccd1 _11041_/C sky130_fd_sc_hd__xnor2_1
XFILLER_131_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12991_ _12991_/A _12991_/B vssd1 vssd1 vccd1 vccd1 _12991_/X sky130_fd_sc_hd__or2_1
XTAP_3611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11942_ _08868_/X _08873_/C _11940_/X _11941_/Y vssd1 vssd1 vccd1 vccd1 _12156_/A
+ sky130_fd_sc_hd__a211o_1
X_14730_ _14731_/A _14731_/B vssd1 vssd1 vccd1 vccd1 _14730_/Y sky130_fd_sc_hd__nand2_1
XFILLER_57_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14661_ _14661_/A _14662_/A vssd1 vssd1 vccd1 vccd1 _14698_/B sky130_fd_sc_hd__nand2_1
XTAP_2954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11873_ _11874_/A _11874_/B vssd1 vssd1 vccd1 vccd1 _12085_/B sky130_fd_sc_hd__nand2_1
XTAP_2965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13612_ _13612_/A _13612_/B vssd1 vssd1 vccd1 vccd1 _13614_/A sky130_fd_sc_hd__nor2_1
XFILLER_44_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16400_ _16579_/A _16400_/B _16400_/C vssd1 vssd1 vccd1 vccd1 _16404_/A sky130_fd_sc_hd__or3_1
X_10824_ _11117_/C _10962_/B vssd1 vssd1 vccd1 vccd1 _10828_/A sky130_fd_sc_hd__nand2_1
XTAP_2987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17380_ input66/X _17424_/A2 _17379_/X _17388_/C1 vssd1 vssd1 vccd1 vccd1 _17518_/D
+ sky130_fd_sc_hd__o211a_1
X_14592_ _14708_/B _14433_/B _14593_/D _14738_/A vssd1 vssd1 vccd1 vccd1 _14594_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_13_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16331_ _16331_/A _16331_/B vssd1 vssd1 vccd1 vccd1 _16344_/A sky130_fd_sc_hd__xor2_1
X_13543_ _13543_/A _13543_/B vssd1 vssd1 vccd1 vccd1 _13545_/C sky130_fd_sc_hd__xnor2_1
X_10755_ _10756_/A _10754_/Y _10993_/C _11841_/B vssd1 vssd1 vccd1 vccd1 _11165_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_9_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16262_ _16262_/A _16681_/C _16262_/C vssd1 vssd1 vccd1 vccd1 _16358_/B sky130_fd_sc_hd__nor3_1
X_13474_ _13353_/A _13355_/B _13353_/B vssd1 vssd1 vccd1 vccd1 _13476_/B sky130_fd_sc_hd__o21ba_1
X_10686_ _10579_/B _10584_/X _10685_/B _10688_/A vssd1 vssd1 vccd1 vccd1 _11768_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_139_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_912 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15213_ _15846_/A _16127_/A _15213_/C vssd1 vssd1 vccd1 vccd1 _15213_/X sky130_fd_sc_hd__and3_1
XFILLER_139_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12425_ _12425_/A _12425_/B vssd1 vssd1 vccd1 vccd1 _12427_/A sky130_fd_sc_hd__nor2_1
XFILLER_173_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16193_ _16089_/A _16089_/B _16081_/A vssd1 vssd1 vccd1 vccd1 _16195_/B sky130_fd_sc_hd__o21a_1
XFILLER_126_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15144_ _11790_/X _14877_/Y _15270_/B _15143_/C _15147_/D vssd1 vssd1 vccd1 vccd1
+ _15144_/X sky130_fd_sc_hd__a2111o_1
X_12356_ _12357_/B _12357_/A vssd1 vssd1 vccd1 vccd1 _12356_/X sky130_fd_sc_hd__and2b_1
XFILLER_126_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11307_ _11364_/A _11364_/B vssd1 vssd1 vccd1 vccd1 _11399_/A sky130_fd_sc_hd__nand2_1
XFILLER_153_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15075_ _17119_/A _15147_/C vssd1 vssd1 vccd1 vccd1 _15075_/X sky130_fd_sc_hd__and2_1
XFILLER_5_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12287_ _12112_/X _12116_/A _12476_/A _12286_/Y vssd1 vssd1 vccd1 vccd1 _12476_/B
+ sky130_fd_sc_hd__o211ai_2
X_14026_ _14027_/A _14027_/B _14025_/Y vssd1 vssd1 vccd1 vccd1 _14119_/B sky130_fd_sc_hd__o21ba_1
X_11238_ _11238_/A _11238_/B vssd1 vssd1 vccd1 vccd1 _11249_/A sky130_fd_sc_hd__xor2_1
XFILLER_171_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11169_ _11168_/A _11168_/B _11167_/X vssd1 vssd1 vccd1 vccd1 _11169_/X sky130_fd_sc_hd__o21ba_1
XFILLER_67_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15977_ _16165_/A _16165_/B _15850_/A _15848_/A vssd1 vssd1 vccd1 vccd1 _15980_/C
+ sky130_fd_sc_hd__a31o_1
XFILLER_83_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14928_ _14929_/A _14933_/B vssd1 vssd1 vccd1 vccd1 _14928_/Y sky130_fd_sc_hd__nor2_1
XFILLER_48_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14859_ _16298_/A _14859_/B _16115_/B vssd1 vssd1 vccd1 vccd1 _16399_/B sky130_fd_sc_hd__and3_1
XFILLER_35_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17578_ fanout938/X _17578_/D vssd1 vssd1 vccd1 vccd1 _17578_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16529_ _16454_/A _16454_/B _16452_/Y vssd1 vssd1 vccd1 vccd1 _16545_/A sky130_fd_sc_hd__a21bo_1
XFILLER_149_536 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09001_ _09001_/A _09001_/B vssd1 vssd1 vccd1 vccd1 _09003_/B sky130_fd_sc_hd__xnor2_1
XFILLER_160_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09903_ _10034_/A _10042_/A _10034_/C vssd1 vssd1 vccd1 vccd1 _10035_/A sky130_fd_sc_hd__o21ai_1
XFILLER_104_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout503 _17519_/Q vssd1 vssd1 vccd1 vccd1 _10271_/A sky130_fd_sc_hd__buf_4
Xfanout514 _09892_/B vssd1 vssd1 vccd1 vccd1 _11895_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_116_48 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout525 _17516_/Q vssd1 vssd1 vccd1 vccd1 _12442_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_86_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout536 _12471_/A vssd1 vssd1 vccd1 vccd1 _09755_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_76_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout547 _14421_/S vssd1 vssd1 vccd1 vccd1 _16012_/S sky130_fd_sc_hd__clkbuf_4
X_09834_ _09866_/A _09866_/B vssd1 vssd1 vccd1 vccd1 _09884_/A sky130_fd_sc_hd__nand2_1
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout558 _10851_/B vssd1 vssd1 vccd1 vccd1 _11122_/B sky130_fd_sc_hd__buf_2
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_171 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout569 _15538_/A vssd1 vssd1 vccd1 vccd1 _11932_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_86_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09765_ _09765_/A _09765_/B _09765_/C vssd1 vssd1 vccd1 vccd1 _09765_/X sky130_fd_sc_hd__and3_1
XFILLER_73_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09696_ _09696_/A _09696_/B _09703_/B vssd1 vssd1 vccd1 vccd1 _09718_/B sky130_fd_sc_hd__or3_1
XTAP_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_818 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10540_ _10540_/A _10540_/B _10540_/C vssd1 vssd1 vccd1 vccd1 _10550_/B sky130_fd_sc_hd__nand3_1
XFILLER_41_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10471_ _10463_/A _10461_/X _10454_/A _10455_/X vssd1 vssd1 vccd1 vccd1 _10471_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_10_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12210_ _12374_/B _12210_/B vssd1 vssd1 vccd1 vccd1 _12210_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_108_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13190_ _13189_/A _13189_/B _13189_/C vssd1 vssd1 vccd1 vccd1 _13190_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_68_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12141_ _12141_/A _12141_/B vssd1 vssd1 vccd1 vccd1 _12143_/A sky130_fd_sc_hd__xnor2_1
XFILLER_68_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12072_ _12239_/B _12072_/B vssd1 vssd1 vccd1 vccd1 _12075_/A sky130_fd_sc_hd__nor2_1
XFILLER_96_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11023_ _11024_/A _11024_/B _11024_/C vssd1 vssd1 vccd1 vccd1 _11041_/A sky130_fd_sc_hd__o21ai_2
X_15900_ _09424_/X _17075_/A2 _15899_/X vssd1 vssd1 vccd1 vccd1 _15900_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_150_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16880_ _16880_/A _16935_/B _16880_/C vssd1 vssd1 vccd1 vccd1 _16882_/A sky130_fd_sc_hd__and3_1
XFILLER_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15831_ _15829_/X _15831_/B vssd1 vssd1 vccd1 vccd1 _15832_/B sky130_fd_sc_hd__and2b_1
XFILLER_66_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15762_ _15762_/A _15762_/B vssd1 vssd1 vccd1 vccd1 _15764_/C sky130_fd_sc_hd__xnor2_1
X_12974_ _12974_/A _12974_/B vssd1 vssd1 vccd1 vccd1 _12975_/B sky130_fd_sc_hd__nand2_1
XFILLER_66_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17501_ fanout946/X _17501_/D vssd1 vssd1 vccd1 vccd1 _17501_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14713_ _14713_/A _14713_/B _14713_/C vssd1 vssd1 vccd1 vccd1 _14742_/A sky130_fd_sc_hd__nand3_1
XTAP_3474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11925_ _12179_/B _11925_/B vssd1 vssd1 vccd1 vccd1 _11941_/A sky130_fd_sc_hd__nor2_1
XTAP_3485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15693_ _15779_/B _15691_/Y _15591_/A _15600_/Y vssd1 vssd1 vccd1 vccd1 _15693_/Y
+ sky130_fd_sc_hd__a211oi_1
XTAP_3496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17432_ input58/X _17476_/D _17433_/S vssd1 vssd1 vccd1 vccd1 _17609_/D sky130_fd_sc_hd__mux2_1
XFILLER_61_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11856_ _11849_/A _11845_/X _13625_/B _11855_/X vssd1 vssd1 vccd1 vccd1 _11856_/X
+ sky130_fd_sc_hd__a211o_1
X_14644_ _14676_/A _14708_/D _14644_/C vssd1 vssd1 vccd1 vccd1 _14678_/B sky130_fd_sc_hd__and3_1
XTAP_2784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10807_ _10807_/A _10807_/B vssd1 vssd1 vccd1 vccd1 _10808_/B sky130_fd_sc_hd__nor2_1
XFILLER_32_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17363_ _17363_/A _17377_/B vssd1 vssd1 vccd1 vccd1 _17363_/Y sky130_fd_sc_hd__nand2_1
X_14575_ _14624_/A _14575_/B vssd1 vssd1 vccd1 vccd1 _14577_/B sky130_fd_sc_hd__nand2_1
X_11787_ _15396_/A _15373_/C vssd1 vssd1 vccd1 vccd1 _14888_/A sky130_fd_sc_hd__or2_1
XFILLER_60_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16314_ _15647_/A _17119_/C _16695_/B _16226_/C vssd1 vssd1 vccd1 vccd1 _16316_/A
+ sky130_fd_sc_hd__a22o_1
X_10738_ _10739_/A _10737_/Y _11117_/C _10933_/D vssd1 vssd1 vccd1 vccd1 _11018_/A
+ sky130_fd_sc_hd__and4bb_1
X_13526_ _13526_/A _13526_/B vssd1 vssd1 vccd1 vccd1 _13527_/C sky130_fd_sc_hd__nand2_1
XFILLER_159_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17294_ input35/X input68/X input69/X vssd1 vssd1 vccd1 vccd1 _17362_/D sky130_fd_sc_hd__nand3_2
XFILLER_12_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16245_ _16245_/A _16245_/B vssd1 vssd1 vccd1 vccd1 _16246_/C sky130_fd_sc_hd__xor2_1
X_13457_ _13457_/A _13576_/A vssd1 vssd1 vccd1 vccd1 _13459_/B sky130_fd_sc_hd__and2_1
XFILLER_12_1023 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10669_ _10669_/A _10669_/B _10661_/A vssd1 vssd1 vccd1 vccd1 _10769_/A sky130_fd_sc_hd__or3b_1
XFILLER_139_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12408_ _12871_/A _13208_/C _12408_/C vssd1 vssd1 vccd1 vccd1 _12561_/B sky130_fd_sc_hd__and3_1
X_16176_ _16177_/A _16177_/B vssd1 vssd1 vccd1 vccd1 _16279_/B sky130_fd_sc_hd__and2b_1
X_13388_ _13508_/B _13388_/B vssd1 vssd1 vccd1 vccd1 _13388_/X sky130_fd_sc_hd__or2_1
XFILLER_142_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput106 _17436_/Q vssd1 vssd1 vccd1 vccd1 o_wb_data[2] sky130_fd_sc_hd__clkbuf_1
XFILLER_115_915 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_723 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12339_ _12339_/A _12339_/B vssd1 vssd1 vccd1 vccd1 _12341_/A sky130_fd_sc_hd__nor2_1
X_15127_ _15126_/A _15125_/Y _15126_/Y vssd1 vssd1 vccd1 vccd1 _15711_/B sky130_fd_sc_hd__o21ai_1
XFILLER_142_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15058_ _15624_/A _15709_/A _15811_/A _15898_/A _15058_/S0 _14954_/A vssd1 vssd1
+ vccd1 vccd1 _15059_/B sky130_fd_sc_hd__mux4_1
XFILLER_99_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14009_ _14254_/A _14008_/B _14008_/C vssd1 vssd1 vccd1 vccd1 _14010_/B sky130_fd_sc_hd__a21o_1
XFILLER_141_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_620 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09550_ _10236_/B _09843_/D _09838_/C _10236_/A vssd1 vssd1 vccd1 vccd1 _09550_/Y
+ sky130_fd_sc_hd__a22oi_1
X_09481_ _09460_/X _09461_/Y _09476_/Y _09480_/X vssd1 vssd1 vccd1 vccd1 _09484_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_70_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_773 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout300 _17369_/A vssd1 vssd1 vccd1 vccd1 _13833_/S sky130_fd_sc_hd__clkbuf_4
Xfanout311 _17612_/Q vssd1 vssd1 vccd1 vccd1 _15147_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_114_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout322 _14290_/A vssd1 vssd1 vccd1 vccd1 _14738_/A sky130_fd_sc_hd__clkbuf_2
Xfanout333 _12770_/B vssd1 vssd1 vccd1 vccd1 _17423_/A sky130_fd_sc_hd__buf_2
Xfanout344 _17538_/Q vssd1 vssd1 vccd1 vccd1 _13227_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_98_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout355 _12804_/B vssd1 vssd1 vccd1 vccd1 _17417_/A sky130_fd_sc_hd__clkbuf_4
Xfanout366 _13080_/A vssd1 vssd1 vccd1 vccd1 _14769_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_59_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout377 fanout380/X vssd1 vssd1 vccd1 vccd1 _17411_/A sky130_fd_sc_hd__buf_2
X_09817_ _09814_/X _09817_/B vssd1 vssd1 vccd1 vccd1 _09828_/B sky130_fd_sc_hd__and2b_1
XFILLER_101_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout388 _13903_/A vssd1 vssd1 vccd1 vccd1 _14176_/A sky130_fd_sc_hd__buf_2
XFILLER_100_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout399 _17531_/Q vssd1 vssd1 vccd1 vccd1 _16644_/C sky130_fd_sc_hd__buf_2
XFILLER_47_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09748_ _09892_/A _09892_/B _10299_/D _10421_/D vssd1 vssd1 vccd1 vccd1 _09751_/A
+ sky130_fd_sc_hd__and4_1
XTAP_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09679_ _09679_/A _09679_/B vssd1 vssd1 vccd1 vccd1 _12016_/A sky130_fd_sc_hd__nor2_1
XTAP_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11710_ _15997_/A _15997_/B _16105_/A _11709_/Y _11708_/B vssd1 vssd1 vccd1 vccd1
+ _16206_/A sky130_fd_sc_hd__a32o_1
XFILLER_54_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12690_ _12689_/A _12689_/B _12689_/C vssd1 vssd1 vccd1 vccd1 _12691_/B sky130_fd_sc_hd__o21a_1
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_979 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11641_ _11641_/A _11664_/A vssd1 vssd1 vccd1 vccd1 _11648_/A sky130_fd_sc_hd__xor2_1
XTAP_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14360_ _14641_/A _14641_/B _16859_/A _14360_/D vssd1 vssd1 vccd1 vccd1 _14440_/A
+ sky130_fd_sc_hd__and4_1
X_11572_ _11572_/A _11576_/B _11572_/C _11572_/D vssd1 vssd1 vccd1 vccd1 _11607_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_10_331 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13311_ _13317_/A vssd1 vssd1 vccd1 vccd1 _13431_/A sky130_fd_sc_hd__inv_2
X_10523_ _10437_/X _10521_/Y _10517_/A _10502_/X vssd1 vssd1 vccd1 vccd1 _10523_/Y
+ sky130_fd_sc_hd__o211ai_1
XFILLER_122_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput19 i_wb_addr[24] vssd1 vssd1 vccd1 vccd1 input19/X sky130_fd_sc_hd__clkbuf_1
X_14291_ _14291_/A _14372_/A vssd1 vssd1 vccd1 vccd1 _14294_/A sky130_fd_sc_hd__or2_1
XFILLER_109_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16030_ _16315_/C _16662_/D vssd1 vssd1 vccd1 vccd1 _16136_/C sky130_fd_sc_hd__nor2_1
X_13242_ _13243_/A _13243_/B vssd1 vssd1 vccd1 vccd1 _13244_/B sky130_fd_sc_hd__nand2_1
XFILLER_171_818 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10454_ _10454_/A _10454_/B vssd1 vssd1 vccd1 vccd1 _10456_/B sky130_fd_sc_hd__nand2_1
XFILLER_170_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_200 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13173_ _13174_/A _13174_/B vssd1 vssd1 vccd1 vccd1 _13314_/B sky130_fd_sc_hd__and2b_1
X_10385_ _10385_/A _10385_/B _10385_/C vssd1 vssd1 vccd1 vccd1 _10385_/Y sky130_fd_sc_hd__nand3_1
XFILLER_163_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12124_ _12121_/X _12122_/Y _11915_/A _11916_/Y vssd1 vssd1 vccd1 vccd1 _12151_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_2_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16932_ _16909_/A _16851_/A _16909_/B vssd1 vssd1 vccd1 vccd1 _16932_/X sky130_fd_sc_hd__a21bo_1
XFILLER_78_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12055_ _10657_/C _14956_/B _12046_/A vssd1 vssd1 vccd1 vccd1 _12055_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_96_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11006_ _11006_/A _11006_/B _11006_/C vssd1 vssd1 vccd1 vccd1 _11006_/X sky130_fd_sc_hd__and3_1
XFILLER_77_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16863_ _16863_/A _16863_/B vssd1 vssd1 vccd1 vccd1 _16863_/Y sky130_fd_sc_hd__nand2_1
XFILLER_65_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15814_ _15792_/X _15794_/X _15813_/X _16494_/B1 _15811_/A vssd1 vssd1 vccd1 vccd1
+ _15815_/A sky130_fd_sc_hd__a32o_1
X_16794_ _16794_/A _16794_/B vssd1 vssd1 vccd1 vccd1 _16795_/B sky130_fd_sc_hd__nand2_1
XFILLER_65_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15745_ _16745_/A _16021_/B vssd1 vssd1 vccd1 vccd1 _16681_/C sky130_fd_sc_hd__nand2_4
XTAP_3271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12957_ _13578_/A _13966_/C vssd1 vssd1 vccd1 vccd1 _12959_/B sky130_fd_sc_hd__nand2_1
XFILLER_80_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11908_ _11908_/A _11908_/B vssd1 vssd1 vccd1 vccd1 _11909_/B sky130_fd_sc_hd__nor2_1
X_15676_ _15676_/A vssd1 vssd1 vccd1 vccd1 _15772_/A sky130_fd_sc_hd__inv_2
XTAP_2570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12888_ _12723_/A _12725_/B _12723_/B vssd1 vssd1 vccd1 vccd1 _12895_/A sky130_fd_sc_hd__o21ba_1
XTAP_2581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17415_ _17415_/A _17425_/B vssd1 vssd1 vccd1 vccd1 _17415_/X sky130_fd_sc_hd__or2_1
XFILLER_60_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14627_ _14627_/A _14627_/B _14627_/C vssd1 vssd1 vccd1 vccd1 _14628_/B sky130_fd_sc_hd__or3_1
X_11839_ _12334_/B _12328_/B _11839_/S vssd1 vssd1 vccd1 vccd1 _11840_/B sky130_fd_sc_hd__mux2_1
XTAP_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17346_ _12258_/B _17356_/A2 _17345_/X _17406_/C1 vssd1 vssd1 vccd1 vccd1 _17502_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_158_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14558_ _14558_/A _14558_/B vssd1 vssd1 vccd1 vccd1 _14560_/A sky130_fd_sc_hd__nor2_1
XFILLER_174_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13509_ _13509_/A _13509_/B vssd1 vssd1 vccd1 vccd1 _13509_/Y sky130_fd_sc_hd__nor2_1
XFILLER_174_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17277_ _17569_/Q _17292_/B vssd1 vssd1 vccd1 vccd1 _17277_/X sky130_fd_sc_hd__and2_1
XFILLER_174_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14489_ _14489_/A _14489_/B vssd1 vssd1 vccd1 vccd1 _14490_/B sky130_fd_sc_hd__and2_1
XFILLER_146_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16228_ _16315_/C _16813_/B vssd1 vssd1 vccd1 vccd1 _16229_/B sky130_fd_sc_hd__nor2_1
XFILLER_155_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16159_ _16036_/A _16036_/B _16047_/X vssd1 vssd1 vccd1 vccd1 _16161_/B sky130_fd_sc_hd__a21oi_2
XFILLER_6_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08981_ _08981_/A vssd1 vssd1 vccd1 vccd1 _08983_/B sky130_fd_sc_hd__inv_2
XFILLER_142_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_835 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09602_ _09602_/A _09610_/A _09602_/C vssd1 vssd1 vccd1 vccd1 _09603_/B sky130_fd_sc_hd__or3_1
XFILLER_83_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09533_ _09487_/X _09530_/B _09531_/X _09532_/Y vssd1 vssd1 vccd1 vccd1 _09540_/A
+ sky130_fd_sc_hd__a211oi_1
XFILLER_36_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_935 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09464_ _09892_/A _09892_/B _10543_/B _10545_/D vssd1 vssd1 vccd1 vccd1 _09473_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_19_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09395_ _09395_/A _09395_/B _09395_/C vssd1 vssd1 vccd1 vccd1 _09395_/X sky130_fd_sc_hd__or3_1
XFILLER_52_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10170_ _10170_/A _10174_/A _10170_/C vssd1 vssd1 vccd1 vccd1 _10177_/B sky130_fd_sc_hd__or3_1
XFILLER_160_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout130 _17187_/Y vssd1 vssd1 vccd1 vccd1 _17225_/A2 sky130_fd_sc_hd__buf_2
Xfanout141 _15088_/B vssd1 vssd1 vccd1 vccd1 _16086_/A sky130_fd_sc_hd__clkbuf_4
Xfanout152 _14911_/X vssd1 vssd1 vccd1 vccd1 _15100_/A sky130_fd_sc_hd__buf_2
Xfanout163 _17308_/A2 vssd1 vssd1 vccd1 vccd1 _17322_/A2 sky130_fd_sc_hd__clkbuf_4
Xfanout174 _16883_/A vssd1 vssd1 vccd1 vccd1 _16938_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_47_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout185 _15854_/B vssd1 vssd1 vccd1 vccd1 _16812_/A sky130_fd_sc_hd__buf_4
XFILLER_75_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout196 _14926_/X vssd1 vssd1 vccd1 vccd1 _16582_/A sky130_fd_sc_hd__clkbuf_4
X_13860_ _13861_/A _13861_/B _13861_/C vssd1 vssd1 vccd1 vccd1 _13964_/A sky130_fd_sc_hd__a21o_1
XFILLER_47_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12811_ _12812_/B _12812_/A vssd1 vssd1 vccd1 vccd1 _12972_/B sky130_fd_sc_hd__and2b_1
XFILLER_34_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13791_ _14387_/A _14426_/D vssd1 vssd1 vccd1 vccd1 _13792_/B sky130_fd_sc_hd__nand2_1
XFILLER_90_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15530_ _15541_/A _16571_/B _15472_/A vssd1 vssd1 vccd1 vccd1 _15620_/A sky130_fd_sc_hd__or3b_1
X_12742_ _12902_/A _12743_/B _12743_/C vssd1 vssd1 vccd1 vccd1 _12744_/A sky130_fd_sc_hd__a21o_1
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12673_ _12673_/A _12673_/B vssd1 vssd1 vccd1 vccd1 _12675_/B sky130_fd_sc_hd__xnor2_1
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15461_ _15628_/A _15460_/X _14962_/B vssd1 vssd1 vccd1 vccd1 _15461_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_15_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17200_ _17434_/Q _17171_/X _17197_/X _17199_/X _17428_/B vssd1 vssd1 vccd1 vccd1
+ _17434_/D sky130_fd_sc_hd__o221a_1
X_11624_ _11624_/A _11624_/B vssd1 vssd1 vccd1 vccd1 _11624_/Y sky130_fd_sc_hd__nand2_1
XFILLER_8_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14412_ _14413_/A _14413_/B _14413_/C vssd1 vssd1 vccd1 vccd1 _14414_/A sky130_fd_sc_hd__o21a_1
XFILLER_129_804 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15392_ _15381_/A _17170_/B1 _15391_/Y vssd1 vssd1 vccd1 vccd1 _17550_/D sky130_fd_sc_hd__a21oi_1
XFILLER_156_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17131_ _17131_/A _17131_/B _17131_/C vssd1 vssd1 vccd1 vccd1 _17131_/X sky130_fd_sc_hd__and3_1
X_11555_ _11555_/A _11555_/B _11637_/A vssd1 vssd1 vccd1 vccd1 _11558_/B sky130_fd_sc_hd__nor3b_1
XFILLER_11_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14343_ _14344_/A _14344_/B _14344_/C vssd1 vssd1 vccd1 vccd1 _14413_/A sky130_fd_sc_hd__o21a_1
XFILLER_156_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10506_ _10963_/A _10963_/B _10736_/D _10875_/C vssd1 vssd1 vccd1 vccd1 _10509_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_7_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17062_ _17062_/A _17062_/B vssd1 vssd1 vccd1 vccd1 _17063_/B sky130_fd_sc_hd__xor2_1
XFILLER_7_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14274_ _14350_/B _14274_/B vssd1 vssd1 vccd1 vccd1 _14274_/X sky130_fd_sc_hd__or2_1
X_11486_ _11477_/A _11477_/C _11514_/A vssd1 vssd1 vccd1 vccd1 _11487_/B sky130_fd_sc_hd__a21oi_1
XFILLER_109_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13225_ _13068_/A _13070_/B _13068_/B vssd1 vssd1 vccd1 vccd1 _13232_/A sky130_fd_sc_hd__o21ba_1
X_16013_ _17143_/A1 _13624_/X _15808_/A _16012_/X vssd1 vssd1 vccd1 vccd1 _16017_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_109_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10437_ _10437_/A _10437_/B _10437_/C vssd1 vssd1 vccd1 vccd1 _10437_/X sky130_fd_sc_hd__and3_1
XFILLER_109_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13156_ _13641_/A _13156_/B _13632_/D _13522_/D vssd1 vssd1 vccd1 vccd1 _13157_/B
+ sky130_fd_sc_hd__and4_1
X_10368_ _10484_/B vssd1 vssd1 vccd1 vccd1 _10369_/B sky130_fd_sc_hd__inv_2
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12107_ _12275_/A _12275_/B _12275_/D _12258_/B vssd1 vssd1 vccd1 vccd1 _12108_/B
+ sky130_fd_sc_hd__and4_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13087_ _13087_/A _13220_/A vssd1 vssd1 vccd1 vccd1 _13088_/C sky130_fd_sc_hd__and2_1
XFILLER_111_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10299_ _10300_/A _10298_/Y _15805_/A _10299_/D vssd1 vssd1 vccd1 vccd1 _10418_/A
+ sky130_fd_sc_hd__and4bb_1
X_12038_ _12028_/X _12037_/Y _13833_/S vssd1 vssd1 vccd1 vccd1 _12038_/X sky130_fd_sc_hd__mux2_1
X_16915_ _16863_/A _16863_/B _16858_/Y vssd1 vssd1 vccd1 vccd1 _16916_/B sky130_fd_sc_hd__a21oi_1
XFILLER_111_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16846_ _16846_/A _16846_/B _16846_/C vssd1 vssd1 vccd1 vccd1 _16847_/B sky130_fd_sc_hd__or3_1
XFILLER_66_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16777_ _16777_/A _16777_/B _16777_/C vssd1 vssd1 vccd1 vccd1 _16778_/B sky130_fd_sc_hd__and3_1
XFILLER_81_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13989_ _14077_/A _13989_/B vssd1 vssd1 vccd1 vccd1 _13990_/B sky130_fd_sc_hd__nor2_1
XFILLER_80_326 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15728_ _15834_/A _15728_/B vssd1 vssd1 vccd1 vccd1 _15730_/B sky130_fd_sc_hd__nor2_1
XFILLER_61_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15659_ _16056_/A _16259_/B vssd1 vssd1 vccd1 vccd1 _15661_/B sky130_fd_sc_hd__nand2_1
XFILLER_21_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09180_ _09358_/A _09345_/B vssd1 vssd1 vccd1 vccd1 _09346_/A sky130_fd_sc_hd__and2_1
XFILLER_105_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17329_ input43/X _17359_/B _17359_/C vssd1 vssd1 vccd1 vccd1 _17329_/X sky130_fd_sc_hd__or3_1
XFILLER_30_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08964_ _09654_/C _17139_/A vssd1 vssd1 vccd1 vccd1 _08993_/C sky130_fd_sc_hd__nand2_1
XFILLER_102_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08895_ _08895_/A _08895_/B vssd1 vssd1 vccd1 vccd1 _08903_/A sky130_fd_sc_hd__xnor2_1
XFILLER_69_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_846 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_24 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09516_ _09517_/A _09515_/Y _09639_/C _10072_/B vssd1 vssd1 vccd1 vccd1 _09636_/A
+ sky130_fd_sc_hd__and4bb_1
XPHY_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09447_ _09447_/A _09583_/A vssd1 vssd1 vccd1 vccd1 _09449_/B sky130_fd_sc_hd__nor2_1
XPHY_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09378_ _09379_/A _09377_/Y _09639_/C _09937_/B vssd1 vssd1 vccd1 vccd1 _09513_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_71_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_34 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11340_ _11340_/A _11340_/B vssd1 vssd1 vccd1 vccd1 _11341_/C sky130_fd_sc_hd__xnor2_1
XFILLER_137_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11271_ _11313_/A _11313_/B vssd1 vssd1 vccd1 vccd1 _11274_/C sky130_fd_sc_hd__nand2_1
XFILLER_3_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13010_ _13268_/A _13010_/B vssd1 vssd1 vccd1 vccd1 _13138_/B sky130_fd_sc_hd__nand2b_1
X_10222_ _10559_/A _09937_/B _09953_/B _09952_/A vssd1 vssd1 vccd1 vccd1 _10226_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_140_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10153_ _10149_/A _10152_/X _10137_/X _10138_/Y vssd1 vssd1 vccd1 vccd1 _10155_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_160_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10084_ _10084_/A _10084_/B vssd1 vssd1 vccd1 vccd1 _10086_/B sky130_fd_sc_hd__nand2_1
X_14961_ _15460_/B _15458_/B _17369_/A vssd1 vssd1 vccd1 vccd1 _14961_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16700_ _16701_/A _16701_/B vssd1 vssd1 vccd1 vccd1 _16777_/B sky130_fd_sc_hd__or2_1
X_13912_ _13912_/A _13912_/B vssd1 vssd1 vccd1 vccd1 _13913_/B sky130_fd_sc_hd__nand2_1
XFILLER_75_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14892_ _16760_/A _15204_/B _16807_/A vssd1 vssd1 vccd1 vccd1 _15208_/C sky130_fd_sc_hd__or3_2
X_16631_ _16711_/A _16631_/B vssd1 vssd1 vccd1 vccd1 _16634_/A sky130_fd_sc_hd__or2_1
XFILLER_47_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13843_ _13948_/B _13844_/C _14008_/B _13948_/A vssd1 vssd1 vccd1 vccd1 _13845_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_74_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwb_buttons_leds_960 vssd1 vssd1 vccd1 vccd1 wb_buttons_leds_960/HI led_enb[2] sky130_fd_sc_hd__conb_1
XFILLER_74_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16562_ _16561_/X _16562_/B _16562_/C vssd1 vssd1 vccd1 vccd1 _16562_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_74_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10986_ _10987_/A _10987_/B vssd1 vssd1 vccd1 vccd1 _11162_/B sky130_fd_sc_hd__nand2_1
X_13774_ _13774_/A _13774_/B vssd1 vssd1 vccd1 vccd1 _13776_/A sky130_fd_sc_hd__nor2_1
XFILLER_16_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15513_ _15514_/A _15514_/B _15514_/C vssd1 vssd1 vccd1 vccd1 _15609_/A sky130_fd_sc_hd__a21oi_1
X_12725_ _12725_/A _12725_/B vssd1 vssd1 vccd1 vccd1 _12727_/B sky130_fd_sc_hd__xnor2_1
X_16493_ _16483_/X _16493_/B _16493_/C vssd1 vssd1 vccd1 vccd1 _16493_/X sky130_fd_sc_hd__and3b_1
XFILLER_70_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15444_ _15442_/Y _15443_/X _16911_/A vssd1 vssd1 vccd1 vccd1 _15444_/Y sky130_fd_sc_hd__o21ai_1
X_12656_ _12804_/B _13194_/D _13067_/D _12804_/A vssd1 vssd1 vccd1 vccd1 _12658_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_157_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11607_ _11607_/A _11607_/B _11607_/C vssd1 vssd1 vccd1 vccd1 _11613_/A sky130_fd_sc_hd__nand3_1
X_12587_ _12588_/A _12588_/B _12588_/C vssd1 vssd1 vccd1 vccd1 _12612_/A sky130_fd_sc_hd__a21oi_4
X_15375_ _15307_/B _15307_/C _15307_/A vssd1 vssd1 vccd1 vccd1 _15375_/X sky130_fd_sc_hd__o21ba_1
XFILLER_12_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17114_ _14828_/Y _16304_/A _17104_/X _17107_/X _17113_/X vssd1 vssd1 vccd1 vccd1
+ _17114_/X sky130_fd_sc_hd__o311a_1
X_14326_ _16723_/A _14450_/B _14326_/C vssd1 vssd1 vccd1 vccd1 _14393_/B sky130_fd_sc_hd__nand3_1
X_11538_ _11538_/A _11538_/B vssd1 vssd1 vccd1 vccd1 _11538_/X sky130_fd_sc_hd__or2_1
XFILLER_116_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17045_ _17046_/A _17046_/B _17046_/C vssd1 vssd1 vccd1 vccd1 _17088_/A sky130_fd_sc_hd__o21a_1
X_11469_ _11553_/B _11561_/D vssd1 vssd1 vccd1 vccd1 _11469_/X sky130_fd_sc_hd__and2_1
X_14257_ _14258_/A _14258_/B vssd1 vssd1 vccd1 vccd1 _14257_/Y sky130_fd_sc_hd__nand2_1
XFILLER_172_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13208_ _14769_/A _13450_/B _13208_/C _13208_/D vssd1 vssd1 vccd1 vccd1 _13339_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_171_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14188_ _14188_/A _14188_/B _14188_/C vssd1 vssd1 vccd1 vccd1 _14189_/B sky130_fd_sc_hd__and3_1
XFILLER_112_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13139_ _13268_/B _13140_/B vssd1 vssd1 vccd1 vccd1 _13139_/X sky130_fd_sc_hd__or2_1
XFILLER_98_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_334 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_676 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16829_ _16829_/A _16829_/B vssd1 vssd1 vccd1 vccd1 _16830_/B sky130_fd_sc_hd__xnor2_1
XFILLER_53_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09301_ _09302_/A _09300_/Y _09730_/C _12077_/C vssd1 vssd1 vccd1 vccd1 _09443_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_55_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09232_ _12804_/B _12129_/B _12127_/C _12804_/A vssd1 vssd1 vccd1 vccd1 _09234_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_22_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09163_ _09164_/A _09163_/B _09654_/C _09350_/B vssd1 vssd1 vccd1 vccd1 _09354_/A
+ sky130_fd_sc_hd__and4b_1
XFILLER_148_954 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09094_ _08973_/B _08971_/C _08993_/C vssd1 vssd1 vccd1 vccd1 _09095_/B sky130_fd_sc_hd__o21a_1
XFILLER_147_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09996_ _09996_/A _09996_/B vssd1 vssd1 vccd1 vccd1 _10003_/A sky130_fd_sc_hd__xnor2_1
XFILLER_48_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08947_ _09078_/A _08947_/B _12256_/C _12256_/D vssd1 vssd1 vccd1 vccd1 _08950_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_29_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08878_ _08883_/A _08883_/B vssd1 vssd1 vccd1 vccd1 _08889_/A sky130_fd_sc_hd__nor2_1
XFILLER_151_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_816 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_698 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_326 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10840_ _11122_/B _10933_/D _10970_/B _10933_/A vssd1 vssd1 vccd1 vccd1 _10841_/B
+ sky130_fd_sc_hd__a22oi_1
XFILLER_71_123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10771_ _10771_/A _10771_/B _10771_/C vssd1 vssd1 vccd1 vccd1 _10772_/B sky130_fd_sc_hd__or3_1
XFILLER_71_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12510_ _12339_/A _12341_/B _12339_/B vssd1 vssd1 vccd1 vccd1 _12511_/B sky130_fd_sc_hd__o21ba_1
XFILLER_44_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13490_ _13607_/A _13490_/B _13490_/C _13490_/D vssd1 vssd1 vccd1 vccd1 _13492_/A
+ sky130_fd_sc_hd__nor4_1
XFILLER_12_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12441_ _12442_/A _12592_/C _12442_/C vssd1 vssd1 vccd1 vccd1 _12443_/A sky130_fd_sc_hd__a21oi_1
XFILLER_40_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12372_ _12373_/A _12373_/B vssd1 vssd1 vccd1 vccd1 _12372_/X sky130_fd_sc_hd__or2_1
X_15160_ _15161_/A _15161_/B vssd1 vssd1 vccd1 vccd1 _15162_/A sky130_fd_sc_hd__or2_1
XFILLER_138_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11323_ _11553_/A _11561_/C _11563_/D _11427_/A vssd1 vssd1 vccd1 vccd1 _11324_/D
+ sky130_fd_sc_hd__a22o_1
X_14111_ _14197_/B _14111_/B vssd1 vssd1 vccd1 vccd1 _14113_/C sky130_fd_sc_hd__nand2_1
XFILLER_165_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15091_ _15091_/A _15091_/B vssd1 vssd1 vccd1 vccd1 _15170_/B sky130_fd_sc_hd__or2_1
XFILLER_153_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11254_ _11139_/A _11139_/B _11139_/C vssd1 vssd1 vccd1 vccd1 _11255_/C sky130_fd_sc_hd__a21oi_1
XFILLER_125_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14042_ _14043_/A _14043_/B vssd1 vssd1 vccd1 vccd1 _14042_/Y sky130_fd_sc_hd__nand2_1
XFILLER_4_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10205_ _10469_/B _10205_/B vssd1 vssd1 vccd1 vccd1 _10331_/B sky130_fd_sc_hd__nor2_1
X_11185_ _11182_/Y _11183_/X _11039_/Y _11041_/Y vssd1 vssd1 vccd1 vccd1 _11186_/D
+ sky130_fd_sc_hd__o211ai_1
XFILLER_79_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10136_ _10136_/A _10136_/B vssd1 vssd1 vccd1 vccd1 _10138_/C sky130_fd_sc_hd__xnor2_1
XFILLER_79_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15993_ _15991_/X _15994_/B vssd1 vssd1 vccd1 vccd1 _15993_/X sky130_fd_sc_hd__and2b_1
XFILLER_48_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10067_ _10321_/B _10067_/B _10067_/C vssd1 vssd1 vccd1 vccd1 _10200_/A sky130_fd_sc_hd__and3_1
X_14944_ _14944_/A _14944_/B _14944_/C vssd1 vssd1 vccd1 vccd1 _14944_/Y sky130_fd_sc_hd__nor3_1
XFILLER_78_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14875_ _14888_/C _14876_/C _14876_/D vssd1 vssd1 vccd1 vccd1 _14875_/X sky130_fd_sc_hd__or3_1
XFILLER_78_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16614_ _16614_/A _16614_/B vssd1 vssd1 vccd1 vccd1 _16616_/C sky130_fd_sc_hd__xnor2_1
XFILLER_35_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13826_ _13824_/A _13824_/B _13827_/A vssd1 vssd1 vccd1 vccd1 _13826_/Y sky130_fd_sc_hd__a21oi_1
X_17594_ fanout933/X _17594_/D vssd1 vssd1 vccd1 vccd1 _17594_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16545_ _16545_/A _16545_/B vssd1 vssd1 vccd1 vccd1 _16547_/B sky130_fd_sc_hd__xnor2_1
XFILLER_16_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13757_ _13756_/B _13757_/B vssd1 vssd1 vccd1 vccd1 _13758_/B sky130_fd_sc_hd__and2b_1
X_10969_ _10969_/A _10969_/B vssd1 vssd1 vccd1 vccd1 _10976_/A sky130_fd_sc_hd__xnor2_1
X_12708_ _12040_/Y _12042_/Y _12397_/B _12061_/Y _12383_/S _16011_/B vssd1 vssd1 vccd1
+ vccd1 _12709_/B sky130_fd_sc_hd__mux4_1
XFILLER_149_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16476_ _11200_/Y _16389_/C _11229_/Y vssd1 vssd1 vccd1 vccd1 _16478_/A sky130_fd_sc_hd__a21oi_1
X_13688_ _13688_/A _13688_/B vssd1 vssd1 vccd1 vccd1 _13707_/A sky130_fd_sc_hd__xor2_1
XFILLER_15_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15427_ _15340_/X _15345_/B _15342_/Y vssd1 vssd1 vccd1 vccd1 _15429_/B sky130_fd_sc_hd__o21ai_1
X_12639_ _12640_/A _12792_/A _12640_/C vssd1 vssd1 vccd1 vccd1 _12641_/A sky130_fd_sc_hd__o21a_1
XFILLER_79_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15358_ _15358_/A _15358_/B vssd1 vssd1 vccd1 vccd1 _15359_/B sky130_fd_sc_hd__xnor2_1
XFILLER_172_721 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14309_ _14309_/A _14309_/B vssd1 vssd1 vccd1 vccd1 _14312_/A sky130_fd_sc_hd__xor2_1
XFILLER_145_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15289_ _16086_/A _16317_/B vssd1 vssd1 vccd1 vccd1 _15291_/B sky130_fd_sc_hd__nand2_1
XFILLER_116_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17028_ _17028_/A _17028_/B vssd1 vssd1 vccd1 vccd1 _17029_/C sky130_fd_sc_hd__nor2_1
XFILLER_104_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout707 _10431_/B vssd1 vssd1 vccd1 vccd1 _10311_/D sky130_fd_sc_hd__buf_2
X_09850_ _09863_/B _09863_/C _09863_/A vssd1 vssd1 vccd1 vccd1 _09865_/A sky130_fd_sc_hd__a21o_1
XFILLER_112_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout718 _13966_/C vssd1 vssd1 vccd1 vccd1 _13334_/C sky130_fd_sc_hd__buf_4
XFILLER_112_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_854 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout729 _12077_/D vssd1 vssd1 vccd1 vccd1 _09446_/D sky130_fd_sc_hd__clkbuf_4
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08801_ _08801_/A _08801_/B _08801_/C vssd1 vssd1 vccd1 vccd1 _08801_/Y sky130_fd_sc_hd__nand3_4
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09781_ _15254_/S _10180_/B _14949_/A vssd1 vssd1 vccd1 vccd1 _09781_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_86_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08732_ _17609_/Q _17610_/Q vssd1 vssd1 vccd1 vccd1 _08732_/X sky130_fd_sc_hd__and2_1
XFILLER_85_248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_679 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09215_ _17411_/A _09555_/D _12338_/D _17413_/A vssd1 vssd1 vccd1 vccd1 _09219_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_6_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09146_ _09147_/B _09231_/B vssd1 vssd1 vccd1 vccd1 _09148_/B sky130_fd_sc_hd__nor2_1
XFILLER_135_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09077_ _09077_/A _09077_/B vssd1 vssd1 vccd1 vccd1 _09091_/A sky130_fd_sc_hd__xnor2_1
XFILLER_107_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_832 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09979_ _09979_/A _10109_/B _09979_/C _10111_/D vssd1 vssd1 vccd1 vccd1 _09982_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_58_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12990_ _12987_/X _12988_/Y _12819_/X _12824_/A vssd1 vssd1 vccd1 vccd1 _12993_/B
+ sky130_fd_sc_hd__o211a_1
XTAP_3612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11941_ _11941_/A _11941_/B vssd1 vssd1 vccd1 vccd1 _11941_/Y sky130_fd_sc_hd__nor2_1
XTAP_2900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14660_ _14661_/A _14660_/B vssd1 vssd1 vccd1 vccd1 _14662_/B sky130_fd_sc_hd__nor2_1
XTAP_2944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11872_ _11872_/A vssd1 vssd1 vccd1 vccd1 _11874_/B sky130_fd_sc_hd__inv_2
XTAP_2955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_98 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13611_ _13718_/B _13609_/X _13495_/A _13497_/X vssd1 vssd1 vccd1 vccd1 _13612_/B
+ sky130_fd_sc_hd__a211oi_1
X_10823_ _10823_/A _10823_/B _10829_/B vssd1 vssd1 vccd1 vccd1 _11072_/B sky130_fd_sc_hd__or3_1
XTAP_2988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14591_ _14735_/A1 _12037_/A _13625_/Y _12853_/X vssd1 vssd1 vccd1 vccd1 _14591_/X
+ sky130_fd_sc_hd__a31o_1
XTAP_2999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16330_ _16239_/A _16239_/B _16231_/Y vssd1 vssd1 vccd1 vccd1 _16331_/B sky130_fd_sc_hd__a21bo_1
XFILLER_125_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13542_ _13542_/A vssd1 vssd1 vccd1 vccd1 _13543_/B sky130_fd_sc_hd__inv_2
XFILLER_71_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10754_ _10753_/A _10993_/D _10543_/C vssd1 vssd1 vccd1 vccd1 _10754_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_9_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_1046 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16261_ _16358_/A _16261_/B vssd1 vssd1 vccd1 vccd1 _16262_/C sky130_fd_sc_hd__or2_1
X_13473_ _13473_/A _13473_/B vssd1 vssd1 vccd1 vccd1 _13476_/A sky130_fd_sc_hd__xnor2_1
XFILLER_9_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10685_ _10685_/A _10685_/B _10685_/C vssd1 vssd1 vccd1 vccd1 _10688_/A sky130_fd_sc_hd__nand3_1
X_15212_ _15493_/A _16410_/A vssd1 vssd1 vccd1 vccd1 _15213_/C sky130_fd_sc_hd__nor2_1
X_12424_ _13035_/A _12734_/B _12877_/C _14063_/C vssd1 vssd1 vccd1 vccd1 _12425_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_173_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16192_ _16192_/A _16192_/B vssd1 vssd1 vccd1 vccd1 _16195_/A sky130_fd_sc_hd__xnor2_1
XFILLER_127_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_272 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15143_ _15147_/D _15270_/B _15143_/C vssd1 vssd1 vccd1 vccd1 _15143_/X sky130_fd_sc_hd__or3_1
X_12355_ _12355_/A _12355_/B vssd1 vssd1 vccd1 vccd1 _12357_/B sky130_fd_sc_hd__xnor2_1
XFILLER_5_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11306_ _11306_/A _11306_/B vssd1 vssd1 vccd1 vccd1 _11364_/B sky130_fd_sc_hd__nor2_1
XFILLER_99_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15074_ _15475_/A _15074_/B vssd1 vssd1 vccd1 vccd1 _15913_/A sky130_fd_sc_hd__nand2_2
XFILLER_126_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12286_ _12286_/A _12286_/B _12286_/C vssd1 vssd1 vccd1 vccd1 _12286_/Y sky130_fd_sc_hd__nand3_1
XFILLER_84_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11237_ _11237_/A _11237_/B vssd1 vssd1 vccd1 vccd1 _11295_/A sky130_fd_sc_hd__nand2_1
X_14025_ _14025_/A _14025_/B vssd1 vssd1 vccd1 vccd1 _14025_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_84_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11168_ _11168_/A _11168_/B _11167_/X vssd1 vssd1 vccd1 vccd1 _11168_/Y sky130_fd_sc_hd__nor3b_2
XFILLER_122_684 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10119_ _10119_/A _10119_/B vssd1 vssd1 vccd1 vccd1 _10232_/B sky130_fd_sc_hd__xnor2_1
X_11099_ _11099_/A _11099_/B _11101_/B vssd1 vssd1 vccd1 vccd1 _11104_/B sky130_fd_sc_hd__or3_1
X_15976_ _15976_/A _15976_/B vssd1 vssd1 vccd1 vccd1 _15984_/A sky130_fd_sc_hd__xnor2_1
XFILLER_64_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14927_ _15715_/A _14919_/X _14923_/Y _16582_/A vssd1 vssd1 vccd1 vccd1 _14927_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_76_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_134 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14858_ _16114_/A _16014_/A _16014_/B vssd1 vssd1 vccd1 vccd1 _16115_/B sky130_fd_sc_hd__and3_1
XFILLER_91_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13809_ _13809_/A _13809_/B vssd1 vssd1 vccd1 vccd1 _13810_/B sky130_fd_sc_hd__and2_1
XFILLER_63_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17577_ fanout939/X _17577_/D vssd1 vssd1 vccd1 vccd1 _17577_/Q sky130_fd_sc_hd__dfxtp_1
X_14789_ _14789_/A _14906_/B vssd1 vssd1 vccd1 vccd1 _15244_/B sky130_fd_sc_hd__nor2_1
XFILLER_90_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16528_ _16630_/A _16528_/B vssd1 vssd1 vccd1 vccd1 _16547_/A sky130_fd_sc_hd__and2_1
XFILLER_50_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16459_ _16459_/A _16459_/B vssd1 vssd1 vccd1 vccd1 _16460_/B sky130_fd_sc_hd__or2_1
X_09000_ _09327_/C _17139_/A vssd1 vssd1 vccd1 vccd1 _09001_/B sky130_fd_sc_hd__nand2_1
XFILLER_145_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09902_ _09902_/A _09902_/B vssd1 vssd1 vccd1 vccd1 _10034_/C sky130_fd_sc_hd__xnor2_1
XFILLER_99_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout504 _17519_/Q vssd1 vssd1 vccd1 vccd1 _15472_/A sky130_fd_sc_hd__buf_4
Xfanout515 _09892_/B vssd1 vssd1 vccd1 vccd1 _08947_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout526 _17516_/Q vssd1 vssd1 vccd1 vccd1 _15305_/C sky130_fd_sc_hd__clkbuf_4
Xfanout537 _09899_/A vssd1 vssd1 vccd1 vccd1 _12471_/A sky130_fd_sc_hd__clkbuf_4
X_09833_ _09720_/A _09719_/C _09719_/B vssd1 vssd1 vccd1 vccd1 _09866_/B sky130_fd_sc_hd__a21o_1
XFILLER_113_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout548 _14925_/A vssd1 vssd1 vccd1 vccd1 _14421_/S sky130_fd_sc_hd__clkbuf_4
Xfanout559 _09899_/B vssd1 vssd1 vccd1 vccd1 _10851_/B sky130_fd_sc_hd__buf_2
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09764_ _09788_/A _09764_/B vssd1 vssd1 vccd1 vccd1 _09765_/C sky130_fd_sc_hd__and2_1
XFILLER_86_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09695_ _09695_/A _09842_/A vssd1 vssd1 vccd1 vccd1 _09703_/B sky130_fd_sc_hd__nor2_1
XFILLER_54_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10470_ _10470_/A _10470_/B vssd1 vssd1 vccd1 vccd1 _10582_/A sky130_fd_sc_hd__or2_1
XFILLER_148_570 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09129_ _09502_/A _09128_/B _09126_/Y _09139_/A vssd1 vssd1 vccd1 vccd1 _09130_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_135_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12140_ _12141_/A _12141_/B vssd1 vssd1 vccd1 vccd1 _12305_/B sky130_fd_sc_hd__nand2_1
XFILLER_2_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_798 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12071_ _12070_/A _13080_/D _12070_/C _12070_/D vssd1 vssd1 vccd1 vccd1 _12072_/B
+ sky130_fd_sc_hd__a22oi_1
XFILLER_132_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11022_ _11022_/A _11022_/B vssd1 vssd1 vccd1 vccd1 _11024_/C sky130_fd_sc_hd__xor2_1
XFILLER_1_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15830_ _16315_/C _15932_/A _16827_/A _16514_/A vssd1 vssd1 vccd1 vccd1 _15831_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_92_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15761_ _15762_/A _15762_/B vssd1 vssd1 vccd1 vccd1 _15868_/A sky130_fd_sc_hd__and2_1
X_12973_ _12974_/A _12974_/B vssd1 vssd1 vccd1 vccd1 _13112_/A sky130_fd_sc_hd__or2_1
XTAP_3431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17500_ fanout946/X _17500_/D vssd1 vssd1 vccd1 vccd1 _17500_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14712_ _14744_/A _14712_/B vssd1 vssd1 vccd1 vccd1 _14713_/C sky130_fd_sc_hd__xnor2_1
XTAP_3464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11924_ _11924_/A _11924_/B vssd1 vssd1 vccd1 vccd1 _11925_/B sky130_fd_sc_hd__and2_1
XFILLER_45_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15692_ _15591_/A _15600_/Y _15779_/B _15691_/Y vssd1 vssd1 vccd1 vccd1 _15786_/A
+ sky130_fd_sc_hd__o211a_1
XTAP_2741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_999 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17431_ input47/X _17608_/Q _17433_/S vssd1 vssd1 vccd1 vccd1 _17608_/D sky130_fd_sc_hd__mux2_1
XTAP_2763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14643_ _14676_/A _14708_/D _14644_/C vssd1 vssd1 vccd1 vccd1 _14645_/A sky130_fd_sc_hd__a21oi_1
XTAP_2774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11855_ _16012_/S _11854_/X _15457_/A vssd1 vssd1 vccd1 vccd1 _11855_/X sky130_fd_sc_hd__o21a_1
XFILLER_72_284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10806_ _11095_/B _11115_/C _17469_/D _11095_/A vssd1 vssd1 vccd1 vccd1 _10807_/B
+ sky130_fd_sc_hd__a22oi_1
X_17362_ _17362_/A _17362_/B _17362_/C _17362_/D vssd1 vssd1 vccd1 vccd1 _17371_/B
+ sky130_fd_sc_hd__or4_4
XFILLER_82_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14574_ _14574_/A vssd1 vssd1 vccd1 vccd1 _14575_/B sky130_fd_sc_hd__inv_2
XFILLER_82_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11786_ _12016_/A _09826_/A _14837_/A _16922_/A vssd1 vssd1 vccd1 vccd1 _11786_/Y
+ sky130_fd_sc_hd__o31ai_1
X_16313_ _16313_/A vssd1 vssd1 vccd1 vccd1 _17560_/D sky130_fd_sc_hd__clkinv_2
X_13525_ _13524_/C _13637_/A _13523_/Y vssd1 vssd1 vccd1 vccd1 _13527_/B sky130_fd_sc_hd__a21bo_1
X_10737_ _11115_/B _10970_/B _10971_/B _11115_/A vssd1 vssd1 vccd1 vccd1 _10737_/Y
+ sky130_fd_sc_hd__a22oi_1
X_17293_ _17465_/Q _17293_/A2 _17291_/X _17292_/X _17293_/C1 vssd1 vssd1 vccd1 vccd1
+ _17465_/D sky130_fd_sc_hd__o221a_1
XFILLER_174_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16244_ _16814_/A _16827_/A vssd1 vssd1 vccd1 vccd1 _16245_/B sky130_fd_sc_hd__nor2_1
X_13456_ _13455_/A _13455_/B _13455_/C vssd1 vssd1 vccd1 vccd1 _13576_/A sky130_fd_sc_hd__o21ai_1
X_10668_ _10667_/A _10667_/Y _10556_/B _10587_/Y vssd1 vssd1 vccd1 vccd1 _10678_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_173_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12407_ _12871_/A _13208_/C _12408_/C vssd1 vssd1 vccd1 vccd1 _12409_/A sky130_fd_sc_hd__a21oi_1
X_16175_ _16175_/A _16175_/B vssd1 vssd1 vccd1 vccd1 _16177_/B sky130_fd_sc_hd__xor2_1
XFILLER_126_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10599_ _10599_/A _10599_/B vssd1 vssd1 vccd1 vccd1 _10711_/A sky130_fd_sc_hd__xor2_2
XFILLER_12_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13387_ _13508_/B _13388_/B vssd1 vssd1 vccd1 vccd1 _13387_/Y sky130_fd_sc_hd__nand2_1
XFILLER_115_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput107 _17464_/Q vssd1 vssd1 vccd1 vccd1 o_wb_data[30] sky130_fd_sc_hd__clkbuf_1
XFILLER_126_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15126_ _15126_/A _15126_/B vssd1 vssd1 vccd1 vccd1 _15126_/Y sky130_fd_sc_hd__nand2_1
XFILLER_115_927 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12338_ _17419_/A _17417_/A _12338_/C _12338_/D vssd1 vssd1 vccd1 vccd1 _12339_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_5_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15057_ _15056_/A _14913_/Y _15056_/Y _15097_/A vssd1 vssd1 vccd1 vccd1 _15057_/X
+ sky130_fd_sc_hd__a211o_1
X_12269_ _12592_/B _12439_/D _12447_/B _12592_/A vssd1 vssd1 vccd1 vccd1 _12271_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_96_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14008_ _14254_/A _14008_/B _14008_/C vssd1 vssd1 vccd1 vccd1 _14115_/B sky130_fd_sc_hd__nand3_1
XFILLER_95_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_354 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15959_ _16355_/A _16061_/B vssd1 vssd1 vccd1 vccd1 _15960_/B sky130_fd_sc_hd__nand2_1
XFILLER_36_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09480_ _09480_/A _09480_/B _09480_/C vssd1 vssd1 vccd1 vccd1 _09480_/X sky130_fd_sc_hd__and3_1
XFILLER_102_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_356 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_919 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout301 _17369_/A vssd1 vssd1 vccd1 vccd1 _13840_/S sky130_fd_sc_hd__clkbuf_2
Xfanout312 _15071_/A vssd1 vssd1 vccd1 vccd1 _15147_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_59_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout323 _14832_/A vssd1 vssd1 vccd1 vccd1 _14290_/A sky130_fd_sc_hd__buf_2
XFILLER_132_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout334 _08988_/B vssd1 vssd1 vccd1 vccd1 _12770_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_98_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout345 _14765_/A vssd1 vssd1 vccd1 vccd1 _14680_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_86_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout356 _09172_/A vssd1 vssd1 vccd1 vccd1 _12804_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_59_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout367 _17535_/Q vssd1 vssd1 vccd1 vccd1 _13080_/A sky130_fd_sc_hd__clkbuf_2
X_09816_ _09668_/Y _09683_/X _09772_/X _09813_/X vssd1 vssd1 vccd1 vccd1 _09817_/B
+ sky130_fd_sc_hd__a211o_1
Xfanout378 _14770_/A vssd1 vssd1 vccd1 vccd1 _09514_/B sky130_fd_sc_hd__buf_2
XFILLER_101_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout389 _16723_/A vssd1 vssd1 vccd1 vccd1 _13903_/A sky130_fd_sc_hd__buf_2
XFILLER_86_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09747_ _09747_/A _09747_/B vssd1 vssd1 vccd1 vccd1 _09762_/A sky130_fd_sc_hd__nand2_1
XFILLER_28_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_56 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09678_ _09678_/A _09678_/B _09681_/A vssd1 vssd1 vccd1 vccd1 _09679_/B sky130_fd_sc_hd__nor3_1
XTAP_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11640_ _11663_/A _11663_/B vssd1 vssd1 vccd1 vccd1 _11664_/A sky130_fd_sc_hd__nor2_1
XTAP_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11571_ _15305_/C _17467_/D _17466_/D _15373_/C vssd1 vssd1 vccd1 vccd1 _11572_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_22_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13310_ _13312_/A _13312_/B _13312_/C vssd1 vssd1 vccd1 vccd1 _13317_/A sky130_fd_sc_hd__o21ai_1
XFILLER_168_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10522_ _10502_/X _10517_/A _10521_/Y _10437_/X vssd1 vssd1 vccd1 vccd1 _10566_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_10_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14290_ _14290_/A _14708_/B _14360_/D _16722_/A vssd1 vssd1 vccd1 vccd1 _14372_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_109_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13241_ _13241_/A _13241_/B vssd1 vssd1 vccd1 vccd1 _13243_/B sky130_fd_sc_hd__xnor2_1
X_10453_ _10453_/A _10453_/B _10453_/C vssd1 vssd1 vccd1 vccd1 _10454_/B sky130_fd_sc_hd__nand3_1
XFILLER_108_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10384_ _10385_/A _10385_/B _10385_/C vssd1 vssd1 vccd1 vccd1 _10384_/X sky130_fd_sc_hd__and3_1
X_13172_ _13172_/A _13172_/B vssd1 vssd1 vccd1 vccd1 _13174_/B sky130_fd_sc_hd__xnor2_1
XFILLER_123_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12123_ _11915_/A _11916_/Y _12121_/X _12122_/Y vssd1 vssd1 vccd1 vccd1 _12316_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_97_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16931_ _16931_/A _16931_/B _16910_/B vssd1 vssd1 vccd1 vccd1 _16931_/X sky130_fd_sc_hd__or3b_1
XFILLER_123_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12054_ _12054_/A _12054_/B vssd1 vssd1 vccd1 vccd1 _14956_/B sky130_fd_sc_hd__and2_1
XFILLER_2_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11005_ _11005_/A _11005_/B vssd1 vssd1 vccd1 vccd1 _11009_/A sky130_fd_sc_hd__nand2_1
XFILLER_78_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16862_ _16863_/A _16863_/B vssd1 vssd1 vccd1 vccd1 _16862_/X sky130_fd_sc_hd__or2_1
XFILLER_93_803 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout890 _10446_/B vssd1 vssd1 vccd1 vccd1 _09362_/D sky130_fd_sc_hd__buf_2
XFILLER_93_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15813_ _16007_/A _15802_/Y _15812_/X _15800_/Y vssd1 vssd1 vccd1 vccd1 _15813_/X
+ sky130_fd_sc_hd__o211a_1
X_16793_ _17156_/B _16793_/B vssd1 vssd1 vccd1 vccd1 _16793_/X sky130_fd_sc_hd__or2_1
XFILLER_18_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15744_ _16745_/A _16021_/B vssd1 vssd1 vccd1 vccd1 _16165_/B sky130_fd_sc_hd__and2_4
XFILLER_19_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12956_ _12956_/A _12956_/B vssd1 vssd1 vccd1 vccd1 _12959_/A sky130_fd_sc_hd__nand2_1
XTAP_3261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11907_ _11908_/A _11908_/B vssd1 vssd1 vccd1 vccd1 _11909_/A sky130_fd_sc_hd__and2_1
X_15675_ _15675_/A _15675_/B vssd1 vssd1 vccd1 vccd1 _15676_/A sky130_fd_sc_hd__nor2_1
XTAP_2560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12887_ _12735_/A _12737_/B _12735_/B vssd1 vssd1 vccd1 vccd1 _12897_/A sky130_fd_sc_hd__o21ba_1
XFILLER_33_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17414_ input53/X _17422_/A2 _17413_/X _17426_/C1 vssd1 vssd1 vccd1 vccd1 _17535_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_2582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14626_ _14627_/A _14627_/B _14627_/C vssd1 vssd1 vccd1 vccd1 _14638_/A sky130_fd_sc_hd__o21ai_1
X_11838_ _11835_/Y _11837_/Y _12212_/S vssd1 vssd1 vccd1 vccd1 _11838_/X sky130_fd_sc_hd__mux2_1
XFILLER_60_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17345_ input52/X _17353_/B _17353_/C vssd1 vssd1 vccd1 vccd1 _17345_/X sky130_fd_sc_hd__or3_1
XTAP_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14557_ _14557_/A _14557_/B _14557_/C vssd1 vssd1 vccd1 vccd1 _14558_/B sky130_fd_sc_hd__nor3_1
XFILLER_159_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11769_ _11768_/A _16866_/A _16866_/B _11767_/X vssd1 vssd1 vccd1 vccd1 _16972_/B
+ sky130_fd_sc_hd__o31ai_4
XFILLER_158_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13508_ _13271_/A _13508_/B vssd1 vssd1 vccd1 vccd1 _13511_/B sky130_fd_sc_hd__and2b_1
X_17276_ _17601_/Q _17282_/A2 _17282_/B1 vssd1 vssd1 vccd1 vccd1 _17276_/X sky130_fd_sc_hd__a21o_1
XFILLER_146_326 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14488_ _14489_/A _14489_/B vssd1 vssd1 vccd1 vccd1 _14557_/B sky130_fd_sc_hd__nor2_1
XFILLER_158_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16227_ _16227_/A _16227_/B vssd1 vssd1 vccd1 vccd1 _16229_/A sky130_fd_sc_hd__nor2_1
XFILLER_9_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13439_ _13586_/B _13439_/B vssd1 vssd1 vccd1 vccd1 _13442_/B sky130_fd_sc_hd__nor2_1
XFILLER_61_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_307 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16158_ _16158_/A _16158_/B vssd1 vssd1 vccd1 vccd1 _16161_/A sky130_fd_sc_hd__xnor2_1
XFILLER_142_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15109_ _11472_/B _14791_/X _14797_/X _15108_/Y vssd1 vssd1 vccd1 vccd1 _15109_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_5_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16089_ _16089_/A _16089_/B vssd1 vssd1 vccd1 vccd1 _16092_/A sky130_fd_sc_hd__xnor2_2
X_08980_ _09238_/B _08980_/B vssd1 vssd1 vccd1 vccd1 _08981_/A sky130_fd_sc_hd__or2_1
XFILLER_87_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_866 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09601_ _09480_/X _09599_/Y _09597_/B _09580_/X vssd1 vssd1 vccd1 vccd1 _09601_/Y
+ sky130_fd_sc_hd__o211ai_1
XFILLER_111_996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09532_ _09393_/X _09398_/Y _09485_/X _09530_/X vssd1 vssd1 vccd1 vccd1 _09532_/Y
+ sky130_fd_sc_hd__a211oi_1
XFILLER_37_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09463_ _09463_/A _09463_/B vssd1 vssd1 vccd1 vccd1 _09478_/A sky130_fd_sc_hd__nand2_1
XFILLER_52_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09394_ _09395_/B _09395_/C _09395_/A vssd1 vssd1 vccd1 vccd1 _12005_/A sky130_fd_sc_hd__o21ai_1
XFILLER_22_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout131 _16760_/B vssd1 vssd1 vccd1 vccd1 _16152_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_59_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout142 _15020_/X vssd1 vssd1 vccd1 vccd1 _16226_/B sky130_fd_sc_hd__clkbuf_4
Xfanout153 _15475_/A vssd1 vssd1 vccd1 vccd1 _15726_/A sky130_fd_sc_hd__buf_2
XFILLER_102_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout164 _17360_/A2 vssd1 vssd1 vccd1 vccd1 _17356_/A2 sky130_fd_sc_hd__buf_2
XFILLER_47_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout175 _15575_/Y vssd1 vssd1 vccd1 vccd1 _16065_/B sky130_fd_sc_hd__buf_4
XFILLER_47_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout186 _16168_/A vssd1 vssd1 vccd1 vccd1 _16619_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_19_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout197 _13841_/A vssd1 vssd1 vccd1 vccd1 _14210_/B sky130_fd_sc_hd__buf_2
X_12810_ _12658_/A _12660_/B _12658_/B vssd1 vssd1 vccd1 vccd1 _12812_/B sky130_fd_sc_hd__o21ba_1
XFILLER_74_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13790_ _13790_/A _13790_/B vssd1 vssd1 vccd1 vccd1 _13792_/A sky130_fd_sc_hd__nor2_1
XFILLER_28_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12741_ _12741_/A _12741_/B vssd1 vssd1 vccd1 vccd1 _12743_/C sky130_fd_sc_hd__xnor2_1
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15460_ _15715_/A _15460_/B vssd1 vssd1 vccd1 vccd1 _15460_/X sky130_fd_sc_hd__or2_1
X_12672_ _12673_/A _12673_/B vssd1 vssd1 vccd1 vccd1 _12672_/X sky130_fd_sc_hd__or2_1
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14411_ _14473_/B _14411_/B vssd1 vssd1 vccd1 vccd1 _14413_/C sky130_fd_sc_hd__and2_1
X_11623_ _11583_/B _11587_/X _11617_/B _11616_/Y vssd1 vssd1 vccd1 vccd1 _11624_/B
+ sky130_fd_sc_hd__a211o_1
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_440 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15391_ _17131_/A _15369_/Y _15390_/Y vssd1 vssd1 vccd1 vccd1 _15391_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_23_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17130_ _17130_/A _17130_/B vssd1 vssd1 vccd1 vccd1 _17131_/C sky130_fd_sc_hd__or2_1
XFILLER_129_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14342_ _14342_/A _14342_/B vssd1 vssd1 vccd1 vccd1 _14344_/C sky130_fd_sc_hd__and2_1
X_11554_ _15116_/A _15274_/A _11506_/X _11507_/Y vssd1 vssd1 vccd1 vccd1 _11555_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_11_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17061_ _17060_/A _17060_/B _17062_/A vssd1 vssd1 vccd1 vccd1 _17096_/B sky130_fd_sc_hd__o21a_1
X_10505_ _10505_/A _10505_/B vssd1 vssd1 vccd1 vccd1 _10511_/A sky130_fd_sc_hd__nor2_1
XFILLER_6_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14273_ _14273_/A _14273_/B _14273_/C vssd1 vssd1 vccd1 vccd1 _14274_/B sky130_fd_sc_hd__and3_1
X_11485_ _11534_/A _11485_/B vssd1 vssd1 vccd1 vccd1 _11485_/X sky130_fd_sc_hd__and2_1
XFILLER_155_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16012_ _16010_/X _16011_/X _16012_/S vssd1 vssd1 vccd1 vccd1 _16012_/X sky130_fd_sc_hd__mux2_1
X_13224_ _13224_/A _13224_/B vssd1 vssd1 vccd1 vccd1 _13243_/A sky130_fd_sc_hd__and2_1
XFILLER_6_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10436_ _10436_/A _10436_/B vssd1 vssd1 vccd1 vccd1 _10437_/C sky130_fd_sc_hd__xnor2_1
X_13155_ _13156_/B _13632_/D _13522_/D _13641_/A vssd1 vssd1 vccd1 vccd1 _13157_/A
+ sky130_fd_sc_hd__a22oi_1
X_10367_ _10370_/C _10367_/B vssd1 vssd1 vccd1 vccd1 _10484_/B sky130_fd_sc_hd__xnor2_1
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12106_ _13051_/B _12275_/D _12258_/B _12275_/A vssd1 vssd1 vccd1 vccd1 _12108_/A
+ sky130_fd_sc_hd__a22oi_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10298_ _10419_/B _10421_/D _10297_/D _14789_/A vssd1 vssd1 vccd1 vccd1 _10298_/Y
+ sky130_fd_sc_hd__a22oi_1
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13086_ _13085_/A _13085_/B _13085_/C vssd1 vssd1 vccd1 vccd1 _13220_/A sky130_fd_sc_hd__o21ai_1
XFILLER_97_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12037_ _12037_/A vssd1 vssd1 vccd1 vccd1 _12037_/Y sky130_fd_sc_hd__clkinv_2
X_16914_ _16914_/A _16914_/B vssd1 vssd1 vccd1 vccd1 _16916_/A sky130_fd_sc_hd__nor2_1
XFILLER_78_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_90 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16845_ _16846_/A _16846_/B _16846_/C vssd1 vssd1 vccd1 vccd1 _16909_/A sky130_fd_sc_hd__o21ai_1
XFILLER_92_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16776_ _16777_/A _16777_/B _16777_/C vssd1 vssd1 vccd1 vccd1 _16846_/A sky130_fd_sc_hd__a21oi_1
XFILLER_65_368 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13988_ _13988_/A _13988_/B vssd1 vssd1 vccd1 vccd1 _13989_/B sky130_fd_sc_hd__and2_1
XFILLER_168_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15727_ _16025_/A _16499_/B _16662_/C _15820_/A vssd1 vssd1 vccd1 vccd1 _15728_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_34_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12939_ _12817_/A _12817_/B _12815_/Y vssd1 vssd1 vccd1 vccd1 _12982_/B sky130_fd_sc_hd__a21bo_1
XFILLER_46_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_338 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15658_ _15709_/A _15658_/B vssd1 vssd1 vccd1 vccd1 _15658_/Y sky130_fd_sc_hd__nand2_2
XFILLER_33_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14609_ _14609_/A _14609_/B vssd1 vssd1 vccd1 vccd1 _14610_/B sky130_fd_sc_hd__and2_1
XFILLER_21_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15589_ _15590_/A _15590_/B _15590_/C vssd1 vssd1 vccd1 vccd1 _15591_/A sky130_fd_sc_hd__a21oi_1
X_17328_ _11861_/B _17360_/A2 _17327_/X _17408_/C1 vssd1 vssd1 vccd1 vccd1 _17493_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_119_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17259_ _17563_/Q _17292_/B vssd1 vssd1 vccd1 vccd1 _17259_/X sky130_fd_sc_hd__and2_1
XFILLER_162_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_917 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08963_ _09654_/C _11932_/B _17139_/A _09493_/A vssd1 vssd1 vccd1 vccd1 _08963_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_97_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08894_ _08895_/A _08895_/B vssd1 vssd1 vccd1 vccd1 _08910_/A sky130_fd_sc_hd__nand2b_1
XFILLER_84_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_143 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_36 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09515_ _09514_/B _10203_/B _10067_/B _09797_/A vssd1 vssd1 vccd1 vccd1 _09515_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_71_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_59 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09446_ _09447_/A _09445_/Y _09730_/C _09446_/D vssd1 vssd1 vccd1 vccd1 _09583_/A
+ sky130_fd_sc_hd__and4bb_1
XPHY_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_438 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09377_ _09514_/B _10072_/B _10203_/B _09942_/A vssd1 vssd1 vccd1 vccd1 _09377_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_33_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_871 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11270_ _11270_/A _11270_/B vssd1 vssd1 vccd1 vccd1 _11313_/B sky130_fd_sc_hd__xnor2_1
XFILLER_152_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10221_ _10223_/B _10223_/A vssd1 vssd1 vccd1 vccd1 _10221_/X sky130_fd_sc_hd__and2b_1
XFILLER_106_554 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10152_ _10265_/A _10265_/B vssd1 vssd1 vccd1 vccd1 _10152_/X sky130_fd_sc_hd__and2_1
XFILLER_0_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10083_ _10209_/A _10083_/B vssd1 vssd1 vccd1 vccd1 _10084_/B sky130_fd_sc_hd__or2_1
XFILLER_94_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14960_ _14955_/X _14959_/X _15103_/S vssd1 vssd1 vccd1 vccd1 _15458_/B sky130_fd_sc_hd__mux2_1
X_13911_ _13912_/A _13912_/B vssd1 vssd1 vccd1 vccd1 _14013_/B sky130_fd_sc_hd__or2_1
XFILLER_48_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14891_ _14881_/X _14889_/X _15275_/C1 vssd1 vssd1 vccd1 vccd1 _15081_/A sky130_fd_sc_hd__a21o_2
XFILLER_48_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16630_ _16630_/A _16630_/B _16630_/C vssd1 vssd1 vccd1 vccd1 _16631_/B sky130_fd_sc_hd__and3_1
XFILLER_47_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13842_ _14842_/A1 _13839_/X _13841_/X _14482_/B1 vssd1 vssd1 vccd1 vccd1 _13842_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_114_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwb_buttons_leds_961 vssd1 vssd1 vccd1 vccd1 wb_buttons_leds_961/HI led_enb[3] sky130_fd_sc_hd__conb_1
XFILLER_74_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16561_ _16563_/B _16564_/A _16385_/A vssd1 vssd1 vccd1 vccd1 _16561_/X sky130_fd_sc_hd__or3b_1
X_13773_ _13977_/A _13977_/B _14141_/D _14050_/D vssd1 vssd1 vccd1 vccd1 _13774_/B
+ sky130_fd_sc_hd__and4_1
X_10985_ _10985_/A _10985_/B vssd1 vssd1 vccd1 vccd1 _10987_/B sky130_fd_sc_hd__xnor2_1
XFILLER_55_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15512_ _15512_/A _15512_/B vssd1 vssd1 vccd1 vccd1 _15514_/C sky130_fd_sc_hd__xor2_1
X_12724_ _13028_/A _12877_/C vssd1 vssd1 vccd1 vccd1 _12725_/B sky130_fd_sc_hd__nand2_1
XFILLER_16_788 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_254 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16492_ _16492_/A _16492_/B _16492_/C vssd1 vssd1 vccd1 vccd1 _16493_/C sky130_fd_sc_hd__and3_1
XFILLER_43_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15443_ _15367_/B _15369_/B _15365_/X vssd1 vssd1 vccd1 vccd1 _15443_/X sky130_fd_sc_hd__a21o_1
X_12655_ _12655_/A _12655_/B vssd1 vssd1 vccd1 vccd1 _12671_/A sky130_fd_sc_hd__and2_1
XFILLER_169_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11606_ _11576_/B _11572_/C _11572_/D _11572_/A vssd1 vssd1 vccd1 vccd1 _11607_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_90_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15374_ _15374_/A _15374_/B vssd1 vssd1 vccd1 vccd1 _15374_/X sky130_fd_sc_hd__or2_1
XFILLER_156_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12586_ _12586_/A _12586_/B vssd1 vssd1 vccd1 vccd1 _12588_/C sky130_fd_sc_hd__or2_1
XFILLER_129_646 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17113_ _17113_/A _17113_/B _17113_/C vssd1 vssd1 vccd1 vccd1 _17113_/X sky130_fd_sc_hd__and3_1
XFILLER_157_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14325_ _14325_/A _14325_/B vssd1 vssd1 vccd1 vccd1 _14326_/C sky130_fd_sc_hd__xnor2_1
X_11537_ _11538_/A _11537_/B _11537_/C vssd1 vssd1 vccd1 vccd1 _11538_/B sky130_fd_sc_hd__nor3_1
XFILLER_156_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17044_ _17044_/A _17085_/B vssd1 vssd1 vccd1 vccd1 _17046_/C sky130_fd_sc_hd__nor2_1
Xmax_cap117 wire118/X vssd1 vssd1 vccd1 vccd1 _13713_/A sky130_fd_sc_hd__clkbuf_1
X_14256_ _14258_/A _14258_/B vssd1 vssd1 vccd1 vccd1 _14256_/X sky130_fd_sc_hd__and2_1
X_11468_ _11506_/A _11506_/B _15042_/B _11468_/D vssd1 vssd1 vccd1 vccd1 _11468_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_125_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13207_ _13450_/B _13208_/C _13208_/D _14769_/A vssd1 vssd1 vccd1 vccd1 _13211_/A
+ sky130_fd_sc_hd__a22oi_1
X_10419_ _14789_/A _10419_/B _10534_/D _10899_/D vssd1 vssd1 vccd1 vccd1 _10422_/A
+ sky130_fd_sc_hd__and4_1
X_14187_ _14188_/A _14188_/B _14188_/C vssd1 vssd1 vccd1 vccd1 _14268_/A sky130_fd_sc_hd__a21oi_1
X_11399_ _11399_/A _11399_/B vssd1 vssd1 vccd1 vccd1 _11400_/C sky130_fd_sc_hd__xnor2_1
XFILLER_125_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13138_ _13002_/A _13138_/B vssd1 vssd1 vccd1 vccd1 _13140_/B sky130_fd_sc_hd__and2b_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13069_ _13069_/A _13321_/D vssd1 vssd1 vccd1 vccd1 _13070_/B sky130_fd_sc_hd__nand2_1
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_143 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16828_ _16828_/A _16828_/B vssd1 vssd1 vccd1 vccd1 _16829_/B sky130_fd_sc_hd__nand2_1
XFILLER_66_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16759_ _16759_/A _16759_/B vssd1 vssd1 vccd1 vccd1 _16761_/A sky130_fd_sc_hd__nor2_1
XFILLER_53_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09300_ _09299_/B _09446_/D _11867_/D _17385_/A vssd1 vssd1 vccd1 vccd1 _09300_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_34_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09231_ _09231_/A _09231_/B vssd1 vssd1 vccd1 vccd1 _09240_/A sky130_fd_sc_hd__or2_1
XFILLER_61_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09162_ _09493_/A _11813_/B _08969_/C vssd1 vssd1 vccd1 vccd1 _09163_/B sky130_fd_sc_hd__a21o_1
XFILLER_21_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_966 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09093_ _09093_/A _09093_/B vssd1 vssd1 vccd1 vccd1 _09314_/A sky130_fd_sc_hd__nand2_1
XFILLER_174_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_26 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09995_ _09996_/A _09996_/B vssd1 vssd1 vccd1 vccd1 _10009_/A sky130_fd_sc_hd__nand2b_1
X_08946_ _08946_/A _08946_/B vssd1 vssd1 vccd1 vccd1 _08962_/A sky130_fd_sc_hd__xnor2_1
XFILLER_88_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08877_ _17401_/A _09272_/D _08808_/A _08806_/Y vssd1 vssd1 vccd1 vccd1 _08883_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_85_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_703 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10770_ _10771_/A _10771_/B _10771_/C vssd1 vssd1 vccd1 vccd1 _10777_/A sky130_fd_sc_hd__o21ai_1
XFILLER_13_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09429_ _16990_/A _17038_/B vssd1 vssd1 vccd1 vccd1 _09430_/B sky130_fd_sc_hd__nand2_1
XFILLER_158_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12440_ _12440_/A _12616_/A vssd1 vssd1 vccd1 vccd1 _12442_/C sky130_fd_sc_hd__nor2_1
XFILLER_139_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12371_ _12371_/A _12371_/B vssd1 vssd1 vccd1 vccd1 _12373_/B sky130_fd_sc_hd__nor2_1
XFILLER_154_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14110_ _14015_/B _14110_/B vssd1 vssd1 vccd1 vccd1 _14111_/B sky130_fd_sc_hd__nand2b_1
X_11322_ _11427_/A _11553_/A _11561_/C _11563_/D vssd1 vssd1 vccd1 vccd1 _11325_/A
+ sky130_fd_sc_hd__nand4_1
X_15090_ _15091_/A _15091_/B vssd1 vssd1 vccd1 vccd1 _15170_/A sky130_fd_sc_hd__nand2_1
XFILLER_158_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14041_ _13947_/Y _13951_/B _14040_/X vssd1 vssd1 vccd1 vccd1 _14043_/B sky130_fd_sc_hd__o21a_1
XFILLER_69_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11253_ _11348_/A _11253_/B vssd1 vssd1 vccd1 vccd1 _11288_/A sky130_fd_sc_hd__xor2_1
XFILLER_106_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10204_ _10560_/B _10203_/B _10203_/C vssd1 vssd1 vccd1 vccd1 _10205_/B sky130_fd_sc_hd__a21oi_1
X_11184_ _11039_/Y _11041_/Y _11182_/Y _11183_/X vssd1 vssd1 vccd1 vccd1 _11218_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_122_844 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_395 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10135_ _10134_/A _10134_/Y _10005_/X _10105_/Y vssd1 vssd1 vccd1 vccd1 _10157_/C
+ sky130_fd_sc_hd__a211o_1
X_15992_ _15992_/A _15992_/B _15990_/Y vssd1 vssd1 vccd1 vccd1 _15994_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10066_ _10198_/A _10066_/B vssd1 vssd1 vccd1 vccd1 _10067_/C sky130_fd_sc_hd__xor2_1
X_14943_ _14941_/X _14942_/X _17156_/B vssd1 vssd1 vccd1 vccd1 _14944_/C sky130_fd_sc_hd__a21oi_1
XFILLER_75_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14874_ _15262_/B _14888_/C _14876_/D vssd1 vssd1 vccd1 vccd1 _14874_/X sky130_fd_sc_hd__or3_1
X_16613_ _16697_/B _16613_/B vssd1 vssd1 vccd1 vccd1 _16614_/B sky130_fd_sc_hd__nor2_1
X_13825_ _13827_/B _13827_/A vssd1 vssd1 vccd1 vccd1 _13825_/Y sky130_fd_sc_hd__nand2b_1
X_17593_ fanout933/X _17593_/D vssd1 vssd1 vccd1 vccd1 _17593_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16544_ _16545_/B _16545_/A vssd1 vssd1 vccd1 vccd1 _16544_/X sky130_fd_sc_hd__and2b_1
XFILLER_90_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13756_ _13757_/B _13756_/B vssd1 vssd1 vccd1 vccd1 _13862_/A sky130_fd_sc_hd__and2b_1
X_10968_ _10969_/B _10969_/A vssd1 vssd1 vccd1 vccd1 _11024_/A sky130_fd_sc_hd__and2b_1
XFILLER_16_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12707_ _12703_/X _12706_/X _16012_/S vssd1 vssd1 vccd1 vccd1 _12707_/X sky130_fd_sc_hd__mux2_1
X_16475_ _16475_/A _16475_/B vssd1 vssd1 vccd1 vccd1 _16475_/X sky130_fd_sc_hd__or2_2
XFILLER_43_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13687_ _13787_/A _13687_/B vssd1 vssd1 vccd1 vccd1 _13688_/B sky130_fd_sc_hd__and2_1
XFILLER_31_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10899_ _10995_/A _10898_/Y _10993_/C _10899_/D vssd1 vssd1 vccd1 vccd1 _10995_/B
+ sky130_fd_sc_hd__and4bb_1
X_15426_ _15426_/A _15426_/B vssd1 vssd1 vccd1 vccd1 _15433_/A sky130_fd_sc_hd__xor2_1
XFILLER_129_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12638_ _12788_/A _12942_/D vssd1 vssd1 vccd1 vccd1 _12640_/C sky130_fd_sc_hd__nand2_1
XFILLER_157_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15357_ _16086_/A _15397_/A vssd1 vssd1 vccd1 vccd1 _15358_/B sky130_fd_sc_hd__nand2_1
X_12569_ _12570_/A _12570_/B vssd1 vssd1 vccd1 vccd1 _12730_/B sky130_fd_sc_hd__nand2_1
XFILLER_157_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14308_ _14309_/B _14309_/A vssd1 vssd1 vccd1 vccd1 _14378_/B sky130_fd_sc_hd__nand2b_1
XFILLER_172_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15288_ _15278_/A _16317_/B _15216_/A _15213_/X vssd1 vssd1 vccd1 vccd1 _15291_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_85_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17027_ _11771_/Y _17025_/Y _17026_/Y vssd1 vssd1 vccd1 vccd1 _17033_/A sky130_fd_sc_hd__a21o_1
X_14239_ _14239_/A _14239_/B vssd1 vssd1 vccd1 vccd1 _14258_/A sky130_fd_sc_hd__nor2_1
XFILLER_116_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout708 _17499_/Q vssd1 vssd1 vccd1 vccd1 _10431_/B sky130_fd_sc_hd__clkbuf_4
Xfanout719 _16480_/A vssd1 vssd1 vccd1 vccd1 _13966_/C sky130_fd_sc_hd__buf_4
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08800_ _08801_/A _08801_/B _08801_/C vssd1 vssd1 vccd1 vccd1 _08800_/X sky130_fd_sc_hd__a21o_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09780_ _15254_/S _11808_/B _14952_/A vssd1 vssd1 vccd1 vccd1 _09783_/A sky130_fd_sc_hd__and3_1
XFILLER_112_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08731_ _08731_/A vssd1 vssd1 vccd1 vccd1 _15262_/C sky130_fd_sc_hd__inv_2
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1004 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_338 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09214_ _09214_/A _09214_/B _09214_/C vssd1 vssd1 vccd1 vccd1 _09342_/A sky130_fd_sc_hd__and3_1
XFILLER_50_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09145_ _17415_/A _12129_/B _09145_/C vssd1 vssd1 vccd1 vccd1 _09231_/B sky130_fd_sc_hd__and3_1
XFILLER_148_774 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09076_ _09076_/A _09076_/B _09076_/C vssd1 vssd1 vccd1 vccd1 _09115_/B sky130_fd_sc_hd__and3_1
XFILLER_107_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_844 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09978_ _09983_/A _09983_/B vssd1 vssd1 vccd1 vccd1 _09989_/A sky130_fd_sc_hd__nor2_1
XFILLER_131_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08929_ _08930_/A _08930_/B _08930_/C vssd1 vssd1 vccd1 vccd1 _08929_/Y sky130_fd_sc_hd__nor3_2
XFILLER_76_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11940_ _11941_/A _11941_/B vssd1 vssd1 vccd1 vccd1 _11940_/X sky130_fd_sc_hd__and2_1
XFILLER_91_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11871_ _11871_/A _11871_/B vssd1 vssd1 vccd1 vccd1 _11872_/A sky130_fd_sc_hd__xor2_1
XFILLER_45_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13610_ _13495_/A _13497_/X _13718_/B _13609_/X vssd1 vssd1 vccd1 vccd1 _13612_/A
+ sky130_fd_sc_hd__o211a_1
X_10822_ _10822_/A _11099_/A vssd1 vssd1 vccd1 vccd1 _10829_/B sky130_fd_sc_hd__nor2_1
XTAP_2967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14590_ _14636_/A _14590_/B vssd1 vssd1 vccd1 vccd1 _14590_/Y sky130_fd_sc_hd__nand2_1
XTAP_2989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13541_ _13541_/A _13541_/B vssd1 vssd1 vccd1 vccd1 _13542_/A sky130_fd_sc_hd__xor2_1
X_10753_ _10753_/A _12054_/B _10897_/C vssd1 vssd1 vccd1 vccd1 _10756_/A sky130_fd_sc_hd__and3_1
XFILLER_111_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_875 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16260_ _16352_/A _16259_/B _16259_/C vssd1 vssd1 vccd1 vccd1 _16261_/B sky130_fd_sc_hd__a21oi_1
XFILLER_125_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13472_ _13473_/A _13473_/B vssd1 vssd1 vccd1 vccd1 _13590_/A sky130_fd_sc_hd__and2b_1
XFILLER_41_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10684_ _10575_/Y _10585_/X _10679_/X _10682_/Y vssd1 vssd1 vccd1 vccd1 _10685_/C
+ sky130_fd_sc_hd__a211o_1
X_15211_ _14881_/X _14889_/X _16410_/A _15275_/C1 vssd1 vssd1 vccd1 vccd1 _15494_/A
+ sky130_fd_sc_hd__a211oi_2
X_12423_ _12734_/B _14065_/B _14063_/C _13035_/A vssd1 vssd1 vccd1 vccd1 _12425_/A
+ sky130_fd_sc_hd__a22oi_1
X_16191_ _16191_/A _16191_/B vssd1 vssd1 vccd1 vccd1 _16192_/B sky130_fd_sc_hd__xnor2_1
XFILLER_138_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15142_ _16021_/A _16317_/A _15147_/A vssd1 vssd1 vccd1 vccd1 _15143_/C sky130_fd_sc_hd__o21a_1
XFILLER_138_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12354_ _12354_/A _12354_/B vssd1 vssd1 vccd1 vccd1 _12355_/B sky130_fd_sc_hd__xnor2_1
XFILLER_154_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11305_ _15472_/A _11240_/C _17466_/D _15262_/B vssd1 vssd1 vccd1 vccd1 _11306_/B
+ sky130_fd_sc_hd__a22oi_1
XFILLER_4_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15073_ _14887_/Y _15071_/Y _15715_/A vssd1 vssd1 vccd1 vccd1 _16315_/B sky130_fd_sc_hd__o21ai_4
X_12285_ _12286_/A _12286_/B _12286_/C vssd1 vssd1 vccd1 vccd1 _12476_/A sky130_fd_sc_hd__a21o_1
XFILLER_4_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14024_ _14025_/A _14025_/B vssd1 vssd1 vccd1 vccd1 _14119_/A sky130_fd_sc_hd__nor2_1
X_11236_ _11146_/B _11143_/C _11143_/D _11144_/A vssd1 vssd1 vccd1 vccd1 _11237_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_141_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11167_ _11204_/A _11167_/B vssd1 vssd1 vccd1 vccd1 _11167_/X sky130_fd_sc_hd__and2_1
XFILLER_67_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10118_ _10118_/A _10118_/B vssd1 vssd1 vccd1 vccd1 _10232_/A sky130_fd_sc_hd__xnor2_1
XFILLER_49_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11098_ _11098_/A _11242_/A vssd1 vssd1 vccd1 vccd1 _11101_/B sky130_fd_sc_hd__nor2_1
X_15975_ _15976_/B _15976_/A vssd1 vssd1 vccd1 vccd1 _15975_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_95_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14926_ _16012_/S _15808_/A vssd1 vssd1 vccd1 vccd1 _14926_/X sky130_fd_sc_hd__or2_1
X_10049_ _10053_/A vssd1 vssd1 vccd1 vccd1 _10054_/A sky130_fd_sc_hd__inv_2
XFILLER_76_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14857_ _16014_/A _16014_/B vssd1 vssd1 vccd1 vccd1 _16114_/B sky130_fd_sc_hd__and2_1
XFILLER_17_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13808_ _13809_/A _13809_/B vssd1 vssd1 vccd1 vccd1 _13923_/A sky130_fd_sc_hd__nor2_1
X_14788_ _14788_/A _14788_/B vssd1 vssd1 vccd1 vccd1 _14801_/B sky130_fd_sc_hd__nor2_1
X_17576_ fanout950/X _17576_/D vssd1 vssd1 vccd1 vccd1 _17576_/Q sky130_fd_sc_hd__dfxtp_1
X_16527_ _16527_/A _16527_/B _16527_/C vssd1 vssd1 vccd1 vccd1 _16528_/B sky130_fd_sc_hd__or3_1
XFILLER_149_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13739_ _13739_/A _13739_/B vssd1 vssd1 vccd1 vccd1 _13741_/C sky130_fd_sc_hd__xnor2_1
XFILLER_91_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16458_ _16459_/A _16459_/B vssd1 vssd1 vccd1 vccd1 _16550_/B sky130_fd_sc_hd__nand2_1
X_15409_ _15501_/A _15418_/B vssd1 vssd1 vccd1 vccd1 _15419_/A sky130_fd_sc_hd__nand2b_1
X_16389_ _16389_/A _16389_/B _16389_/C vssd1 vssd1 vccd1 vccd1 _16389_/Y sky130_fd_sc_hd__nand3_2
XFILLER_118_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09901_ _10034_/A _09900_/Y _10045_/C _10311_/D vssd1 vssd1 vccd1 vccd1 _10042_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_125_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout505 _09892_/A vssd1 vssd1 vccd1 vccd1 _17379_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_116_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout516 _12592_/B vssd1 vssd1 vccd1 vccd1 _09892_/B sky130_fd_sc_hd__buf_4
Xfanout527 _17516_/Q vssd1 vssd1 vccd1 vccd1 _11423_/B sky130_fd_sc_hd__clkbuf_2
X_09832_ _09832_/A _09832_/B vssd1 vssd1 vccd1 vccd1 _09914_/A sky130_fd_sc_hd__nor2_1
XFILLER_98_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout538 _15237_/A1 vssd1 vssd1 vccd1 vccd1 _14924_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_86_514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout549 _17514_/Q vssd1 vssd1 vccd1 vccd1 _14925_/A sky130_fd_sc_hd__buf_2
XFILLER_98_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_696 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09763_ _09656_/A _09656_/B _09656_/C vssd1 vssd1 vccd1 vccd1 _09764_/B sky130_fd_sc_hd__o21ai_1
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09694_ _09695_/A _09693_/Y _10366_/A _09838_/C vssd1 vssd1 vccd1 vccd1 _09842_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_55_934 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_820 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_672 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09128_ _09139_/A _09128_/B _17415_/A _09128_/D vssd1 vssd1 vccd1 vccd1 _09139_/B
+ sky130_fd_sc_hd__and4b_1
XFILLER_109_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09059_ _17383_/A _12077_/C _12077_/D _17385_/A vssd1 vssd1 vccd1 vccd1 _09059_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_123_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12070_ _12070_/A _13080_/D _12070_/C _12070_/D vssd1 vssd1 vccd1 vccd1 _12239_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_2_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11021_ _11022_/A _11022_/B vssd1 vssd1 vccd1 vccd1 _11021_/X sky130_fd_sc_hd__or2_1
XFILLER_150_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_94 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15760_ _15760_/A _15760_/B vssd1 vssd1 vccd1 vccd1 _15762_/B sky130_fd_sc_hd__xor2_1
XFILLER_64_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12972_ _12972_/A _12972_/B vssd1 vssd1 vccd1 vccd1 _12974_/B sky130_fd_sc_hd__nor2_1
XTAP_3421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11923_ _11924_/A _11924_/B vssd1 vssd1 vccd1 vccd1 _12179_/B sky130_fd_sc_hd__nor2_1
X_14711_ _14736_/A _14744_/B vssd1 vssd1 vccd1 vccd1 _14712_/B sky130_fd_sc_hd__nor2_1
XTAP_3454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15691_ _15690_/A _15690_/B _15690_/C vssd1 vssd1 vccd1 vccd1 _15691_/Y sky130_fd_sc_hd__o21ai_1
XTAP_3465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17430_ input36/X _17607_/Q _17433_/S vssd1 vssd1 vccd1 vccd1 _17607_/D sky130_fd_sc_hd__mux2_1
X_14642_ _14642_/A _14678_/A vssd1 vssd1 vccd1 vccd1 _14644_/C sky130_fd_sc_hd__nor2_1
XTAP_2764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11854_ _13516_/S _12845_/S _11854_/C vssd1 vssd1 vccd1 vccd1 _11854_/X sky130_fd_sc_hd__or3_2
XFILLER_82_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10805_ _11095_/A _11095_/B _11115_/C _10805_/D vssd1 vssd1 vccd1 vccd1 _10807_/A
+ sky130_fd_sc_hd__and4_1
XTAP_2797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17361_ _17362_/A _17362_/B _17362_/C _17362_/D vssd1 vssd1 vccd1 vccd1 _17361_/Y
+ sky130_fd_sc_hd__nor4_4
X_14573_ _14621_/B _14571_/X _14517_/Y _14519_/X vssd1 vssd1 vccd1 vccd1 _14574_/A
+ sky130_fd_sc_hd__a211oi_1
X_11785_ _09826_/A _14837_/A _12016_/A vssd1 vssd1 vccd1 vccd1 _11785_/X sky130_fd_sc_hd__o21a_1
X_13524_ _13523_/Y _13637_/A _13524_/C vssd1 vssd1 vccd1 vccd1 _13637_/B sky130_fd_sc_hd__nand3b_1
X_16312_ _16298_/A _16494_/B1 _16296_/Y _16311_/X vssd1 vssd1 vccd1 vccd1 _16313_/A
+ sky130_fd_sc_hd__a22o_1
X_10736_ _11115_/A _11115_/B _10970_/B _10736_/D vssd1 vssd1 vccd1 vccd1 _10739_/A
+ sky130_fd_sc_hd__and4_1
X_17292_ _17574_/Q _17292_/B vssd1 vssd1 vccd1 vccd1 _17292_/X sky130_fd_sc_hd__and2_1
XFILLER_40_171 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16243_ _16149_/X _16153_/B _16245_/A _16040_/B vssd1 vssd1 vccd1 vccd1 _16252_/A
+ sky130_fd_sc_hd__a2bb2o_1
X_13455_ _13455_/A _13455_/B _13455_/C vssd1 vssd1 vccd1 vccd1 _13457_/A sky130_fd_sc_hd__or3_1
XFILLER_51_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10667_ _10667_/A _10667_/B _10667_/C vssd1 vssd1 vccd1 vccd1 _10667_/Y sky130_fd_sc_hd__nor3_2
XFILLER_9_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12406_ _12406_/A _12561_/A vssd1 vssd1 vccd1 vccd1 _12408_/C sky130_fd_sc_hd__nor2_1
X_16174_ _16174_/A _16174_/B vssd1 vssd1 vccd1 vccd1 _16175_/B sky130_fd_sc_hd__xor2_1
X_13386_ _13509_/A _13386_/B vssd1 vssd1 vccd1 vccd1 _13388_/B sky130_fd_sc_hd__nand2_1
X_10598_ _10599_/A _10599_/B vssd1 vssd1 vccd1 vccd1 _10598_/X sky130_fd_sc_hd__or2_1
X_15125_ _15131_/A _15125_/B vssd1 vssd1 vccd1 vccd1 _15125_/Y sky130_fd_sc_hd__nand2_1
Xoutput108 _17465_/Q vssd1 vssd1 vccd1 vccd1 o_wb_data[31] sky130_fd_sc_hd__clkbuf_1
X_12337_ _17417_/A _12338_/C _12338_/D _17419_/A vssd1 vssd1 vccd1 vccd1 _12339_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_154_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15056_ _15056_/A _15056_/B vssd1 vssd1 vccd1 vccd1 _15056_/Y sky130_fd_sc_hd__nor2_1
X_12268_ _12268_/A _12268_/B _12268_/C vssd1 vssd1 vccd1 vccd1 _12268_/X sky130_fd_sc_hd__and3_1
XFILLER_142_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14007_ _14007_/A _14007_/B vssd1 vssd1 vccd1 vccd1 _14008_/C sky130_fd_sc_hd__xnor2_1
X_11219_ _11220_/A _11220_/B vssd1 vssd1 vccd1 vccd1 _11219_/Y sky130_fd_sc_hd__nand2_1
XFILLER_141_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12199_ _12198_/A _12198_/B _12198_/C vssd1 vssd1 vccd1 vccd1 _12201_/B sky130_fd_sc_hd__o21ai_1
Xoutput90 _17449_/Q vssd1 vssd1 vccd1 vccd1 o_wb_data[15] sky130_fd_sc_hd__clkbuf_1
XFILLER_150_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_366 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15958_ _15853_/B _15955_/Y _15957_/X vssd1 vssd1 vccd1 vccd1 _15960_/A sky130_fd_sc_hd__a21o_1
XFILLER_37_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14909_ _15553_/A _15553_/B vssd1 vssd1 vccd1 vccd1 _15820_/A sky130_fd_sc_hd__or2_2
X_15889_ _15889_/A _15889_/B vssd1 vssd1 vccd1 vccd1 _15889_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_91_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17559_ fanout952/X _17559_/D vssd1 vssd1 vccd1 vccd1 _17559_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_834 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_703 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_254 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout302 _17369_/A vssd1 vssd1 vccd1 vccd1 _15901_/S sky130_fd_sc_hd__buf_2
XFILLER_87_812 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout313 _15270_/A vssd1 vssd1 vccd1 vccd1 _08731_/A sky130_fd_sc_hd__buf_2
XFILLER_101_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout324 _17541_/Q vssd1 vssd1 vccd1 vccd1 _14832_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_99_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout335 _17540_/Q vssd1 vssd1 vccd1 vccd1 _08988_/B sky130_fd_sc_hd__buf_4
XFILLER_59_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_791 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout346 _17538_/Q vssd1 vssd1 vccd1 vccd1 _14765_/A sky130_fd_sc_hd__clkbuf_4
Xfanout357 _17537_/Q vssd1 vssd1 vccd1 vccd1 _09172_/A sky130_fd_sc_hd__buf_2
X_09815_ _09811_/A _09811_/B _09777_/A vssd1 vssd1 vccd1 vccd1 _09828_/A sky130_fd_sc_hd__a21o_1
XFILLER_113_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout368 _17535_/Q vssd1 vssd1 vccd1 vccd1 _17413_/A sky130_fd_sc_hd__clkbuf_4
Xfanout379 fanout380/X vssd1 vssd1 vccd1 vccd1 _14770_/A sky130_fd_sc_hd__buf_2
XFILLER_115_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09746_ _09746_/A _09754_/A _09746_/C vssd1 vssd1 vccd1 vccd1 _09747_/B sky130_fd_sc_hd__or3_1
XFILLER_39_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09677_ _09677_/A vssd1 vssd1 vccd1 vccd1 _09679_/A sky130_fd_sc_hd__inv_2
XTAP_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11570_ _11526_/B _11552_/X _11557_/X _11603_/A vssd1 vssd1 vccd1 vccd1 _11572_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_35_1047 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_666 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10521_ _10437_/A _10437_/B _10437_/C vssd1 vssd1 vccd1 vccd1 _10521_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_11_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13240_ _13241_/A _13241_/B vssd1 vssd1 vccd1 vccd1 _13240_/Y sky130_fd_sc_hd__nand2b_1
X_10452_ _10453_/A _10453_/B _10453_/C vssd1 vssd1 vccd1 vccd1 _10454_/A sky130_fd_sc_hd__a21o_1
XFILLER_164_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13171_ _13302_/A _14181_/B vssd1 vssd1 vccd1 vccd1 _13172_/B sky130_fd_sc_hd__nand2_1
X_10383_ _10383_/A _10383_/B _10383_/C vssd1 vssd1 vccd1 vccd1 _10385_/C sky130_fd_sc_hd__nand3_1
XFILLER_151_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12122_ _12122_/A _12122_/B _12309_/B _12122_/D vssd1 vssd1 vccd1 vccd1 _12122_/Y
+ sky130_fd_sc_hd__nand4_4
XFILLER_124_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16930_ _16911_/Y _16917_/Y _16929_/X _17170_/B1 _13993_/B vssd1 vssd1 vccd1 vccd1
+ _17568_/D sky130_fd_sc_hd__a32oi_1
X_12053_ _14911_/B _12053_/B vssd1 vssd1 vccd1 vccd1 _12053_/Y sky130_fd_sc_hd__nand2_1
XFILLER_77_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11004_ _11157_/A _11002_/Y _10941_/Y _10946_/X vssd1 vssd1 vccd1 vccd1 _11055_/B
+ sky130_fd_sc_hd__a211o_1
X_16861_ _16792_/A _16792_/B _16788_/Y vssd1 vssd1 vccd1 vccd1 _16863_/B sky130_fd_sc_hd__a21o_1
XFILLER_77_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_366 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout880 _11427_/C vssd1 vssd1 vccd1 vccd1 _15110_/A sky130_fd_sc_hd__clkbuf_4
Xfanout891 _10111_/D vssd1 vssd1 vccd1 vccd1 _10446_/B sky130_fd_sc_hd__clkbuf_4
X_15812_ _16015_/A _15898_/B _15811_/Y _15810_/X vssd1 vssd1 vccd1 vccd1 _15812_/X
+ sky130_fd_sc_hd__o31a_1
X_16792_ _16792_/A _16792_/B vssd1 vssd1 vccd1 vccd1 _16793_/B sky130_fd_sc_hd__xnor2_1
XFILLER_18_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15743_ _15743_/A _15743_/B vssd1 vssd1 vccd1 vccd1 _15765_/A sky130_fd_sc_hd__xor2_1
X_12955_ _12954_/B _12955_/B vssd1 vssd1 vccd1 vccd1 _12956_/B sky130_fd_sc_hd__nand2b_1
XTAP_3251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_252 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11906_ _11906_/A _11906_/B vssd1 vssd1 vccd1 vccd1 _11908_/B sky130_fd_sc_hd__xnor2_1
XTAP_3284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15674_ _15675_/A _15675_/B vssd1 vssd1 vccd1 vccd1 _15674_/X sky130_fd_sc_hd__and2_1
X_12886_ _12886_/A _12886_/B _12886_/C vssd1 vssd1 vccd1 vccd1 _12899_/B sky130_fd_sc_hd__or3_1
XTAP_2550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17413_ _17413_/A _17421_/B vssd1 vssd1 vccd1 vccd1 _17413_/X sky130_fd_sc_hd__or2_1
XFILLER_33_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11837_ _11837_/A _11837_/B vssd1 vssd1 vccd1 vccd1 _11837_/Y sky130_fd_sc_hd__nand2_1
X_14625_ _14660_/B _14625_/B vssd1 vssd1 vccd1 vccd1 _14627_/C sky130_fd_sc_hd__nor2_1
XTAP_2594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17344_ _11900_/D _17356_/A2 _17343_/X _17406_/C1 vssd1 vssd1 vccd1 vccd1 _17501_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14556_ _14557_/A _14557_/B _14557_/C vssd1 vssd1 vccd1 vccd1 _14558_/A sky130_fd_sc_hd__o21a_1
X_11768_ _11768_/A _11768_/B vssd1 vssd1 vccd1 vccd1 _16921_/A sky130_fd_sc_hd__or2_1
XFILLER_159_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10719_ _10720_/A _10718_/Y _10719_/C _10875_/C vssd1 vssd1 vccd1 vccd1 _11013_/A
+ sky130_fd_sc_hd__and4bb_1
X_13507_ _13619_/A _13507_/B vssd1 vssd1 vccd1 vccd1 _13514_/A sky130_fd_sc_hd__nand2_1
XFILLER_158_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17275_ _17459_/Q _17275_/A2 _17273_/X _17274_/X _17275_/C1 vssd1 vssd1 vccd1 vccd1
+ _17459_/D sky130_fd_sc_hd__o221a_1
X_14487_ _14676_/A _14593_/D vssd1 vssd1 vccd1 vccd1 _14489_/B sky130_fd_sc_hd__nand2_1
X_11699_ _11586_/A _11586_/C _11586_/B vssd1 vssd1 vccd1 vccd1 _11700_/C sky130_fd_sc_hd__a21o_1
XFILLER_173_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16226_ _16880_/A _16226_/B _16226_/C _17119_/C vssd1 vssd1 vccd1 vccd1 _16227_/B
+ sky130_fd_sc_hd__and4_1
X_13438_ _13438_/A _13438_/B vssd1 vssd1 vccd1 vccd1 _13439_/B sky130_fd_sc_hd__and2_1
XFILLER_139_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16157_ _16157_/A _16157_/B vssd1 vssd1 vccd1 vccd1 _16158_/B sky130_fd_sc_hd__xnor2_1
XFILLER_6_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13369_ _13369_/A _13369_/B _13369_/C vssd1 vssd1 vccd1 vccd1 _13496_/A sky130_fd_sc_hd__and3_1
XFILLER_154_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15108_ _15108_/A _15108_/B vssd1 vssd1 vccd1 vccd1 _15108_/Y sky130_fd_sc_hd__nand2_1
X_16088_ _16197_/B _16088_/B vssd1 vssd1 vccd1 vccd1 _16089_/B sky130_fd_sc_hd__or2_1
XFILLER_103_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15039_ _15056_/A _14956_/Y _15038_/Y _15097_/A vssd1 vssd1 vccd1 vccd1 _15039_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_102_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_878 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09600_ _09580_/X _09597_/B _09599_/Y _09480_/X vssd1 vssd1 vccd1 vccd1 _09629_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_68_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09531_ _09485_/X _09530_/X _09393_/X _09398_/Y vssd1 vssd1 vccd1 vccd1 _09531_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_3_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09462_ _09462_/A _09468_/A _09462_/C vssd1 vssd1 vccd1 vccd1 _09463_/B sky130_fd_sc_hd__or3_1
XFILLER_51_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09393_ _09395_/B _09393_/B _09393_/C _09393_/D vssd1 vssd1 vccd1 vccd1 _09393_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_33_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout132 _16606_/B vssd1 vssd1 vccd1 vccd1 _16760_/B sky130_fd_sc_hd__clkbuf_4
Xfanout143 _15020_/X vssd1 vssd1 vccd1 vccd1 _16129_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_86_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout154 _15846_/A vssd1 vssd1 vccd1 vccd1 _16056_/A sky130_fd_sc_hd__buf_2
Xfanout165 _17308_/A2 vssd1 vssd1 vccd1 vccd1 _17360_/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_86_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout176 _15575_/Y vssd1 vssd1 vccd1 vccd1 _16814_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_101_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout187 _16595_/A vssd1 vssd1 vccd1 vccd1 _16416_/A sky130_fd_sc_hd__clkbuf_4
Xfanout198 _14758_/A vssd1 vssd1 vccd1 vccd1 _14482_/B1 sky130_fd_sc_hd__buf_2
XFILLER_86_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09729_ _09728_/B _10036_/D _10016_/D _09873_/A vssd1 vssd1 vccd1 vccd1 _09729_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_28_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12740_ _12741_/A _12741_/B vssd1 vssd1 vccd1 vccd1 _12903_/B sky130_fd_sc_hd__and2b_1
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_22 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12671_ _12671_/A _12671_/B vssd1 vssd1 vccd1 vccd1 _12673_/B sky130_fd_sc_hd__xnor2_1
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14410_ _14473_/A _14409_/C _14409_/A vssd1 vssd1 vccd1 vccd1 _14411_/B sky130_fd_sc_hd__a21o_1
X_11622_ _11622_/A _11622_/B vssd1 vssd1 vccd1 vccd1 _15614_/A sky130_fd_sc_hd__or2_1
XFILLER_24_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15390_ _15390_/A _15390_/B vssd1 vssd1 vccd1 vccd1 _15390_/Y sky130_fd_sc_hd__nand2_1
XFILLER_11_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14341_ _14340_/B _14340_/C _14340_/A vssd1 vssd1 vccd1 vccd1 _14342_/B sky130_fd_sc_hd__a21o_1
X_11553_ _11553_/A _11553_/B _11629_/D _11605_/B vssd1 vssd1 vccd1 vccd1 _11637_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_7_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17060_ _17060_/A _17060_/B vssd1 vssd1 vccd1 vccd1 _17062_/B sky130_fd_sc_hd__nor2_1
X_10504_ _10719_/C _10525_/D _10395_/A _10393_/Y vssd1 vssd1 vccd1 vccd1 _10505_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_155_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14272_ _14273_/A _14273_/B _14273_/C vssd1 vssd1 vccd1 vccd1 _14350_/B sky130_fd_sc_hd__a21oi_1
XFILLER_155_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11484_ _11484_/A _11484_/B _11522_/A vssd1 vssd1 vccd1 vccd1 _11485_/B sky130_fd_sc_hd__or3_1
XFILLER_144_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16011_ _16011_/A _16011_/B _16011_/C vssd1 vssd1 vccd1 vccd1 _16011_/X sky130_fd_sc_hd__or3_1
XFILLER_171_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13223_ _16649_/A _13223_/B vssd1 vssd1 vccd1 vccd1 _13224_/B sky130_fd_sc_hd__nand2_1
XFILLER_6_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10435_ _10436_/B _10436_/A vssd1 vssd1 vccd1 vccd1 _10563_/A sky130_fd_sc_hd__and2b_1
XFILLER_124_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13154_ _13154_/A _13154_/B vssd1 vssd1 vccd1 vccd1 _13161_/A sky130_fd_sc_hd__xnor2_1
X_10366_ _10366_/A _11027_/C _10709_/A vssd1 vssd1 vccd1 vccd1 _10367_/B sky130_fd_sc_hd__and3_1
XFILLER_3_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12105_ _12105_/A _12105_/B vssd1 vssd1 vccd1 vccd1 _12115_/A sky130_fd_sc_hd__xnor2_1
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13085_ _13085_/A _13085_/B _13085_/C vssd1 vssd1 vccd1 vccd1 _13087_/A sky130_fd_sc_hd__or3_1
XFILLER_88_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10297_ _14789_/A _10419_/B _10421_/D _10297_/D vssd1 vssd1 vccd1 vccd1 _10300_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_33_8 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12036_ _15384_/S _12034_/X _12035_/X vssd1 vssd1 vccd1 vccd1 _12037_/A sky130_fd_sc_hd__o21ai_2
X_16913_ _13993_/B _16965_/B _16913_/C vssd1 vssd1 vccd1 vccd1 _16914_/B sky130_fd_sc_hd__and3b_1
XFILLER_78_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16844_ _16906_/B _16844_/B vssd1 vssd1 vccd1 vccd1 _16846_/C sky130_fd_sc_hd__and2_1
XFILLER_78_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16775_ _16775_/A _16775_/B vssd1 vssd1 vccd1 vccd1 _16777_/C sky130_fd_sc_hd__xnor2_1
X_13987_ _13988_/A _13988_/B vssd1 vssd1 vccd1 vccd1 _14077_/A sky130_fd_sc_hd__nor2_1
XFILLER_92_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15726_ _15726_/A _15918_/A _16591_/B _16743_/C vssd1 vssd1 vccd1 vccd1 _15834_/A
+ sky130_fd_sc_hd__and4_1
XTAP_3081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12938_ _12938_/A _12938_/B _12938_/C vssd1 vssd1 vccd1 vccd1 _12985_/B sky130_fd_sc_hd__and3_1
XFILLER_33_200 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15657_ _15709_/A _15658_/B vssd1 vssd1 vccd1 vccd1 _16743_/B sky130_fd_sc_hd__and2_2
XFILLER_22_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12869_ _12869_/A _13348_/B _12869_/C vssd1 vssd1 vccd1 vccd1 _12870_/B sky130_fd_sc_hd__and3_1
XTAP_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14608_ _14609_/A _14609_/B vssd1 vssd1 vccd1 vccd1 _14683_/A sky130_fd_sc_hd__nor2_1
XTAP_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15588_ _15588_/A _15588_/B vssd1 vssd1 vccd1 vccd1 _15590_/C sky130_fd_sc_hd__xnor2_1
X_17327_ input42/X _17359_/B _17359_/C vssd1 vssd1 vccd1 vccd1 _17327_/X sky130_fd_sc_hd__or3_1
XFILLER_147_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14539_ _14629_/A _14629_/B vssd1 vssd1 vccd1 vccd1 _14585_/B sky130_fd_sc_hd__nand2_1
XFILLER_146_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17258_ _17595_/Q _17291_/A2 _17291_/B1 vssd1 vssd1 vccd1 vccd1 _17258_/X sky130_fd_sc_hd__a21o_1
XFILLER_174_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16209_ _14859_/B _16209_/B _16209_/C vssd1 vssd1 vccd1 vccd1 _16210_/B sky130_fd_sc_hd__and3b_1
XFILLER_128_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17189_ input30/X input34/X input5/X input4/X vssd1 vssd1 vccd1 vccd1 _17191_/C sky130_fd_sc_hd__or4_1
XFILLER_108_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_929 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08962_ _08962_/A _08962_/B _08962_/C vssd1 vssd1 vccd1 vccd1 _08985_/B sky130_fd_sc_hd__and3_1
XFILLER_102_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08893_ _08893_/A _08893_/B vssd1 vssd1 vccd1 vccd1 _08895_/B sky130_fd_sc_hd__xnor2_1
XFILLER_57_804 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_995 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09514_ _09797_/A _09514_/B _10203_/B _10067_/B vssd1 vssd1 vccd1 vccd1 _09517_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_140_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_188 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09445_ _09728_/B _09042_/B _12500_/B _09873_/A vssd1 vssd1 vccd1 vccd1 _09445_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_24_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09376_ _09942_/A _09514_/B _10072_/B _10203_/B vssd1 vssd1 vccd1 vccd1 _09379_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_166_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_883 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10220_ _10219_/A _10342_/A vssd1 vssd1 vccd1 vccd1 _10223_/B sky130_fd_sc_hd__and2b_1
XFILLER_106_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10151_ _10151_/A _10151_/B vssd1 vssd1 vccd1 vccd1 _10265_/B sky130_fd_sc_hd__nor2_1
X_10082_ _10209_/A _10083_/B vssd1 vssd1 vccd1 vccd1 _10084_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13910_ _14027_/B _13910_/B vssd1 vssd1 vccd1 vccd1 _13912_/B sky130_fd_sc_hd__or2_1
XFILLER_87_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14890_ _14881_/X _14889_/X _15275_/C1 vssd1 vssd1 vccd1 vccd1 _14890_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_75_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13841_ _13841_/A _14839_/B vssd1 vssd1 vccd1 vccd1 _13841_/X sky130_fd_sc_hd__or2_1
XFILLER_114_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xwb_buttons_leds_962 vssd1 vssd1 vccd1 vccd1 wb_buttons_leds_962/HI led_enb[4] sky130_fd_sc_hd__conb_1
XFILLER_56_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16560_ _16560_/A _16560_/B vssd1 vssd1 vccd1 vccd1 _16566_/A sky130_fd_sc_hd__nand2_2
X_13772_ _13977_/B _14141_/D _14050_/D _13977_/A vssd1 vssd1 vccd1 vccd1 _13774_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_74_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10984_ _10984_/A _10985_/A _10984_/C vssd1 vssd1 vccd1 vccd1 _11162_/A sky130_fd_sc_hd__or3_1
XFILLER_15_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15511_ _15512_/A _15512_/B vssd1 vssd1 vccd1 vccd1 _15511_/X sky130_fd_sc_hd__and2b_1
XFILLER_16_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12723_ _12723_/A _12723_/B vssd1 vssd1 vccd1 vccd1 _12725_/A sky130_fd_sc_hd__nor2_1
XFILLER_43_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16491_ _17143_/A1 _14127_/X _16582_/A _15104_/X vssd1 vssd1 vccd1 vccd1 _16492_/C
+ sky130_fd_sc_hd__o22a_1
XFILLER_15_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12654_ _12654_/A _12654_/B vssd1 vssd1 vccd1 vccd1 _12655_/B sky130_fd_sc_hd__nand2_1
XFILLER_43_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15442_ _15442_/A _15442_/B vssd1 vssd1 vccd1 vccd1 _15442_/Y sky130_fd_sc_hd__xnor2_1
X_11605_ _15305_/C _11605_/B _11610_/B _11605_/D vssd1 vssd1 vccd1 vccd1 _11607_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_169_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12585_ _12585_/A _12585_/B _12585_/C vssd1 vssd1 vccd1 vccd1 _12586_/B sky130_fd_sc_hd__and3_1
X_15373_ _15381_/A _15373_/B _15373_/C vssd1 vssd1 vccd1 vccd1 _15374_/B sky130_fd_sc_hd__and3b_1
XFILLER_157_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17112_ _17112_/A1 _17164_/C _15252_/X _17143_/A1 _14705_/B vssd1 vssd1 vccd1 vccd1
+ _17113_/C sky130_fd_sc_hd__o32a_1
X_11536_ _11532_/A _11532_/B _11574_/A vssd1 vssd1 vccd1 vccd1 _11537_/C sky130_fd_sc_hd__o21ba_1
XFILLER_129_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14324_ _14324_/A _14389_/B _14325_/B vssd1 vssd1 vccd1 vccd1 _14393_/A sky130_fd_sc_hd__or3_1
XFILLER_23_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_966 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_606 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17043_ _17119_/A _17043_/B _17043_/C vssd1 vssd1 vccd1 vccd1 _17085_/B sky130_fd_sc_hd__and3_1
X_14255_ _14255_/A _14255_/B vssd1 vssd1 vccd1 vccd1 _14258_/B sky130_fd_sc_hd__xnor2_1
X_11467_ _11506_/A _11506_/B _11592_/B _11468_/D vssd1 vssd1 vccd1 vccd1 _11472_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_7_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13206_ _13578_/A _13564_/C vssd1 vssd1 vccd1 vccd1 _16649_/A sky130_fd_sc_hd__nand2_2
XFILLER_109_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10418_ _10418_/A _10423_/A _10418_/C vssd1 vssd1 vccd1 vccd1 _10427_/B sky130_fd_sc_hd__or3_1
X_14186_ _14186_/A _14186_/B vssd1 vssd1 vccd1 vccd1 _14188_/C sky130_fd_sc_hd__or2_1
X_11398_ _11403_/A _11368_/Y _11384_/Y _11396_/X vssd1 vssd1 vccd1 vccd1 _11400_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_140_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13137_ _13137_/A _13137_/B vssd1 vssd1 vccd1 vccd1 _13268_/B sky130_fd_sc_hd__nand2_1
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10349_ _10349_/A _10349_/B vssd1 vssd1 vccd1 vccd1 _10350_/B sky130_fd_sc_hd__and2_1
XFILLER_97_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_247 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13068_ _13068_/A _13068_/B vssd1 vssd1 vccd1 vccd1 _13070_/A sky130_fd_sc_hd__nor2_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12019_ _12025_/A _10308_/B _14956_/A vssd1 vssd1 vccd1 vccd1 _12020_/B sky130_fd_sc_hd__a21o_1
XFILLER_94_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16827_ _16827_/A _16827_/B _16827_/C _16827_/D vssd1 vssd1 vccd1 vccd1 _16828_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_65_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16758_ _16758_/A _16758_/B _16758_/C vssd1 vssd1 vccd1 vccd1 _16759_/B sky130_fd_sc_hd__and3_1
XFILLER_0_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15709_ _15709_/A _15709_/B vssd1 vssd1 vccd1 vccd1 _15710_/C sky130_fd_sc_hd__nor2_1
X_16689_ _16690_/A _16690_/B vssd1 vssd1 vccd1 vccd1 _16770_/B sky130_fd_sc_hd__and2b_1
XFILLER_110_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09230_ _09230_/A _09230_/B vssd1 vssd1 vccd1 vccd1 _09248_/A sky130_fd_sc_hd__xnor2_1
XFILLER_167_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09161_ _09164_/A vssd1 vssd1 vccd1 vccd1 _09161_/Y sky130_fd_sc_hd__inv_2
XFILLER_119_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09092_ _09092_/A vssd1 vssd1 vccd1 vccd1 _09093_/B sky130_fd_sc_hd__inv_2
XFILLER_135_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09994_ _09994_/A _16809_/B vssd1 vssd1 vccd1 vccd1 _09996_/B sky130_fd_sc_hd__xnor2_2
XFILLER_115_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_878 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08945_ _08945_/A _08945_/B vssd1 vssd1 vccd1 vccd1 _08946_/B sky130_fd_sc_hd__xnor2_1
X_08876_ _08876_/A _08876_/B vssd1 vssd1 vccd1 vccd1 _08904_/A sky130_fd_sc_hd__xnor2_1
XFILLER_151_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09428_ _10255_/A _10899_/D vssd1 vssd1 vccd1 vccd1 _16990_/B sky130_fd_sc_hd__nand2_2
XFILLER_40_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09359_ _09366_/A _09366_/B _09366_/C vssd1 vssd1 vccd1 vccd1 _09370_/B sky130_fd_sc_hd__a21o_1
XFILLER_139_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12370_ _12370_/A _12370_/B vssd1 vssd1 vccd1 vccd1 _12373_/A sky130_fd_sc_hd__xnor2_1
XFILLER_121_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11321_ _14889_/C _15151_/B vssd1 vssd1 vccd1 vccd1 _11321_/X sky130_fd_sc_hd__and2_1
XFILLER_158_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14040_ _13950_/A _13948_/C _14181_/B _13948_/A vssd1 vssd1 vccd1 vccd1 _14040_/X
+ sky130_fd_sc_hd__a22o_1
X_11252_ _11252_/A _11252_/B vssd1 vssd1 vccd1 vccd1 _11253_/B sky130_fd_sc_hd__xnor2_1
XFILLER_158_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_83 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10203_ _10560_/B _10203_/B _10203_/C vssd1 vssd1 vccd1 vccd1 _10469_/B sky130_fd_sc_hd__and3_1
XFILLER_106_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11183_ _11182_/A _11182_/B _11182_/C vssd1 vssd1 vccd1 vccd1 _11183_/X sky130_fd_sc_hd__o21a_1
XFILLER_134_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10134_ _10134_/A _10134_/B _10134_/C vssd1 vssd1 vccd1 vccd1 _10134_/Y sky130_fd_sc_hd__nand3_2
XFILLER_0_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15991_ _15992_/A _15992_/B _15990_/Y vssd1 vssd1 vccd1 vccd1 _15991_/X sky130_fd_sc_hd__o21ba_1
XFILLER_48_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10065_ _10198_/A _10066_/B vssd1 vssd1 vccd1 vccd1 _10069_/B sky130_fd_sc_hd__and2_1
X_14942_ _14942_/A _15553_/A _15450_/B vssd1 vssd1 vccd1 vccd1 _14942_/X sky130_fd_sc_hd__or3_1
XFILLER_47_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14873_ _16021_/A _14873_/B _17613_/Q vssd1 vssd1 vccd1 vccd1 _14876_/D sky130_fd_sc_hd__or3b_1
XFILLER_63_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_86 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16612_ _16611_/B _16612_/B vssd1 vssd1 vccd1 vccd1 _16613_/B sky130_fd_sc_hd__and2b_1
XFILLER_29_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13824_ _13824_/A _13824_/B vssd1 vssd1 vccd1 vccd1 _13827_/B sky130_fd_sc_hd__nand2_1
X_17592_ fanout933/X _17592_/D vssd1 vssd1 vccd1 vccd1 _17592_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16543_ _16543_/A _16543_/B vssd1 vssd1 vccd1 vccd1 _16545_/B sky130_fd_sc_hd__xnor2_1
XFILLER_16_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10967_ _10915_/A _10914_/B _10914_/A vssd1 vssd1 vccd1 vccd1 _10969_/B sky130_fd_sc_hd__o21ba_1
X_13755_ _13650_/B _13652_/B _13648_/X vssd1 vssd1 vccd1 vccd1 _13757_/B sky130_fd_sc_hd__a21oi_1
XFILLER_50_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12706_ _12704_/X _12705_/X _13627_/S vssd1 vssd1 vccd1 vccd1 _12706_/X sky130_fd_sc_hd__mux2_1
XFILLER_149_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16474_ _16563_/A _16384_/Y _16472_/X _15523_/A vssd1 vssd1 vccd1 vccd1 _16475_/B
+ sky130_fd_sc_hd__a31o_1
X_10898_ _10991_/A _10897_/B _10897_/C vssd1 vssd1 vccd1 vccd1 _10898_/Y sky130_fd_sc_hd__a21oi_1
X_13686_ _13686_/A _13686_/B vssd1 vssd1 vccd1 vccd1 _13687_/B sky130_fd_sc_hd__nand2_1
X_15425_ _15426_/A _15426_/B vssd1 vssd1 vccd1 vccd1 _15514_/A sky130_fd_sc_hd__nand2_1
X_12637_ _17413_/A _12787_/B _12787_/D _12637_/D vssd1 vssd1 vccd1 vccd1 _12792_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_15_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_904 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12568_ _12568_/A _12568_/B vssd1 vssd1 vccd1 vccd1 _12570_/B sky130_fd_sc_hd__xnor2_1
X_15356_ _15356_/A _15356_/B vssd1 vssd1 vccd1 vccd1 _15358_/A sky130_fd_sc_hd__nand2_1
XFILLER_172_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_926 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11519_ _11518_/B _11518_/C _11563_/D _11518_/A vssd1 vssd1 vccd1 vccd1 _11519_/Y
+ sky130_fd_sc_hd__a22oi_1
X_14307_ _14225_/A _16970_/A _14225_/B vssd1 vssd1 vccd1 vccd1 _14309_/B sky130_fd_sc_hd__o21ba_1
XFILLER_171_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12499_ _12499_/A _12499_/B vssd1 vssd1 vccd1 vccd1 _12501_/A sky130_fd_sc_hd__nor2_1
X_15287_ _15287_/A _15287_/B vssd1 vssd1 vccd1 vccd1 _15292_/A sky130_fd_sc_hd__xor2_1
XFILLER_172_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17026_ _11771_/Y _17025_/Y _16922_/A vssd1 vssd1 vccd1 vccd1 _17026_/Y sky130_fd_sc_hd__o21ai_1
X_14238_ _14237_/A _14237_/B _14236_/X vssd1 vssd1 vccd1 vccd1 _14239_/B sky130_fd_sc_hd__o21ba_1
XFILLER_125_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_160 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14169_ _14170_/A _14245_/A _14170_/C vssd1 vssd1 vccd1 vccd1 _14171_/A sky130_fd_sc_hd__o21a_1
XFILLER_98_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout709 _13968_/B vssd1 vssd1 vccd1 vccd1 _14141_/D sky130_fd_sc_hd__clkbuf_4
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08730_ input70/X vssd1 vssd1 vccd1 vccd1 _17428_/B sky130_fd_sc_hd__clkinv_4
XFILLER_61_1032 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09213_ _09213_/A _09213_/B vssd1 vssd1 vccd1 vccd1 _09214_/C sky130_fd_sc_hd__xnor2_1
XFILLER_22_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09144_ _09502_/A _12129_/B _09145_/C vssd1 vssd1 vccd1 vccd1 _09147_/B sky130_fd_sc_hd__a21oi_1
XFILLER_163_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_606 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09075_ _09076_/A _09076_/B _09076_/C vssd1 vssd1 vccd1 vccd1 _09115_/A sky130_fd_sc_hd__a21oi_2
XFILLER_30_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_918 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09977_ _10111_/C _09979_/C _09841_/A _09839_/Y vssd1 vssd1 vccd1 vccd1 _09983_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_39_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08928_ _08832_/Y _08875_/X _08905_/A _09051_/A vssd1 vssd1 vccd1 vccd1 _08930_/C
+ sky130_fd_sc_hd__o211a_1
XTAP_3603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08859_ _08859_/A _08859_/B vssd1 vssd1 vccd1 vccd1 _08861_/A sky130_fd_sc_hd__nor2_1
XFILLER_45_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11870_ _17393_/A _12077_/C _11871_/A vssd1 vssd1 vccd1 vccd1 _12093_/B sky130_fd_sc_hd__and3_1
XFILLER_45_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10821_ _10822_/A _10820_/Y _11097_/C _17469_/D vssd1 vssd1 vccd1 vccd1 _11099_/A
+ sky130_fd_sc_hd__and4bb_1
XTAP_2957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_990 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10752_ _11651_/A _10993_/D vssd1 vssd1 vccd1 vccd1 _10897_/C sky130_fd_sc_hd__and2_2
X_13540_ _13658_/A _13852_/B _13657_/B vssd1 vssd1 vccd1 vccd1 _13541_/B sky130_fd_sc_hd__and3_1
XFILLER_71_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13471_ _13471_/A _13471_/B vssd1 vssd1 vccd1 vccd1 _13473_/B sky130_fd_sc_hd__xnor2_1
XFILLER_41_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10683_ _10679_/X _10682_/Y _10575_/Y _10585_/X vssd1 vssd1 vccd1 vccd1 _10685_/B
+ sky130_fd_sc_hd__o211ai_2
X_15210_ _15203_/X _15208_/X _14906_/B vssd1 vssd1 vccd1 vccd1 _16138_/A sky130_fd_sc_hd__a21bo_2
X_12422_ _12257_/A _12259_/B _12257_/B vssd1 vssd1 vccd1 vccd1 _12432_/A sky130_fd_sc_hd__o21ba_1
XFILLER_40_386 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16190_ _16281_/A _16533_/B vssd1 vssd1 vccd1 vccd1 _16191_/B sky130_fd_sc_hd__nand2_1
XFILLER_154_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15141_ _15270_/A _15270_/B vssd1 vssd1 vccd1 vccd1 _15393_/B sky130_fd_sc_hd__or2_1
XFILLER_5_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12353_ _12353_/A _12353_/B vssd1 vssd1 vccd1 vccd1 _12354_/B sky130_fd_sc_hd__and2_1
X_11304_ _11304_/A _11304_/B vssd1 vssd1 vccd1 vccd1 _11364_/A sky130_fd_sc_hd__nor2_1
XFILLER_5_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15072_ _14887_/Y _15071_/Y _15715_/A vssd1 vssd1 vccd1 vccd1 _15074_/B sky130_fd_sc_hd__o21a_1
X_12284_ _12284_/A _12284_/B vssd1 vssd1 vccd1 vccd1 _12286_/C sky130_fd_sc_hd__or2_1
XFILLER_153_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14023_ _13809_/A _13809_/B _13923_/B _13922_/A vssd1 vssd1 vccd1 vccd1 _14025_/B
+ sky130_fd_sc_hd__o31a_1
X_11235_ _11153_/B _11151_/C _11151_/B vssd1 vssd1 vccd1 vccd1 _11235_/X sky130_fd_sc_hd__o21a_1
XFILLER_106_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_171 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11166_ _11165_/A _11165_/B _11165_/C vssd1 vssd1 vccd1 vccd1 _11167_/B sky130_fd_sc_hd__o21ai_1
XFILLER_1_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10117_ _10244_/A _10799_/B vssd1 vssd1 vccd1 vccd1 _10118_/B sky130_fd_sc_hd__nand2_1
XFILLER_96_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11097_ _11098_/A _11096_/Y _11097_/C _17468_/D vssd1 vssd1 vccd1 vccd1 _11242_/A
+ sky130_fd_sc_hd__and4bb_1
X_15974_ _15840_/Y _15864_/B _15839_/Y vssd1 vssd1 vccd1 vccd1 _15976_/B sky130_fd_sc_hd__a21oi_1
XFILLER_49_976 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14925_ _14925_/A _15808_/A vssd1 vssd1 vccd1 vccd1 _14925_/Y sky130_fd_sc_hd__nor2_1
X_10048_ _10050_/B _10163_/A _10050_/A vssd1 vssd1 vccd1 vccd1 _10053_/A sky130_fd_sc_hd__a21o_1
XFILLER_48_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14856_ _15898_/A _15811_/A _15811_/B vssd1 vssd1 vccd1 vccd1 _16014_/B sky130_fd_sc_hd__and3_1
XFILLER_90_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13807_ _13688_/A _13688_/B _13706_/Y vssd1 vssd1 vccd1 vccd1 _13809_/B sky130_fd_sc_hd__a21boi_1
XFILLER_90_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17575_ fanout941/X _17575_/D vssd1 vssd1 vccd1 vccd1 _17575_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14787_ _14787_/A _15381_/A vssd1 vssd1 vccd1 vccd1 _14803_/A sky130_fd_sc_hd__nor2_1
XFILLER_16_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11999_ _11998_/A _11998_/B _12197_/B _11998_/D vssd1 vssd1 vccd1 vccd1 _11999_/Y
+ sky130_fd_sc_hd__o22ai_1
XFILLER_50_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16526_ _16527_/A _16527_/B _16527_/C vssd1 vssd1 vccd1 vccd1 _16630_/A sky130_fd_sc_hd__o21ai_1
X_13738_ _13846_/A _13738_/B _13739_/A vssd1 vssd1 vccd1 vccd1 _13849_/B sky130_fd_sc_hd__and3_1
X_16457_ _16457_/A _16457_/B vssd1 vssd1 vccd1 vccd1 _16459_/B sky130_fd_sc_hd__xnor2_1
X_13669_ _13778_/B _13669_/B vssd1 vssd1 vccd1 vccd1 _13671_/C sky130_fd_sc_hd__nor2_1
XFILLER_84_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15408_ _15408_/A _15408_/B _15408_/C vssd1 vssd1 vccd1 vccd1 _15418_/B sky130_fd_sc_hd__or3_1
XFILLER_118_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16388_ _16387_/B _16387_/C _16387_/A vssd1 vssd1 vccd1 vccd1 _16389_/C sky130_fd_sc_hd__o21ai_1
XFILLER_157_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15339_ _15206_/X _15338_/Y _15381_/A vssd1 vssd1 vccd1 vccd1 _15339_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_144_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17009_ _17037_/A _17009_/B vssd1 vssd1 vccd1 vccd1 _17010_/B sky130_fd_sc_hd__nand2_1
X_09900_ _10419_/B _10543_/B _10657_/B _14789_/A vssd1 vssd1 vccd1 vccd1 _09900_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_104_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout506 _09892_/A vssd1 vssd1 vccd1 vccd1 _09078_/A sky130_fd_sc_hd__clkbuf_2
Xfanout517 _17517_/Q vssd1 vssd1 vccd1 vccd1 _12592_/B sky130_fd_sc_hd__buf_4
X_09831_ _09740_/A _09740_/B _09740_/C vssd1 vssd1 vccd1 vccd1 _09832_/B sky130_fd_sc_hd__a21oi_1
Xfanout528 _10970_/A vssd1 vssd1 vccd1 vccd1 _14788_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_112_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout539 _15237_/A1 vssd1 vssd1 vccd1 vccd1 _11427_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_59_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09762_ _09762_/A _09762_/B _09891_/A vssd1 vssd1 vccd1 vccd1 _09765_/B sky130_fd_sc_hd__nand3_1
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09693_ _10236_/B _09937_/B _09979_/C _10236_/A vssd1 vssd1 vccd1 vccd1 _09693_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_66_272 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_915 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09127_ _17419_/A _17417_/A _12127_/D _11920_/D vssd1 vssd1 vccd1 vccd1 _09139_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_135_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09058_ _17385_/A _17383_/A _09058_/C _12077_/D vssd1 vssd1 vccd1 vccd1 _09061_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_135_255 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11020_ _11020_/A _11020_/B vssd1 vssd1 vccd1 vccd1 _11022_/B sky130_fd_sc_hd__xnor2_1
XFILLER_150_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1041 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12971_ _12971_/A _12971_/B vssd1 vssd1 vccd1 vccd1 _12974_/A sky130_fd_sc_hd__xor2_1
XTAP_3422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14710_ _14719_/A _14710_/B _14710_/C vssd1 vssd1 vccd1 vccd1 _14744_/B sky130_fd_sc_hd__and3b_1
XTAP_3444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11922_ _11922_/A _12127_/C vssd1 vssd1 vccd1 vccd1 _11924_/B sky130_fd_sc_hd__nand2_1
XFILLER_85_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15690_ _15690_/A _15690_/B _15690_/C vssd1 vssd1 vccd1 vccd1 _15779_/B sky130_fd_sc_hd__or3_1
XTAP_3466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14641_ _14641_/A _14641_/B _14641_/C _14641_/D vssd1 vssd1 vccd1 vccd1 _14678_/A
+ sky130_fd_sc_hd__and4_1
XTAP_3499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11853_ _14757_/S _13626_/B vssd1 vssd1 vccd1 vccd1 _11853_/Y sky130_fd_sc_hd__nand2_1
XTAP_2765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10804_ _11097_/C _11117_/D vssd1 vssd1 vccd1 vccd1 _10808_/A sky130_fd_sc_hd__nand2_1
X_17360_ _12592_/C _17360_/A2 _17359_/X _17426_/C1 vssd1 vssd1 vccd1 vccd1 _17509_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_82_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14572_ _14517_/Y _14519_/X _14621_/B _14571_/X vssd1 vssd1 vccd1 vccd1 _14624_/A
+ sky130_fd_sc_hd__o211ai_1
X_11784_ _14872_/A _14924_/C vssd1 vssd1 vccd1 vccd1 _11784_/X sky130_fd_sc_hd__or2_1
XFILLER_159_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16311_ _08743_/A _16293_/Y _16301_/Y _16111_/A _16310_/X vssd1 vssd1 vccd1 vccd1
+ _16311_/X sky130_fd_sc_hd__o221a_1
X_13523_ _13846_/A _13632_/D vssd1 vssd1 vccd1 vccd1 _13523_/Y sky130_fd_sc_hd__nand2_1
X_10735_ _10735_/A _10735_/B vssd1 vssd1 vccd1 vccd1 _10750_/A sky130_fd_sc_hd__xnor2_1
XFILLER_15_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17291_ _17606_/Q _17291_/A2 _17291_/B1 vssd1 vssd1 vccd1 vccd1 _17291_/X sky130_fd_sc_hd__a21o_1
X_16242_ _16347_/A _16242_/B vssd1 vssd1 vccd1 vccd1 _16254_/A sky130_fd_sc_hd__nand2b_1
XFILLER_40_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10666_ _10519_/Y _10588_/X _10632_/A _10632_/Y vssd1 vssd1 vccd1 vccd1 _10667_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_40_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13454_ _13454_/A _13569_/B vssd1 vssd1 vccd1 vccd1 _13455_/C sky130_fd_sc_hd__nor2_1
XFILLER_139_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12405_ _12714_/A _12869_/A _13334_/C _13208_/D vssd1 vssd1 vccd1 vccd1 _12561_/A
+ sky130_fd_sc_hd__and4_1
X_16173_ _16355_/A _16065_/B _16066_/A _16064_/A vssd1 vssd1 vccd1 vccd1 _16174_/B
+ sky130_fd_sc_hd__a31o_1
X_13385_ _13509_/B _13385_/B vssd1 vssd1 vccd1 vccd1 _13508_/B sky130_fd_sc_hd__nor2_1
XFILLER_154_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10597_ _10597_/A _10597_/B vssd1 vssd1 vccd1 vccd1 _10599_/B sky130_fd_sc_hd__xnor2_1
XFILLER_12_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15124_ _10142_/B _10014_/D _10146_/B _10016_/D _14914_/S _10545_/C vssd1 vssd1 vccd1
+ vccd1 _15125_/B sky130_fd_sc_hd__mux4_1
Xoutput109 _17437_/Q vssd1 vssd1 vccd1 vccd1 o_wb_data[3] sky130_fd_sc_hd__clkbuf_1
X_12336_ _12336_/A _12336_/B vssd1 vssd1 vccd1 vccd1 _12354_/A sky130_fd_sc_hd__nor2_1
XFILLER_5_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_91 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12267_ _12268_/A _12268_/B _12268_/C vssd1 vssd1 vccd1 vccd1 _12267_/Y sky130_fd_sc_hd__a21oi_2
X_15055_ _15628_/A _16219_/A1 _12063_/X _15054_/X vssd1 vssd1 vccd1 vccd1 _15055_/X
+ sky130_fd_sc_hd__o31a_1
X_11218_ _11218_/A _11218_/B vssd1 vssd1 vccd1 vccd1 _11220_/B sky130_fd_sc_hd__nand2_1
X_14006_ _14007_/A _14007_/B vssd1 vssd1 vccd1 vccd1 _14115_/A sky130_fd_sc_hd__nand2b_1
X_12198_ _12198_/A _12198_/B _12198_/C vssd1 vssd1 vccd1 vccd1 _12367_/B sky130_fd_sc_hd__or3_1
XFILLER_68_504 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput80 _17473_/Q vssd1 vssd1 vccd1 vccd1 leds[7] sky130_fd_sc_hd__clkbuf_1
Xoutput91 _17450_/Q vssd1 vssd1 vccd1 vccd1 o_wb_data[16] sky130_fd_sc_hd__clkbuf_1
XFILLER_122_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11149_ _11154_/A _11149_/B vssd1 vssd1 vccd1 vccd1 _11151_/B sky130_fd_sc_hd__nand2_1
XFILLER_95_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15957_ _16168_/A _16667_/A _16062_/C vssd1 vssd1 vccd1 vccd1 _15957_/X sky130_fd_sc_hd__o21ba_1
XFILLER_95_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14908_ _15553_/A _15553_/B vssd1 vssd1 vccd1 vccd1 _15475_/A sky130_fd_sc_hd__nor2_1
X_15888_ _15888_/A _15888_/B vssd1 vssd1 vccd1 vccd1 _15889_/B sky130_fd_sc_hd__nand2_1
XFILLER_64_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14839_ _14925_/A _14839_/B vssd1 vssd1 vccd1 vccd1 _14839_/Y sky130_fd_sc_hd__nor2_1
XFILLER_91_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_139 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17558_ fanout954/X _17558_/D vssd1 vssd1 vccd1 vccd1 _17558_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16509_ _16509_/A _16509_/B _16509_/C vssd1 vssd1 vccd1 vccd1 _16510_/B sky130_fd_sc_hd__and3_1
XFILLER_20_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17489_ fanout943/X _17489_/D vssd1 vssd1 vccd1 vccd1 _17489_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_846 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout303 _15116_/A vssd1 vssd1 vccd1 vccd1 _17369_/A sky130_fd_sc_hd__clkbuf_4
Xfanout314 _15071_/A vssd1 vssd1 vccd1 vccd1 _15270_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_99_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout325 _12770_/A vssd1 vssd1 vccd1 vccd1 _17425_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_59_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout336 _13069_/A vssd1 vssd1 vccd1 vccd1 _14215_/A sky130_fd_sc_hd__clkbuf_4
Xfanout347 _12804_/A vssd1 vssd1 vccd1 vccd1 _17419_/A sky130_fd_sc_hd__clkbuf_4
X_09814_ _09772_/X _09813_/X _09668_/Y _09683_/X vssd1 vssd1 vccd1 vccd1 _09814_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_100_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout358 _16965_/C vssd1 vssd1 vccd1 vccd1 _14155_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_140_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout369 _12487_/A vssd1 vssd1 vccd1 vccd1 _09942_/A sky130_fd_sc_hd__buf_2
XFILLER_28_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09745_ _09621_/X _09743_/Y _09740_/B _09724_/X vssd1 vssd1 vccd1 vccd1 _09745_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_39_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09676_ _09678_/B _09681_/A _09678_/A vssd1 vssd1 vccd1 vccd1 _09677_/A sky130_fd_sc_hd__o21ai_1
XFILLER_28_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10520_ _10519_/A _10519_/Y _10406_/B _10474_/Y vssd1 vssd1 vccd1 vccd1 _10555_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_168_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10451_ _10451_/A _10451_/B vssd1 vssd1 vccd1 vccd1 _10453_/C sky130_fd_sc_hd__or2_1
XFILLER_6_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13170_ _13170_/A _13170_/B vssd1 vssd1 vccd1 vccd1 _13172_/A sky130_fd_sc_hd__nor2_1
XFILLER_109_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10382_ _10382_/A _10382_/B vssd1 vssd1 vccd1 vccd1 _10385_/B sky130_fd_sc_hd__xnor2_1
X_12121_ _12122_/A _12122_/B _12309_/B _12122_/D vssd1 vssd1 vccd1 vccd1 _12121_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_123_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12052_ _12025_/A _10993_/D _10991_/C vssd1 vssd1 vccd1 vccd1 _12053_/B sky130_fd_sc_hd__a21o_1
XFILLER_78_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11003_ _10941_/Y _10946_/X _11157_/A _11002_/Y vssd1 vssd1 vccd1 vccd1 _11157_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_78_846 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16860_ _14383_/A _16859_/Y _16858_/Y vssd1 vssd1 vccd1 vccd1 _16863_/A sky130_fd_sc_hd__a21oi_2
XFILLER_104_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout870 fanout874/X vssd1 vssd1 vccd1 vccd1 _11563_/D sky130_fd_sc_hd__buf_2
X_15811_ _15811_/A _15811_/B vssd1 vssd1 vccd1 vccd1 _15811_/Y sky130_fd_sc_hd__nor2_1
Xfanout881 _11427_/C vssd1 vssd1 vccd1 vccd1 _11561_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_77_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout892 _17480_/Q vssd1 vssd1 vccd1 vccd1 _10111_/D sky130_fd_sc_hd__clkbuf_4
X_16791_ _16791_/A _16791_/B vssd1 vssd1 vccd1 vccd1 _16792_/B sky130_fd_sc_hd__nand2_1
XFILLER_46_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15742_ _15742_/A _15742_/B _15743_/B vssd1 vssd1 vccd1 vccd1 _15866_/A sky130_fd_sc_hd__nor3_1
XTAP_3241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12954_ _12955_/B _12954_/B vssd1 vssd1 vccd1 vccd1 _12956_/A sky130_fd_sc_hd__nand2b_1
XFILLER_18_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11905_ _11906_/B _11906_/A vssd1 vssd1 vccd1 vccd1 _11905_/X sky130_fd_sc_hd__and2b_1
XTAP_3285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15673_ _15673_/A _15673_/B vssd1 vssd1 vccd1 vccd1 _15675_/B sky130_fd_sc_hd__xnor2_1
XFILLER_45_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12885_ _12886_/A _12886_/B _12886_/C vssd1 vssd1 vccd1 vccd1 _13049_/A sky130_fd_sc_hd__o21ai_2
XTAP_2551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17412_ input52/X _17426_/A2 _17411_/X _17426_/C1 vssd1 vssd1 vccd1 vccd1 _17534_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_45_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14624_ _14624_/A _14624_/B vssd1 vssd1 vccd1 vccd1 _14625_/B sky130_fd_sc_hd__and2_1
XTAP_2573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11836_ _12637_/D _12487_/D _11839_/S vssd1 vssd1 vccd1 vccd1 _11837_/B sky130_fd_sc_hd__mux2_1
XTAP_2584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17343_ input51/X _17353_/B _17353_/C vssd1 vssd1 vccd1 vccd1 _17343_/X sky130_fd_sc_hd__or3_1
XTAP_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14555_ _14555_/A _14555_/B vssd1 vssd1 vccd1 vccd1 _14557_/C sky130_fd_sc_hd__xnor2_1
XTAP_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11767_ _11768_/A _11767_/B vssd1 vssd1 vccd1 vccd1 _11767_/X sky130_fd_sc_hd__or2_1
XFILLER_9_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13506_ _13506_/A _13506_/B vssd1 vssd1 vccd1 vccd1 _13507_/B sky130_fd_sc_hd__or2_1
X_10718_ _09299_/B _10962_/B _14849_/A _10142_/A vssd1 vssd1 vccd1 vccd1 _10718_/Y
+ sky130_fd_sc_hd__a22oi_1
X_17274_ _17568_/Q _17274_/B vssd1 vssd1 vccd1 vccd1 _17274_/X sky130_fd_sc_hd__and2_1
X_14486_ _14486_/A _14557_/A vssd1 vssd1 vccd1 vccd1 _14489_/A sky130_fd_sc_hd__or2_1
X_11698_ _11622_/B _15614_/B _11622_/A vssd1 vssd1 vccd1 vccd1 _11700_/B sky130_fd_sc_hd__o21bai_1
XFILLER_158_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16225_ _16315_/B _16827_/C _16938_/D _15734_/A vssd1 vssd1 vccd1 vccd1 _16227_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_173_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13437_ _13438_/A _13438_/B vssd1 vssd1 vccd1 vccd1 _13586_/B sky130_fd_sc_hd__nor2_1
X_10649_ _10649_/A _10649_/B vssd1 vssd1 vccd1 vccd1 _10735_/B sky130_fd_sc_hd__xnor2_1
XFILLER_6_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16156_ _16157_/B _16157_/A vssd1 vssd1 vccd1 vccd1 _16270_/B sky130_fd_sc_hd__and2b_1
X_13368_ _13368_/A _13368_/B vssd1 vssd1 vccd1 vccd1 _13369_/C sky130_fd_sc_hd__or2_1
XFILLER_155_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15107_ _11472_/B _14791_/X _14797_/X vssd1 vssd1 vccd1 vccd1 _15108_/B sky130_fd_sc_hd__a21o_1
X_12319_ _12787_/B _12487_/D _12320_/D _17413_/A vssd1 vssd1 vccd1 vccd1 _12323_/A
+ sky130_fd_sc_hd__a22oi_1
X_16087_ _16281_/A _16355_/B _16086_/C vssd1 vssd1 vccd1 vccd1 _16088_/B sky130_fd_sc_hd__a21oi_1
XFILLER_115_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13299_ _13658_/A _14094_/B _13657_/B vssd1 vssd1 vccd1 vccd1 _13301_/A sky130_fd_sc_hd__a21boi_1
XFILLER_5_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15038_ _15056_/A _15038_/B vssd1 vssd1 vccd1 vccd1 _15038_/Y sky130_fd_sc_hd__nor2_1
XFILLER_142_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16989_ _16989_/A _16989_/B vssd1 vssd1 vccd1 vccd1 _16991_/C sky130_fd_sc_hd__or2_1
XFILLER_110_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09530_ _09485_/X _09530_/B _09530_/C _09530_/D vssd1 vssd1 vccd1 vccd1 _09530_/X
+ sky130_fd_sc_hd__and4b_1
XFILLER_3_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09461_ _09335_/A _09459_/Y _09455_/B _09440_/X vssd1 vssd1 vccd1 vccd1 _09461_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_25_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09392_ _09395_/B _09393_/B _09393_/C _09393_/D vssd1 vssd1 vccd1 vccd1 _09395_/C
+ sky130_fd_sc_hd__nor4_1
XFILLER_52_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_895 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout133 _15755_/B vssd1 vssd1 vccd1 vccd1 _16667_/A sky130_fd_sc_hd__clkbuf_4
Xfanout144 _16165_/A vssd1 vssd1 vccd1 vccd1 _15750_/A sky130_fd_sc_hd__clkbuf_4
Xfanout155 _14890_/Y vssd1 vssd1 vccd1 vccd1 _15846_/A sky130_fd_sc_hd__buf_2
Xfanout166 _17296_/Y vssd1 vssd1 vccd1 vccd1 _17308_/A2 sky130_fd_sc_hd__clkbuf_4
Xfanout177 _16514_/A vssd1 vssd1 vccd1 vccd1 _16827_/B sky130_fd_sc_hd__buf_2
XFILLER_86_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout188 _15263_/Y vssd1 vssd1 vccd1 vccd1 _16533_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_47_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout199 _15457_/B vssd1 vssd1 vccd1 vccd1 _12710_/A sky130_fd_sc_hd__buf_2
XFILLER_28_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09728_ _09873_/A _09728_/B _10036_/D _10532_/D vssd1 vssd1 vccd1 vccd1 _09731_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_16_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09659_ _09788_/A _09788_/B vssd1 vssd1 vccd1 vccd1 _09789_/A sky130_fd_sc_hd__nor2_2
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_34 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12670_ _12670_/A _12670_/B vssd1 vssd1 vccd1 vccd1 _12671_/B sky130_fd_sc_hd__xor2_1
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_919 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11621_ _11620_/A _11620_/C _11624_/A vssd1 vssd1 vccd1 vccd1 _11622_/B sky130_fd_sc_hd__o21a_1
XFILLER_30_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_470 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14340_ _14340_/A _14340_/B _14340_/C vssd1 vssd1 vccd1 vccd1 _14342_/A sky130_fd_sc_hd__nand3_1
X_11552_ _11526_/A _11525_/C _11525_/B vssd1 vssd1 vccd1 vccd1 _11552_/X sky130_fd_sc_hd__a21o_1
XFILLER_128_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10503_ _10503_/A _10503_/B _10503_/C vssd1 vssd1 vccd1 vccd1 _10503_/Y sky130_fd_sc_hd__nand3_1
XFILLER_10_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11483_ _11484_/B _11522_/A _11484_/A vssd1 vssd1 vccd1 vccd1 _11534_/A sky130_fd_sc_hd__o21ai_1
XFILLER_7_636 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14271_ _14350_/A _14271_/B vssd1 vssd1 vccd1 vccd1 _14273_/C sky130_fd_sc_hd__or2_1
XFILLER_137_851 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16010_ _15034_/Y _15037_/X _15039_/X _15057_/X _15312_/S _15901_/S vssd1 vssd1 vccd1
+ vccd1 _16010_/X sky130_fd_sc_hd__mux4_1
XFILLER_155_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13222_ _16649_/A _13223_/B vssd1 vssd1 vccd1 vccd1 _13224_/A sky130_fd_sc_hd__or2_1
X_10434_ _10434_/A _10547_/A vssd1 vssd1 vccd1 vccd1 _10436_/B sky130_fd_sc_hd__nor2_1
XFILLER_171_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13153_ _13154_/B _13154_/A vssd1 vssd1 vccd1 vccd1 _13295_/A sky130_fd_sc_hd__nand2b_1
X_10365_ _10236_/X _10365_/B vssd1 vssd1 vccd1 vccd1 _10370_/C sky130_fd_sc_hd__and2b_1
XFILLER_98_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12104_ _17375_/A _12439_/D vssd1 vssd1 vccd1 vccd1 _12105_/B sky130_fd_sc_hd__nand2_1
XFILLER_2_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13084_ _13084_/A _13213_/B vssd1 vssd1 vccd1 vccd1 _13085_/C sky130_fd_sc_hd__nor2_1
XFILLER_124_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10296_ _10296_/A _10301_/A _10296_/C vssd1 vssd1 vccd1 vccd1 _10305_/B sky130_fd_sc_hd__or3_1
XFILLER_151_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12035_ _12845_/S _14948_/A _12035_/C vssd1 vssd1 vccd1 vccd1 _12035_/X sky130_fd_sc_hd__or3_1
X_16912_ _16913_/C _16965_/B _13993_/B vssd1 vssd1 vccd1 vccd1 _16914_/A sky130_fd_sc_hd__a21boi_1
XFILLER_78_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16843_ _16843_/A _16843_/B vssd1 vssd1 vccd1 vccd1 _16844_/B sky130_fd_sc_hd__or2_1
XFILLER_65_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16774_ _16774_/A _16774_/B vssd1 vssd1 vccd1 vccd1 _16775_/B sky130_fd_sc_hd__xnor2_1
XFILLER_168_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13986_ _13986_/A _13986_/B vssd1 vssd1 vccd1 vccd1 _13988_/B sky130_fd_sc_hd__nor2_1
XFILLER_46_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15725_ _16136_/A _16054_/B vssd1 vssd1 vccd1 vccd1 _16497_/C sky130_fd_sc_hd__nand2_1
XFILLER_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12937_ _12985_/A vssd1 vssd1 vccd1 vccd1 _13125_/A sky130_fd_sc_hd__inv_2
XTAP_3071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15656_ _15656_/A _15656_/B vssd1 vssd1 vccd1 vccd1 _15679_/A sky130_fd_sc_hd__xnor2_1
X_12868_ _12869_/A _13348_/B _12869_/C vssd1 vssd1 vccd1 vccd1 _12870_/A sky130_fd_sc_hd__a21oi_1
XTAP_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14607_ _14558_/B _14560_/B _14558_/A vssd1 vssd1 vccd1 vccd1 _14609_/B sky130_fd_sc_hd__o21ba_1
X_11819_ _17367_/A _12700_/B _12546_/C _11818_/Y vssd1 vssd1 vccd1 vccd1 _11820_/A
+ sky130_fd_sc_hd__a31o_2
XFILLER_33_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15587_ _15685_/B _15587_/B vssd1 vssd1 vccd1 vccd1 _15588_/B sky130_fd_sc_hd__xnor2_1
X_12799_ _12799_/A _12799_/B vssd1 vssd1 vccd1 vccd1 _12801_/A sky130_fd_sc_hd__nor2_1
XTAP_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17326_ _11859_/D _17360_/A2 _17325_/X _17408_/C1 vssd1 vssd1 vccd1 vccd1 _17492_/D
+ sky130_fd_sc_hd__o211a_1
X_14538_ _14629_/A _14629_/B vssd1 vssd1 vccd1 vccd1 _14538_/X sky130_fd_sc_hd__or2_1
XFILLER_174_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17257_ _17453_/Q _17290_/A2 _17255_/X _17256_/X _17293_/C1 vssd1 vssd1 vccd1 vccd1
+ _17453_/D sky130_fd_sc_hd__o221a_1
XFILLER_174_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14469_ _14469_/A _14469_/B vssd1 vssd1 vccd1 vccd1 _14471_/B sky130_fd_sc_hd__xnor2_1
XFILLER_88_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16208_ _16209_/C _16209_/B _14859_/B vssd1 vssd1 vccd1 vccd1 _16300_/A sky130_fd_sc_hd__a21boi_1
XFILLER_134_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17188_ input15/X input20/X input22/X input21/X vssd1 vssd1 vccd1 vccd1 _17191_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_108_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16139_ _16140_/A _16140_/B vssd1 vssd1 vccd1 vccd1 _16250_/B sky130_fd_sc_hd__and2b_1
XFILLER_143_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08961_ _08962_/B _08962_/C _08962_/A vssd1 vssd1 vccd1 vccd1 _08985_/A sky130_fd_sc_hd__a21oi_1
XFILLER_103_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_1014 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08892_ _16315_/A _08887_/A _08887_/B vssd1 vssd1 vccd1 vccd1 _08895_/A sky130_fd_sc_hd__o21ba_1
XFILLER_151_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09513_ _09513_/A _09513_/B vssd1 vssd1 vccd1 vccd1 _09519_/A sky130_fd_sc_hd__nor2_1
XFILLER_37_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09444_ _09873_/A _09728_/B _11867_/D _12500_/B vssd1 vssd1 vccd1 vccd1 _09447_/A
+ sky130_fd_sc_hd__and4_1
XPHY_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09375_ _09375_/A _09375_/B vssd1 vssd1 vccd1 vccd1 _09381_/A sky130_fd_sc_hd__nor2_1
XFILLER_71_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10150_ _14788_/A _11841_/B _10039_/A _10037_/Y vssd1 vssd1 vccd1 vccd1 _10151_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_161_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_695 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10081_ _10081_/A _10081_/B vssd1 vssd1 vccd1 vccd1 _10083_/B sky130_fd_sc_hd__and2_1
XFILLER_0_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13840_ _12862_/X _12866_/B _13840_/S vssd1 vssd1 vccd1 vccd1 _14839_/B sky130_fd_sc_hd__mux2_1
XFILLER_28_551 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwb_buttons_leds_963 vssd1 vssd1 vccd1 vccd1 wb_buttons_leds_963/HI led_enb[5] sky130_fd_sc_hd__conb_1
XFILLER_16_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13771_ _13921_/A _13771_/B vssd1 vssd1 vccd1 vccd1 _13812_/A sky130_fd_sc_hd__nand2_1
X_10983_ _10984_/A _10984_/C vssd1 vssd1 vccd1 vccd1 _10985_/B sky130_fd_sc_hd__nor2_1
XFILLER_15_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_1002 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15510_ _15510_/A _15510_/B vssd1 vssd1 vccd1 vccd1 _15512_/B sky130_fd_sc_hd__xor2_1
XFILLER_16_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12722_ _12722_/A _12722_/B _13464_/B _13348_/B vssd1 vssd1 vccd1 vccd1 _12723_/B
+ sky130_fd_sc_hd__and4_1
X_16490_ _12560_/A _17163_/A2 _16489_/X vssd1 vssd1 vccd1 vccd1 _16492_/B sky130_fd_sc_hd__o21ba_1
XFILLER_128_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15441_ _15442_/A _15442_/B vssd1 vssd1 vccd1 vccd1 _15441_/X sky130_fd_sc_hd__and2b_1
XFILLER_130_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12653_ _12654_/A _12654_/B vssd1 vssd1 vccd1 vccd1 _12655_/A sky130_fd_sc_hd__or2_1
XFILLER_169_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11604_ _11603_/A _11603_/C _11603_/B vssd1 vssd1 vccd1 vccd1 _11605_/D sky130_fd_sc_hd__o21ai_1
XFILLER_129_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15372_ _17377_/A _15450_/B _15381_/A vssd1 vssd1 vccd1 vccd1 _15374_/A sky130_fd_sc_hd__o21a_1
X_12584_ _12585_/A _12585_/B _12585_/C vssd1 vssd1 vccd1 vccd1 _12586_/A sky130_fd_sc_hd__a21oi_1
XFILLER_30_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17111_ _14596_/Y _17163_/A2 _17110_/X _16977_/A vssd1 vssd1 vccd1 vccd1 _17113_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_90_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14323_ _14242_/A _14244_/B _14242_/B vssd1 vssd1 vccd1 vccd1 _14325_/B sky130_fd_sc_hd__o21ba_1
X_11535_ _11541_/A _11535_/B vssd1 vssd1 vccd1 vccd1 _11537_/B sky130_fd_sc_hd__nand2_1
XFILLER_11_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_618 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17042_ _17119_/A _16987_/B _17043_/C vssd1 vssd1 vccd1 vccd1 _17044_/A sky130_fd_sc_hd__a21oi_1
XFILLER_7_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14254_ _14254_/A _14450_/B vssd1 vssd1 vccd1 vccd1 _14255_/B sky130_fd_sc_hd__nand2_1
X_11466_ _11444_/A _11444_/C _11444_/B vssd1 vssd1 vccd1 vccd1 _11466_/X sky130_fd_sc_hd__a21o_1
XFILLER_156_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xmax_cap119 _13494_/B vssd1 vssd1 vccd1 vccd1 _13376_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_99_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13205_ _13201_/Y _13203_/A _13075_/A _13075_/Y vssd1 vssd1 vccd1 vccd1 _13249_/B
+ sky130_fd_sc_hd__o211ai_2
X_10417_ _10418_/A _10418_/C vssd1 vssd1 vccd1 vccd1 _10423_/B sky130_fd_sc_hd__nor2_1
X_11397_ _11384_/Y _11396_/X _11403_/A _11368_/Y vssd1 vssd1 vccd1 vccd1 _11403_/B
+ sky130_fd_sc_hd__o211ai_1
X_14185_ _14185_/A _14185_/B vssd1 vssd1 vccd1 vccd1 _14186_/B sky130_fd_sc_hd__nor2_1
XFILLER_125_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13136_ _13136_/A vssd1 vssd1 vccd1 vccd1 _13137_/B sky130_fd_sc_hd__inv_2
XFILLER_140_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10348_ _10348_/A _10348_/B _10348_/C vssd1 vssd1 vccd1 vccd1 _11775_/B sky130_fd_sc_hd__or3_1
XFILLER_124_386 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13067_ _13434_/A _14050_/B _13194_/D _13067_/D vssd1 vssd1 vccd1 vccd1 _13068_/B
+ sky130_fd_sc_hd__and4_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10279_ _10387_/A _10387_/B vssd1 vssd1 vccd1 vccd1 _10388_/A sky130_fd_sc_hd__and2_1
X_12018_ _12374_/A _12018_/B vssd1 vssd1 vccd1 vccd1 _12018_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_66_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16826_ _16880_/A _16758_/B _16695_/B _16604_/B vssd1 vssd1 vccd1 vccd1 _16828_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_19_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_988 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16757_ _16758_/A _15551_/Y _16758_/C vssd1 vssd1 vccd1 vccd1 _16759_/A sky130_fd_sc_hd__a21oi_1
XFILLER_19_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13969_ _13969_/A _13969_/B vssd1 vssd1 vccd1 vccd1 _13971_/B sky130_fd_sc_hd__xnor2_1
XFILLER_47_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15708_ _15707_/A _15707_/B _15707_/C vssd1 vssd1 vccd1 vccd1 _15708_/X sky130_fd_sc_hd__a21o_1
XFILLER_94_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16688_ _16688_/A _16688_/B vssd1 vssd1 vccd1 vccd1 _16690_/B sky130_fd_sc_hd__xor2_1
XFILLER_22_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15639_ _16315_/D _15639_/B vssd1 vssd1 vccd1 vccd1 _16499_/B sky130_fd_sc_hd__or2_4
XFILLER_34_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09160_ _10180_/A _11815_/B _14948_/B vssd1 vssd1 vccd1 vccd1 _09164_/A sky130_fd_sc_hd__and3_1
XFILLER_9_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17309_ input64/X _17321_/B _17321_/C vssd1 vssd1 vccd1 vccd1 _17309_/X sky130_fd_sc_hd__or3_1
X_09091_ _09091_/A _09091_/B _09318_/A vssd1 vssd1 vccd1 vccd1 _09092_/A sky130_fd_sc_hd__and3_1
XFILLER_119_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_802 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_898 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09993_ _09986_/A _09988_/B _09986_/B vssd1 vssd1 vccd1 vccd1 _09996_/A sky130_fd_sc_hd__o21ba_1
XFILLER_88_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08944_ _08945_/A _08945_/B vssd1 vssd1 vccd1 vccd1 _08944_/X sky130_fd_sc_hd__and2b_1
XFILLER_130_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08875_ _08832_/A _08832_/C _08832_/B vssd1 vssd1 vccd1 vccd1 _08875_/X sky130_fd_sc_hd__o21a_1
XFILLER_97_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_359 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09427_ _17119_/B _16933_/A vssd1 vssd1 vccd1 vccd1 _09427_/Y sky130_fd_sc_hd__nor2_1
XFILLER_40_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09358_ _09358_/A _09358_/B vssd1 vssd1 vccd1 vccd1 _09366_/C sky130_fd_sc_hd__or2_1
XFILLER_60_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09289_ _09289_/A _09289_/B vssd1 vssd1 vccd1 vccd1 _09291_/B sky130_fd_sc_hd__xnor2_1
XFILLER_5_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11320_ _11320_/A _11320_/B _11320_/C vssd1 vssd1 vccd1 vccd1 _11331_/B sky130_fd_sc_hd__or3_2
XFILLER_153_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11251_ _11347_/A _11347_/B vssd1 vssd1 vccd1 vccd1 _11348_/A sky130_fd_sc_hd__or2_1
XFILLER_4_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10202_ _10202_/A _10202_/B vssd1 vssd1 vccd1 vccd1 _10203_/C sky130_fd_sc_hd__xnor2_1
XFILLER_109_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11182_ _11182_/A _11182_/B _11182_/C vssd1 vssd1 vccd1 vccd1 _11182_/Y sky130_fd_sc_hd__nor3_1
XFILLER_133_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10133_ _10133_/A _10133_/B _10133_/C vssd1 vssd1 vccd1 vccd1 _10134_/C sky130_fd_sc_hd__nand3_1
XFILLER_133_194 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15990_ _16096_/B _15990_/B vssd1 vssd1 vccd1 vccd1 _15990_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_782 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10064_ _10064_/A _10064_/B vssd1 vssd1 vccd1 vccd1 _10066_/B sky130_fd_sc_hd__nor2_1
X_14941_ _12054_/A _15373_/B _10062_/B vssd1 vssd1 vccd1 vccd1 _14941_/X sky130_fd_sc_hd__a21o_1
XFILLER_75_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14872_ _14872_/A _14933_/B vssd1 vssd1 vccd1 vccd1 _16977_/A sky130_fd_sc_hd__or2_4
X_16611_ _16612_/B _16611_/B vssd1 vssd1 vccd1 vccd1 _16697_/B sky130_fd_sc_hd__and2b_1
XFILLER_85_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13823_ _13823_/A _13823_/B vssd1 vssd1 vccd1 vccd1 _13827_/A sky130_fd_sc_hd__xor2_2
X_17591_ fanout935/X _17591_/D vssd1 vssd1 vccd1 vccd1 _17591_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16542_ _16542_/A _16542_/B vssd1 vssd1 vccd1 vccd1 _16543_/B sky130_fd_sc_hd__nor2_1
XFILLER_141_82 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13754_ _13754_/A _13754_/B vssd1 vssd1 vccd1 vccd1 _13756_/B sky130_fd_sc_hd__xnor2_1
XFILLER_90_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10966_ _10966_/A _10966_/B vssd1 vssd1 vccd1 vccd1 _10969_/A sky130_fd_sc_hd__xnor2_1
X_12705_ _12044_/Y _12046_/Y _12049_/Y _12051_/Y _12383_/S _12865_/S vssd1 vssd1 vccd1
+ vccd1 _12705_/X sky130_fd_sc_hd__mux4_1
X_16473_ _16563_/A _16384_/Y _16472_/X vssd1 vssd1 vccd1 vccd1 _16475_/A sky130_fd_sc_hd__a21oi_1
XFILLER_43_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13685_ _13686_/A _13686_/B vssd1 vssd1 vccd1 vccd1 _13787_/A sky130_fd_sc_hd__or2_1
XFILLER_31_524 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10897_ _10991_/A _10897_/B _10897_/C vssd1 vssd1 vccd1 vccd1 _10995_/A sky130_fd_sc_hd__and3_1
XFILLER_31_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15424_ _15424_/A _15424_/B vssd1 vssd1 vccd1 vccd1 _15426_/B sky130_fd_sc_hd__xor2_1
XFILLER_31_568 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12636_ _12787_/B _12787_/D _12637_/D _12487_/A vssd1 vssd1 vccd1 vccd1 _12640_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_141_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15355_ _15355_/A _15355_/B vssd1 vssd1 vccd1 vccd1 _15356_/B sky130_fd_sc_hd__or2_1
XFILLER_15_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12567_ _13028_/A _13464_/B vssd1 vssd1 vccd1 vccd1 _12568_/B sky130_fd_sc_hd__nand2_1
XFILLER_156_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14306_ _14306_/A _14306_/B vssd1 vssd1 vccd1 vccd1 _14309_/A sky130_fd_sc_hd__xnor2_1
XFILLER_172_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11518_ _11518_/A _11518_/B _11518_/C _11563_/D vssd1 vssd1 vccd1 vccd1 _11521_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_171_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15286_ _15287_/A _15287_/B vssd1 vssd1 vccd1 vccd1 _15286_/Y sky130_fd_sc_hd__nor2_1
XFILLER_116_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12498_ _12498_/A _12498_/B _12498_/C vssd1 vssd1 vccd1 vccd1 _12499_/B sky130_fd_sc_hd__and3_1
XFILLER_116_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17025_ _16972_/A _16972_/B _10583_/A vssd1 vssd1 vccd1 vccd1 _17025_/Y sky130_fd_sc_hd__a21boi_1
X_14237_ _14237_/A _14237_/B _14236_/X vssd1 vssd1 vccd1 vccd1 _14239_/A sky130_fd_sc_hd__nor3b_1
X_11449_ _11453_/B _11449_/B _11449_/C vssd1 vssd1 vccd1 vccd1 _11495_/A sky130_fd_sc_hd__and3_1
XFILLER_109_191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14168_ _14387_/A _14433_/B vssd1 vssd1 vccd1 vccd1 _14170_/C sky130_fd_sc_hd__nand2_1
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13119_ _13120_/B _13120_/A vssd1 vssd1 vccd1 vccd1 _13119_/Y sky130_fd_sc_hd__nand2b_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14099_ _14188_/B _14101_/B vssd1 vssd1 vccd1 vccd1 _14194_/A sky130_fd_sc_hd__nand2_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1044 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16809_ _16809_/A _16809_/B _16809_/C vssd1 vssd1 vccd1 vccd1 _16809_/X sky130_fd_sc_hd__and3_1
XFILLER_121_19 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09212_ _09212_/A _09212_/B vssd1 vssd1 vccd1 vccd1 _09213_/B sky130_fd_sc_hd__nor2_1
X_09143_ _09143_/A _09231_/A vssd1 vssd1 vccd1 vccd1 _09145_/C sky130_fd_sc_hd__nor2_1
XFILLER_148_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09074_ _09074_/A _09074_/B vssd1 vssd1 vccd1 vccd1 _09076_/C sky130_fd_sc_hd__nand2_1
XFILLER_162_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09976_ _09976_/A _09976_/B vssd1 vssd1 vccd1 vccd1 _10004_/A sky130_fd_sc_hd__xnor2_1
XFILLER_104_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08927_ _08927_/A _09012_/B vssd1 vssd1 vccd1 vccd1 _08930_/B sky130_fd_sc_hd__nand2_1
XFILLER_130_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08858_ _17385_/A _17383_/A _11900_/D _09321_/D vssd1 vssd1 vccd1 vccd1 _08859_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_17_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08789_ _08791_/B _09319_/D _09058_/C _08791_/A vssd1 vssd1 vccd1 vccd1 _08792_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_55_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10820_ _11095_/B _17468_/D _17467_/D _11095_/A vssd1 vssd1 vccd1 vccd1 _10820_/Y
+ sky130_fd_sc_hd__a22oi_1
XTAP_2947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10751_ _10993_/C _12054_/B _10660_/A _10658_/Y vssd1 vssd1 vccd1 vccd1 _10757_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_40_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13470_ _14155_/A _13966_/D vssd1 vssd1 vccd1 vccd1 _13471_/B sky130_fd_sc_hd__nand2_1
XFILLER_40_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10682_ _10690_/A _10690_/B vssd1 vssd1 vccd1 vccd1 _10682_/Y sky130_fd_sc_hd__nor2_1
XFILLER_139_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12421_ _12421_/A _12421_/B _12421_/C vssd1 vssd1 vccd1 vccd1 _12434_/B sky130_fd_sc_hd__nand3_1
XFILLER_40_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15140_ _15270_/A _15270_/B vssd1 vssd1 vccd1 vccd1 _15140_/Y sky130_fd_sc_hd__nor2_1
X_12352_ _12351_/A _12351_/B _12350_/X vssd1 vssd1 vccd1 vccd1 _12353_/B sky130_fd_sc_hd__o21bai_1
XFILLER_166_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11303_ _11423_/B fanout874/X _11261_/A _11259_/Y vssd1 vssd1 vccd1 vccd1 _11304_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_154_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15071_ _15071_/A _15071_/B vssd1 vssd1 vccd1 vccd1 _15071_/Y sky130_fd_sc_hd__nor2_1
X_12283_ _12283_/A _12283_/B vssd1 vssd1 vccd1 vccd1 _12284_/B sky130_fd_sc_hd__nor2_1
XFILLER_135_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14022_ _14113_/B _14022_/B vssd1 vssd1 vccd1 vccd1 _14025_/A sky130_fd_sc_hd__nand2_1
XFILLER_107_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11234_ _11234_/A _11234_/B vssd1 vssd1 vccd1 vccd1 _11711_/A sky130_fd_sc_hd__or2_1
XFILLER_135_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_963 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11165_ _11165_/A _11165_/B _11165_/C vssd1 vssd1 vccd1 vccd1 _11204_/A sky130_fd_sc_hd__or3_1
XFILLER_95_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10116_ _10116_/A _10116_/B vssd1 vssd1 vccd1 vccd1 _10118_/A sky130_fd_sc_hd__nor2_1
X_11096_ _11095_/B _11240_/C _11095_/D _11095_/A vssd1 vssd1 vccd1 vccd1 _11096_/Y
+ sky130_fd_sc_hd__a22oi_1
X_15973_ _16080_/B _15973_/B vssd1 vssd1 vccd1 vccd1 _15976_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_443 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10047_ _10162_/A _10170_/A _10162_/C vssd1 vssd1 vccd1 vccd1 _10163_/A sky130_fd_sc_hd__o21ai_1
X_14924_ _14924_/A _14929_/A _14924_/C vssd1 vssd1 vccd1 vccd1 _14962_/B sky130_fd_sc_hd__or3_2
XFILLER_64_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14855_ _15811_/A _15709_/A _15709_/B vssd1 vssd1 vccd1 vccd1 _15898_/B sky130_fd_sc_hd__and3_1
XFILLER_17_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13806_ _13915_/B _13806_/B vssd1 vssd1 vccd1 vccd1 _13809_/A sky130_fd_sc_hd__or2_1
X_17574_ fanout936/X _17574_/D vssd1 vssd1 vccd1 vccd1 _17574_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14786_ _14786_/A _14851_/A vssd1 vssd1 vccd1 vccd1 _14805_/B sky130_fd_sc_hd__or2_1
X_11998_ _11998_/A _11998_/B _12197_/B _11998_/D vssd1 vssd1 vccd1 vccd1 _11998_/X
+ sky130_fd_sc_hd__or4_1
X_16525_ _16616_/B _16525_/B vssd1 vssd1 vccd1 vccd1 _16527_/C sky130_fd_sc_hd__nor2_1
XFILLER_32_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13737_ _13846_/A _13738_/B vssd1 vssd1 vccd1 vccd1 _13739_/B sky130_fd_sc_hd__nand2_1
X_10949_ _10946_/X _10947_/Y _10927_/X _11059_/A vssd1 vssd1 vccd1 vccd1 _10949_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_16_384 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16456_ _16457_/B _16457_/A vssd1 vssd1 vccd1 vccd1 _16456_/Y sky130_fd_sc_hd__nand2b_1
X_13668_ _13668_/A _13668_/B vssd1 vssd1 vccd1 vccd1 _13669_/B sky130_fd_sc_hd__and2_1
X_15407_ _15408_/A _15408_/B _15408_/C vssd1 vssd1 vccd1 vccd1 _15501_/A sky130_fd_sc_hd__o21a_1
X_12619_ _12619_/A _12619_/B vssd1 vssd1 vccd1 vccd1 _12621_/A sky130_fd_sc_hd__nor2_1
X_16387_ _16387_/A _16387_/B _16387_/C vssd1 vssd1 vccd1 vccd1 _16389_/B sky130_fd_sc_hd__or3_1
X_13599_ _13600_/A _13600_/B vssd1 vssd1 vccd1 vccd1 _13601_/A sky130_fd_sc_hd__nor2_1
XFILLER_145_702 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15338_ _16935_/A _15147_/A _15393_/B vssd1 vssd1 vccd1 vccd1 _15338_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_144_223 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15269_ _16935_/A _15204_/B _15147_/A vssd1 vssd1 vccd1 vccd1 _15270_/C sky130_fd_sc_hd__o21a_1
XFILLER_6_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17008_ _17008_/A _17012_/B vssd1 vssd1 vccd1 vccd1 _17009_/B sky130_fd_sc_hd__or2_1
XFILLER_132_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout507 _12592_/A vssd1 vssd1 vccd1 vccd1 _09892_/A sky130_fd_sc_hd__buf_4
X_09830_ _09769_/B _09776_/B _09769_/D _09769_/A vssd1 vssd1 vccd1 vccd1 _09830_/X
+ sky130_fd_sc_hd__a22o_1
Xfanout518 _17517_/Q vssd1 vssd1 vccd1 vccd1 _15373_/C sky130_fd_sc_hd__clkbuf_4
Xfanout529 _10970_/A vssd1 vssd1 vccd1 vccd1 _11117_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_98_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09761_ _09761_/A vssd1 vssd1 vccd1 vccd1 _09765_/A sky130_fd_sc_hd__inv_2
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09692_ _10236_/A _10236_/B _09985_/D _09979_/C vssd1 vssd1 vccd1 vccd1 _09695_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_132_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_722 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_254 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_927 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09126_ _09128_/D vssd1 vssd1 vccd1 vccd1 _09126_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_136_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09057_ _09057_/A _09057_/B vssd1 vssd1 vccd1 vccd1 _09063_/A sky130_fd_sc_hd__nor2_1
XFILLER_135_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09959_ _09960_/A _09960_/B _09960_/C vssd1 vssd1 vccd1 vccd1 _09959_/X sky130_fd_sc_hd__and3_1
XFILLER_106_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12970_ _12971_/B _12971_/A vssd1 vssd1 vccd1 vccd1 _13107_/B sky130_fd_sc_hd__and2b_1
XFILLER_46_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11921_ _11921_/A _12179_/A vssd1 vssd1 vccd1 vccd1 _11924_/A sky130_fd_sc_hd__or2_1
XFILLER_57_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_947 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14640_ _14738_/A _14641_/C vssd1 vssd1 vccd1 vccd1 _14675_/A sky130_fd_sc_hd__nand2_1
XTAP_3489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11852_ _12700_/B _11852_/B vssd1 vssd1 vccd1 vccd1 _11854_/C sky130_fd_sc_hd__or2_1
XTAP_2755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10803_ _10803_/A _10803_/B vssd1 vssd1 vccd1 vccd1 _10816_/A sky130_fd_sc_hd__xnor2_1
XTAP_2777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14571_ _14621_/A _14570_/C _14570_/A vssd1 vssd1 vccd1 vccd1 _14571_/X sky130_fd_sc_hd__a21o_1
XTAP_2799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11783_ _14872_/A _14924_/C vssd1 vssd1 vccd1 vccd1 _11783_/Y sky130_fd_sc_hd__nor2_1
XFILLER_25_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16310_ _16310_/A _16310_/B _16310_/C _16310_/D vssd1 vssd1 vccd1 vccd1 _16310_/X
+ sky130_fd_sc_hd__and4_1
X_13522_ _13632_/A _13735_/B _13735_/D _13522_/D vssd1 vssd1 vccd1 vccd1 _13637_/A
+ sky130_fd_sc_hd__nand4_1
X_10734_ _10662_/X _10732_/Y _10728_/B _10714_/X vssd1 vssd1 vccd1 vccd1 _10734_/X
+ sky130_fd_sc_hd__o211a_1
X_17290_ _17464_/Q _17290_/A2 _17288_/X _17289_/X _17293_/C1 vssd1 vssd1 vccd1 vccd1
+ _17464_/D sky130_fd_sc_hd__o221a_1
XFILLER_14_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16241_ _16241_/A _16241_/B _16239_/Y vssd1 vssd1 vccd1 vccd1 _16242_/B sky130_fd_sc_hd__or3b_1
X_13453_ _13897_/A _13564_/C _13453_/C vssd1 vssd1 vccd1 vccd1 _13569_/B sky130_fd_sc_hd__and3_1
XFILLER_51_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10665_ _10670_/B _10665_/B vssd1 vssd1 vccd1 vccd1 _10667_/B sky130_fd_sc_hd__nand2_1
XFILLER_127_702 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12404_ _12869_/A _13334_/C _13208_/D _12714_/A vssd1 vssd1 vccd1 vccd1 _12406_/A
+ sky130_fd_sc_hd__a22oi_1
X_16172_ _16172_/A _16172_/B vssd1 vssd1 vccd1 vccd1 _16174_/A sky130_fd_sc_hd__xor2_1
XFILLER_12_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13384_ _13261_/A _13263_/A _13504_/B _13382_/X vssd1 vssd1 vccd1 vccd1 _13385_/B
+ sky130_fd_sc_hd__a211oi_1
X_10596_ _10709_/A _10709_/B vssd1 vssd1 vccd1 vccd1 _10599_/A sky130_fd_sc_hd__or2_1
XFILLER_166_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15123_ _15126_/B vssd1 vssd1 vccd1 vccd1 _15123_/Y sky130_fd_sc_hd__inv_2
X_12335_ _17405_/A _12334_/B _12334_/C vssd1 vssd1 vccd1 vccd1 _12336_/B sky130_fd_sc_hd__a21oi_1
XFILLER_31_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15054_ _16207_/B _15053_/X _15051_/X _15049_/X vssd1 vssd1 vccd1 vccd1 _15054_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_114_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12266_ _12266_/A _12437_/B vssd1 vssd1 vccd1 vccd1 _12268_/C sky130_fd_sc_hd__nand2_1
XFILLER_107_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14005_ _13904_/A _13904_/B _13902_/B vssd1 vssd1 vccd1 vccd1 _14007_/B sky130_fd_sc_hd__o21ai_1
X_11217_ _11217_/A _11217_/B vssd1 vssd1 vccd1 vccd1 _11220_/A sky130_fd_sc_hd__xnor2_1
XFILLER_123_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12197_ _12197_/A _12197_/B vssd1 vssd1 vccd1 vccd1 _12198_/C sky130_fd_sc_hd__nor2_1
XFILLER_123_985 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput81 _17474_/Q vssd1 vssd1 vccd1 vccd1 leds[8] sky130_fd_sc_hd__clkbuf_1
XFILLER_68_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput92 _17451_/Q vssd1 vssd1 vccd1 vccd1 o_wb_data[17] sky130_fd_sc_hd__clkbuf_1
X_11148_ _11148_/A _11148_/B vssd1 vssd1 vccd1 vccd1 _11149_/B sky130_fd_sc_hd__nand2_1
XFILLER_96_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11079_ _11077_/A _11077_/C _11110_/A vssd1 vssd1 vccd1 vccd1 _11080_/D sky130_fd_sc_hd__o21ai_1
X_15956_ _16446_/A _16814_/A vssd1 vssd1 vccd1 vccd1 _16062_/C sky130_fd_sc_hd__nor2_1
XFILLER_110_679 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14907_ _14899_/C _14906_/X _14905_/X _14903_/X vssd1 vssd1 vccd1 vccd1 _15553_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_37_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15887_ _15884_/Y _15885_/Y _15886_/Y vssd1 vssd1 vccd1 vccd1 _15887_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_48_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14838_ _12016_/B _11781_/B _14837_/Y vssd1 vssd1 vccd1 vccd1 _14838_/X sky130_fd_sc_hd__o21a_1
XFILLER_51_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14769_ _14769_/A _14865_/B vssd1 vssd1 vccd1 vccd1 _16918_/B sky130_fd_sc_hd__or2_1
X_17557_ fanout951/X _17557_/D vssd1 vssd1 vccd1 vccd1 _17557_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16508_ _16509_/A _16509_/B _16509_/C vssd1 vssd1 vccd1 vccd1 _16616_/A sky130_fd_sc_hd__a21oi_1
XFILLER_60_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17488_ fanout942/X _17488_/D vssd1 vssd1 vccd1 vccd1 _17488_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16439_ _16439_/A _16439_/B vssd1 vssd1 vccd1 vccd1 _16442_/A sky130_fd_sc_hd__xor2_1
XFILLER_20_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout304 _08720_/Y vssd1 vssd1 vccd1 vccd1 _15116_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_59_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout315 _17611_/Q vssd1 vssd1 vccd1 vccd1 _15071_/A sky130_fd_sc_hd__clkbuf_2
Xfanout326 _17541_/Q vssd1 vssd1 vccd1 vccd1 _12770_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_141_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout337 _17100_/C vssd1 vssd1 vccd1 vccd1 _14676_/A sky130_fd_sc_hd__clkbuf_4
X_09813_ _09813_/A _09813_/B _09813_/C vssd1 vssd1 vccd1 vccd1 _09813_/X sky130_fd_sc_hd__and3_1
Xfanout348 _09360_/A vssd1 vssd1 vccd1 vccd1 _12804_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_101_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout359 _16965_/C vssd1 vssd1 vccd1 vccd1 _14554_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_98_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09744_ _09724_/X _09740_/B _09743_/Y _09621_/X vssd1 vssd1 vccd1 vccd1 _09776_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_28_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09675_ _09678_/B _09675_/B _09675_/C vssd1 vssd1 vccd1 vccd1 _09681_/A sky130_fd_sc_hd__nor3_1
XFILLER_67_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10450_ _10450_/A _10450_/B vssd1 vssd1 vccd1 vccd1 _10451_/B sky130_fd_sc_hd__nor2_1
XFILLER_108_223 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09109_ _09110_/A _09110_/B vssd1 vssd1 vccd1 vccd1 _09153_/B sky130_fd_sc_hd__and2_1
XFILLER_109_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10381_ _10382_/B _10382_/A vssd1 vssd1 vccd1 vccd1 _10390_/B sky130_fd_sc_hd__nand2b_1
X_12120_ _12309_/A _12118_/Y _11905_/X _11909_/A vssd1 vssd1 vccd1 vccd1 _12122_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_105_930 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12051_ _14911_/B _12051_/B vssd1 vssd1 vccd1 vccd1 _12051_/Y sky130_fd_sc_hd__nand2_1
XFILLER_151_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11002_ _10999_/X _11000_/Y _10977_/X _11051_/A vssd1 vssd1 vccd1 vccd1 _11002_/Y
+ sky130_fd_sc_hd__o211ai_1
XFILLER_2_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout860 _10359_/B vssd1 vssd1 vccd1 vccd1 _11117_/D sky130_fd_sc_hd__buf_2
Xfanout871 _10479_/B vssd1 vssd1 vccd1 vccd1 _11115_/C sky130_fd_sc_hd__buf_2
XFILLER_120_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15810_ _14924_/A _15457_/B _13390_/X _15804_/Y _15809_/Y vssd1 vssd1 vccd1 vccd1
+ _15810_/X sky130_fd_sc_hd__o311a_1
Xfanout882 _10805_/D vssd1 vssd1 vccd1 vccd1 _17469_/D sky130_fd_sc_hd__buf_2
X_16790_ _13689_/A _16789_/Y _16788_/Y vssd1 vssd1 vccd1 vccd1 _16792_/A sky130_fd_sc_hd__a21oi_1
Xfanout893 _17480_/Q vssd1 vssd1 vccd1 vccd1 _17468_/D sky130_fd_sc_hd__buf_2
XFILLER_19_914 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15741_ _15741_/A _15741_/B vssd1 vssd1 vccd1 vccd1 _15743_/B sky130_fd_sc_hd__xnor2_2
XFILLER_46_722 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12953_ _12795_/A _13080_/C _12796_/A _12794_/B vssd1 vssd1 vccd1 vccd1 _12954_/B
+ sky130_fd_sc_hd__a31o_1
XTAP_3231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11904_ _08859_/A _08861_/B _08859_/B vssd1 vssd1 vccd1 vccd1 _11906_/B sky130_fd_sc_hd__o21ba_1
XTAP_3264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15672_ _15673_/A _15673_/B vssd1 vssd1 vccd1 vccd1 _15764_/B sky130_fd_sc_hd__nand2_1
XFILLER_18_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12884_ _12884_/A _12884_/B vssd1 vssd1 vccd1 vccd1 _12886_/C sky130_fd_sc_hd__xnor2_1
XFILLER_33_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17411_ _17411_/A _17425_/B vssd1 vssd1 vccd1 vccd1 _17411_/X sky130_fd_sc_hd__or2_1
X_14623_ _14624_/A _14624_/B vssd1 vssd1 vccd1 vccd1 _14660_/B sky130_fd_sc_hd__nor2_1
XTAP_2563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11835_ _11837_/A _11835_/B vssd1 vssd1 vccd1 vccd1 _11835_/Y sky130_fd_sc_hd__nand2_1
XTAP_2574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17342_ _09321_/D _17356_/A2 _17341_/X _17406_/C1 vssd1 vssd1 vccd1 vccd1 _17500_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14554_ _14554_/A _14738_/B vssd1 vssd1 vccd1 vccd1 _14555_/B sky130_fd_sc_hd__nand2_1
XTAP_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11766_ _16866_/A _16866_/B vssd1 vssd1 vccd1 vccd1 _11766_/X sky130_fd_sc_hd__or2_1
XFILLER_42_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13505_ _13506_/A _13506_/B vssd1 vssd1 vccd1 vccd1 _13619_/A sky130_fd_sc_hd__nand2_1
X_10717_ _11095_/A _11095_/B _10962_/B _14849_/A vssd1 vssd1 vccd1 vccd1 _10720_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_147_808 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17273_ _17600_/Q _17273_/A2 _17273_/B1 vssd1 vssd1 vccd1 vccd1 _17273_/X sky130_fd_sc_hd__a21o_1
XFILLER_9_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14485_ _14641_/A _14641_/B _14545_/D _14485_/D vssd1 vssd1 vccd1 vccd1 _14557_/A
+ sky130_fd_sc_hd__and4_1
X_11697_ _15614_/A _15614_/B vssd1 vssd1 vccd1 vccd1 _15615_/A sky130_fd_sc_hd__nor2_1
X_16224_ _16224_/A vssd1 vssd1 vccd1 vccd1 _17559_/D sky130_fd_sc_hd__inv_2
X_13436_ _14215_/A _13664_/D vssd1 vssd1 vccd1 vccd1 _13438_/B sky130_fd_sc_hd__nand2_1
XFILLER_174_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10648_ _10648_/A _10742_/A vssd1 vssd1 vccd1 vccd1 _10735_/A sky130_fd_sc_hd__or2_1
XFILLER_9_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_532 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16155_ _16155_/A _16155_/B vssd1 vssd1 vccd1 vccd1 _16157_/B sky130_fd_sc_hd__xnor2_1
X_13367_ _13368_/A _13368_/B vssd1 vssd1 vccd1 vccd1 _13369_/B sky130_fd_sc_hd__nand2_1
XFILLER_155_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10579_ _10579_/A _10579_/B vssd1 vssd1 vccd1 vccd1 _10582_/B sky130_fd_sc_hd__nor2_1
XFILLER_170_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15106_ _15106_/A _15106_/B vssd1 vssd1 vccd1 vccd1 _15106_/Y sky130_fd_sc_hd__nand2_1
XFILLER_115_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12318_ _12150_/A _12149_/B _12149_/A vssd1 vssd1 vccd1 vccd1 _12355_/A sky130_fd_sc_hd__o21ba_1
X_16086_ _16086_/A _16355_/B _16086_/C vssd1 vssd1 vccd1 vccd1 _16197_/B sky130_fd_sc_hd__and3_1
X_13298_ _13414_/B _13844_/C vssd1 vssd1 vccd1 vccd1 _13657_/B sky130_fd_sc_hd__nand2_1
XFILLER_138_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15037_ _15097_/A _15037_/B vssd1 vssd1 vccd1 vccd1 _15037_/X sky130_fd_sc_hd__or2_1
X_12249_ _12250_/A _12250_/B vssd1 vssd1 vccd1 vccd1 _12421_/B sky130_fd_sc_hd__nand2b_1
XFILLER_123_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_847 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16988_ _16989_/A _16989_/B vssd1 vssd1 vccd1 vccd1 _17049_/A sky130_fd_sc_hd__nor2_1
X_15939_ _15939_/A _15939_/B vssd1 vssd1 vccd1 vccd1 _15940_/B sky130_fd_sc_hd__nor2_1
XFILLER_36_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09460_ _09440_/X _09455_/B _09459_/Y _09335_/A vssd1 vssd1 vccd1 vccd1 _09460_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_64_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17609_ fanout950/X _17609_/D vssd1 vssd1 vccd1 vccd1 _17609_/Q sky130_fd_sc_hd__dfxtp_2
X_09391_ _09391_/A _09391_/B _09391_/C vssd1 vssd1 vccd1 vccd1 _09393_/D sky130_fd_sc_hd__and3_1
XFILLER_91_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_830 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout123 _17244_/B vssd1 vssd1 vccd1 vccd1 _17274_/B sky130_fd_sc_hd__buf_2
Xfanout134 _15755_/B vssd1 vssd1 vccd1 vccd1 _16497_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_87_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout145 _16165_/A vssd1 vssd1 vccd1 vccd1 _15278_/A sky130_fd_sc_hd__clkbuf_2
Xfanout156 _17426_/A2 vssd1 vssd1 vccd1 vccd1 _17422_/A2 sky130_fd_sc_hd__buf_2
Xfanout167 _16595_/B vssd1 vssd1 vccd1 vccd1 _16938_/D sky130_fd_sc_hd__buf_2
Xfanout178 _15552_/X vssd1 vssd1 vccd1 vccd1 _16514_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_102_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout189 _15263_/Y vssd1 vssd1 vccd1 vccd1 _16352_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_102_999 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09727_ _09727_/A _09727_/B vssd1 vssd1 vccd1 vccd1 _09733_/A sky130_fd_sc_hd__nor2_1
XFILLER_28_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09658_ _09658_/A _09658_/B vssd1 vssd1 vccd1 vccd1 _09788_/B sky130_fd_sc_hd__or2_1
XFILLER_15_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09589_ _09589_/A _09589_/B vssd1 vssd1 vccd1 vccd1 _09722_/A sky130_fd_sc_hd__xnor2_1
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11620_ _11620_/A _11624_/A _11620_/C vssd1 vssd1 vccd1 vccd1 _11622_/A sky130_fd_sc_hd__nor3_1
XFILLER_24_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11551_ _11538_/A _11537_/C _11537_/B vssd1 vssd1 vccd1 vccd1 _11551_/X sky130_fd_sc_hd__o21a_1
XFILLER_168_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10502_ _10503_/A _10503_/B _10503_/C vssd1 vssd1 vccd1 vccd1 _10502_/X sky130_fd_sc_hd__a21o_1
X_14270_ _14270_/A _14270_/B _14270_/C vssd1 vssd1 vccd1 vccd1 _14271_/B sky130_fd_sc_hd__and3_1
X_11482_ _11484_/B _11481_/Y _11520_/C _11518_/C vssd1 vssd1 vccd1 vccd1 _11522_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_7_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13221_ _13221_/A _13221_/B vssd1 vssd1 vccd1 vccd1 _13223_/B sky130_fd_sc_hd__nand2_1
XFILLER_137_863 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10433_ _10434_/A _10432_/Y _10545_/C _10543_/B vssd1 vssd1 vccd1 vccd1 _10547_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_94 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13152_ _13019_/A _13021_/B _13019_/B vssd1 vssd1 vccd1 vccd1 _13154_/B sky130_fd_sc_hd__o21ba_1
X_10364_ _10364_/A _10364_/B vssd1 vssd1 vccd1 vccd1 _10484_/A sky130_fd_sc_hd__xor2_1
XFILLER_163_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12103_ _12103_/A _12103_/B vssd1 vssd1 vccd1 vccd1 _12105_/A sky130_fd_sc_hd__nor2_1
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13083_ _13083_/A _13213_/A _13083_/C vssd1 vssd1 vccd1 vccd1 _13213_/B sky130_fd_sc_hd__nor3_1
X_10295_ _10296_/A _10296_/C vssd1 vssd1 vccd1 vccd1 _10301_/B sky130_fd_sc_hd__nor2_1
XFILLER_105_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16911_ _16911_/A _16911_/B vssd1 vssd1 vccd1 vccd1 _16911_/Y sky130_fd_sc_hd__nand2_2
X_12034_ _12031_/Y _12033_/Y _14948_/A vssd1 vssd1 vccd1 vccd1 _12034_/X sky130_fd_sc_hd__mux2_1
XFILLER_105_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16842_ _16843_/A _16843_/B vssd1 vssd1 vccd1 vccd1 _16906_/B sky130_fd_sc_hd__nand2_1
XFILLER_144_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout690 _17501_/Q vssd1 vssd1 vccd1 vccd1 fanout690/X sky130_fd_sc_hd__buf_6
XFILLER_92_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16773_ _16774_/A _16774_/B vssd1 vssd1 vccd1 vccd1 _16843_/A sky130_fd_sc_hd__and2b_1
X_13985_ _13985_/A _13985_/B vssd1 vssd1 vccd1 vccd1 _13988_/A sky130_fd_sc_hd__xor2_1
XFILLER_18_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15724_ _16136_/A _17083_/A vssd1 vssd1 vccd1 vccd1 _15724_/X sky130_fd_sc_hd__and2_1
X_12936_ _12938_/A _12938_/B _12938_/C vssd1 vssd1 vccd1 vccd1 _12985_/A sky130_fd_sc_hd__a21oi_2
XFILLER_19_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_522 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12867_ _14356_/S _12864_/Y _12866_/Y _13831_/S _15457_/A vssd1 vssd1 vccd1 vccd1
+ _12867_/X sky130_fd_sc_hd__a221o_1
XTAP_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15655_ _15655_/A _15655_/B _15656_/B vssd1 vssd1 vccd1 vccd1 _15769_/A sky130_fd_sc_hd__and3_1
XTAP_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11818_ _12848_/S _11818_/B vssd1 vssd1 vccd1 vccd1 _11818_/Y sky130_fd_sc_hd__nor2_1
X_14606_ _14606_/A _14606_/B vssd1 vssd1 vccd1 vccd1 _14609_/A sky130_fd_sc_hd__xor2_1
XFILLER_33_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15586_ _15685_/B _15587_/B vssd1 vssd1 vccd1 vccd1 _15686_/A sky130_fd_sc_hd__and2b_1
XFILLER_144_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12798_ _12798_/A _12798_/B _12798_/C vssd1 vssd1 vccd1 vccd1 _12799_/B sky130_fd_sc_hd__and3_1
XTAP_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17325_ input41/X _17359_/B _17359_/C vssd1 vssd1 vccd1 vccd1 _17325_/X sky130_fd_sc_hd__or3_1
X_14537_ wire116/X _14281_/Y _14534_/Y _14535_/Y _14536_/X vssd1 vssd1 vccd1 vccd1
+ _14629_/B sky130_fd_sc_hd__o311ai_2
X_11749_ _11749_/A _11749_/B vssd1 vssd1 vccd1 vccd1 _11750_/B sky130_fd_sc_hd__xnor2_2
XFILLER_30_997 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14468_ _14469_/A _14469_/B vssd1 vssd1 vccd1 vccd1 _14531_/A sky130_fd_sc_hd__nor2_1
X_17256_ _17562_/Q _17292_/B vssd1 vssd1 vccd1 vccd1 _17256_/X sky130_fd_sc_hd__and2_1
XFILLER_105_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16207_ _16294_/B _16207_/B _16207_/C vssd1 vssd1 vccd1 vccd1 _16207_/X sky130_fd_sc_hd__or3_2
X_13419_ _13420_/A _13420_/B vssd1 vssd1 vccd1 vccd1 _13419_/Y sky130_fd_sc_hd__nand2b_1
X_17187_ input28/X _17362_/B _17429_/B vssd1 vssd1 vccd1 vccd1 _17187_/Y sky130_fd_sc_hd__nor3_4
X_14399_ _14466_/A _14400_/C _14400_/A vssd1 vssd1 vccd1 vccd1 _14399_/X sky130_fd_sc_hd__a21o_1
XFILLER_143_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16138_ _16138_/A _16499_/B vssd1 vssd1 vccd1 vccd1 _16140_/B sky130_fd_sc_hd__nor2_1
XFILLER_155_693 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16069_ _16070_/A _16070_/B vssd1 vssd1 vccd1 vccd1 _16069_/Y sky130_fd_sc_hd__nand2b_1
X_08960_ _09077_/A _09077_/B vssd1 vssd1 vccd1 vccd1 _08962_/C sky130_fd_sc_hd__nand2_1
XFILLER_142_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08891_ _08904_/B _08904_/C _08904_/A vssd1 vssd1 vccd1 vccd1 _08905_/A sky130_fd_sc_hd__a21o_1
XFILLER_97_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09512_ _09639_/C _09937_/B _09379_/A _09377_/Y vssd1 vssd1 vccd1 vccd1 _09513_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_71_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09443_ _09443_/A _09443_/B vssd1 vssd1 vccd1 vccd1 _09449_/A sky130_fd_sc_hd__nor2_1
XFILLER_64_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_544 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09374_ _09639_/C _09843_/D _09206_/A _09204_/Y vssd1 vssd1 vccd1 vccd1 _09375_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_21_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_1019 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10080_ _10080_/A _10080_/B vssd1 vssd1 vccd1 vccd1 _10081_/B sky130_fd_sc_hd__or2_1
XFILLER_99_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_763 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_796 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13770_ _13770_/A _13770_/B _13770_/C vssd1 vssd1 vccd1 vccd1 _13771_/B sky130_fd_sc_hd__or3_1
Xwb_buttons_leds_964 vssd1 vssd1 vccd1 vccd1 wb_buttons_leds_964/HI led_enb[6] sky130_fd_sc_hd__conb_1
X_10982_ _10745_/C _10532_/D _10746_/A _10744_/Y vssd1 vssd1 vccd1 vccd1 _10984_/C
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_62_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12721_ _12722_/B _13464_/B _13348_/B _12722_/A vssd1 vssd1 vccd1 vccd1 _12723_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_55_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_1014 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15440_ _15363_/A _15363_/B _15361_/Y vssd1 vssd1 vccd1 vccd1 _15442_/B sky130_fd_sc_hd__a21bo_1
X_12652_ _17405_/A _13080_/C vssd1 vssd1 vccd1 vccd1 _12654_/B sky130_fd_sc_hd__nand2_1
XFILLER_70_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11603_ _11603_/A _11603_/B _11603_/C vssd1 vssd1 vccd1 vccd1 _11610_/B sky130_fd_sc_hd__or3_1
X_15371_ _15303_/A _15370_/X _15998_/A _11691_/Y vssd1 vssd1 vccd1 vccd1 _15390_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_30_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12583_ _12583_/A _12583_/B vssd1 vssd1 vccd1 vccd1 _12585_/C sky130_fd_sc_hd__xnor2_1
XFILLER_30_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14322_ _14324_/A _14389_/B vssd1 vssd1 vccd1 vccd1 _14325_/A sky130_fd_sc_hd__nor2_1
X_17110_ _14867_/A _16974_/B _14929_/X _14827_/Y vssd1 vssd1 vccd1 vccd1 _17110_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_11534_ _11534_/A _11534_/B vssd1 vssd1 vccd1 vccd1 _11535_/B sky130_fd_sc_hd__nand2_1
XFILLER_156_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17041_ _16982_/A _17119_/B _17039_/X _17085_/A vssd1 vssd1 vccd1 vccd1 _17043_/C
+ sky130_fd_sc_hd__a211oi_1
XFILLER_7_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14253_ _14253_/A _14253_/B vssd1 vssd1 vccd1 vccd1 _14255_/A sky130_fd_sc_hd__nor2_1
XFILLER_171_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11465_ _11465_/A _11465_/B vssd1 vssd1 vccd1 vccd1 _15997_/A sky130_fd_sc_hd__xor2_1
XFILLER_125_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13204_ _13075_/A _13075_/Y _13201_/Y _13203_/A vssd1 vssd1 vccd1 vccd1 _13249_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_143_129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10416_ _15805_/A _10299_/D _10300_/A _10298_/Y vssd1 vssd1 vccd1 vccd1 _10418_/C
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_171_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14184_ _14185_/A _14273_/B _14184_/C vssd1 vssd1 vccd1 vccd1 _14186_/A sky130_fd_sc_hd__and3_1
X_11396_ _11396_/A _11396_/B _11396_/C vssd1 vssd1 vccd1 vccd1 _11396_/X sky130_fd_sc_hd__and3_1
XFILLER_124_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13135_ _13264_/B _13132_/X _12993_/X _12999_/A vssd1 vssd1 vccd1 vccd1 _13136_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_48_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10347_ _10349_/A _10349_/B vssd1 vssd1 vccd1 vccd1 _10347_/X sky130_fd_sc_hd__or2_1
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_931 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13066_ _14050_/B _13194_/D _13067_/D _14213_/A vssd1 vssd1 vccd1 vccd1 _13068_/A
+ sky130_fd_sc_hd__a22oi_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10278_ _10278_/A _10278_/B vssd1 vssd1 vccd1 vccd1 _10387_/B sky130_fd_sc_hd__nor2_1
XFILLER_2_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12017_ _11780_/Y _12377_/A _12015_/Y vssd1 vssd1 vccd1 vccd1 _12018_/B sky130_fd_sc_hd__o21ai_1
XFILLER_78_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16825_ _16938_/A _16935_/B _16746_/A _16744_/B vssd1 vssd1 vccd1 vccd1 _16829_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_65_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_861 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16756_ _16827_/A _16827_/C vssd1 vssd1 vccd1 vccd1 _16758_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13968_ _14215_/A _13968_/B vssd1 vssd1 vccd1 vccd1 _13969_/B sky130_fd_sc_hd__nand2_1
XFILLER_19_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_511 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_596 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15707_ _15707_/A _15707_/B _15707_/C vssd1 vssd1 vccd1 vccd1 _15707_/Y sky130_fd_sc_hd__nand3_1
X_12919_ _12919_/A _13065_/B vssd1 vssd1 vccd1 vccd1 _12920_/C sky130_fd_sc_hd__nand2_1
X_16687_ _16685_/X _16687_/B vssd1 vssd1 vccd1 vccd1 _16688_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13899_ _13790_/A _13792_/B _13790_/B vssd1 vssd1 vccd1 vccd1 _13900_/B sky130_fd_sc_hd__o21ba_1
X_15638_ _16315_/D _15639_/B vssd1 vssd1 vccd1 vccd1 _15638_/Y sky130_fd_sc_hd__nor2_1
XTAP_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15569_ _16262_/A _16410_/A vssd1 vssd1 vccd1 vccd1 _15570_/B sky130_fd_sc_hd__nor2_1
X_17308_ _12127_/C _17308_/A2 _17307_/X _17358_/C1 vssd1 vssd1 vccd1 vccd1 _17483_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_147_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09090_ _09091_/B _09318_/A _09091_/A vssd1 vssd1 vccd1 vccd1 _09093_/A sky130_fd_sc_hd__a21o_1
XFILLER_174_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17239_ _17447_/Q _17293_/A2 _17237_/X _17238_/X _17284_/C1 vssd1 vssd1 vccd1 vccd1
+ _17447_/D sky130_fd_sc_hd__o221a_1
XFILLER_174_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_990 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_814 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09992_ _10004_/B _10004_/C _10004_/A vssd1 vssd1 vccd1 vccd1 _10005_/A sky130_fd_sc_hd__a21o_1
XFILLER_103_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08943_ _08943_/A _08943_/B vssd1 vssd1 vccd1 vccd1 _08945_/B sky130_fd_sc_hd__xnor2_1
XFILLER_142_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08874_ _08874_/A _08874_/B _08873_/C _08873_/D vssd1 vssd1 vccd1 vccd1 _08874_/X
+ sky130_fd_sc_hd__or4bb_2
XFILLER_97_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_566 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09426_ _10254_/A _10932_/B vssd1 vssd1 vccd1 vccd1 _17038_/B sky130_fd_sc_hd__nand2_2
XFILLER_53_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_683 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_396 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09357_ _09357_/A _09364_/A _09357_/C vssd1 vssd1 vccd1 vccd1 _09358_/B sky130_fd_sc_hd__nor3_1
XFILLER_100_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09288_ _09289_/B _09289_/A vssd1 vssd1 vccd1 vccd1 _09296_/B sky130_fd_sc_hd__nand2b_1
XFILLER_166_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_58 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_416 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11250_ _11255_/B _11250_/B vssd1 vssd1 vccd1 vccd1 _11347_/B sky130_fd_sc_hd__nand2_1
XFILLER_158_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10201_ _10202_/A _10202_/B vssd1 vssd1 vccd1 vccd1 _10469_/A sky130_fd_sc_hd__and2b_1
X_11181_ _11181_/A _11181_/B vssd1 vssd1 vccd1 vccd1 _11182_/C sky130_fd_sc_hd__xnor2_1
XFILLER_106_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10132_ _10132_/A _10132_/B vssd1 vssd1 vccd1 vccd1 _10134_/B sky130_fd_sc_hd__xnor2_1
XFILLER_121_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10063_ _10321_/A _10446_/B _09945_/A _09943_/Y vssd1 vssd1 vccd1 vccd1 _10064_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_14940_ _17607_/Q _17477_/D _17476_/D _17608_/Q vssd1 vssd1 vccd1 vccd1 _14940_/X
+ sky130_fd_sc_hd__or4bb_1
XFILLER_76_934 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14871_ _14872_/A _14933_/B vssd1 vssd1 vccd1 vccd1 _14871_/Y sky130_fd_sc_hd__nor2_1
XFILLER_48_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16610_ _16697_/A _16610_/B vssd1 vssd1 vccd1 vccd1 _16612_/B sky130_fd_sc_hd__or2_1
XFILLER_63_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13822_ _13823_/A _13823_/B vssd1 vssd1 vccd1 vccd1 _13930_/B sky130_fd_sc_hd__and2b_1
XFILLER_35_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17590_ fanout940/X _17590_/D vssd1 vssd1 vccd1 vccd1 _17590_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16541_ _16541_/A _16541_/B vssd1 vssd1 vccd1 vccd1 _16542_/B sky130_fd_sc_hd__nor2_1
X_13753_ _13754_/B _13754_/A vssd1 vssd1 vccd1 vccd1 _13861_/B sky130_fd_sc_hd__nand2b_1
XFILLER_16_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10965_ _10965_/A _10965_/B vssd1 vssd1 vccd1 vccd1 _10966_/B sky130_fd_sc_hd__nor2_1
XFILLER_62_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_94 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12704_ _12020_/Y _12022_/Y _12053_/Y _12055_/Y _14948_/A _16011_/B vssd1 vssd1 vccd1
+ vccd1 _12704_/X sky130_fd_sc_hd__mux4_1
X_16472_ _16563_/B _16564_/A vssd1 vssd1 vccd1 vccd1 _16472_/X sky130_fd_sc_hd__or2_1
X_13684_ _13587_/B _13589_/B _13587_/A vssd1 vssd1 vccd1 vccd1 _13686_/B sky130_fd_sc_hd__o21ba_1
X_10896_ _11082_/A _11082_/B vssd1 vssd1 vccd1 vccd1 _11088_/A sky130_fd_sc_hd__or2_1
XFILLER_31_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12635_ _12478_/A _12478_/B _12477_/A vssd1 vssd1 vccd1 vccd1 _12673_/A sky130_fd_sc_hd__a21oi_1
X_15423_ _15424_/A _15424_/B vssd1 vssd1 vccd1 vccd1 _15505_/A sky130_fd_sc_hd__nor2_1
XFILLER_157_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_424 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15354_ _15355_/A _15355_/B vssd1 vssd1 vccd1 vccd1 _15356_/A sky130_fd_sc_hd__nand2_1
XFILLER_141_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12566_ _12566_/A _12566_/B vssd1 vssd1 vccd1 vccd1 _12568_/A sky130_fd_sc_hd__nor2_1
XFILLER_156_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11517_ _11629_/B _15175_/B vssd1 vssd1 vccd1 vccd1 _11595_/A sky130_fd_sc_hd__nand2_1
X_14305_ _14306_/A _14306_/B vssd1 vssd1 vccd1 vccd1 _14378_/A sky130_fd_sc_hd__nand2b_1
XFILLER_8_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15285_ _15285_/A _15285_/B vssd1 vssd1 vccd1 vccd1 _15287_/B sky130_fd_sc_hd__xnor2_1
X_12497_ _12498_/A _12498_/B _12498_/C vssd1 vssd1 vccd1 vccd1 _12499_/A sky130_fd_sc_hd__a21oi_1
XFILLER_7_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14236_ _14315_/A _14236_/B vssd1 vssd1 vccd1 vccd1 _14236_/X sky130_fd_sc_hd__and2_1
X_17024_ _17024_/A _17024_/B vssd1 vssd1 vccd1 vccd1 _17024_/X sky130_fd_sc_hd__xor2_1
XFILLER_116_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11448_ _11448_/A _11448_/B vssd1 vssd1 vccd1 vccd1 _11449_/C sky130_fd_sc_hd__and2_1
XFILLER_172_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14167_ _14167_/A _14318_/B _14366_/B _14301_/C vssd1 vssd1 vccd1 vccd1 _14245_/A
+ sky130_fd_sc_hd__and4_1
X_11379_ _11553_/A _11563_/D _11561_/D _11427_/A vssd1 vssd1 vccd1 vccd1 _11380_/C
+ sky130_fd_sc_hd__a22oi_1
XFILLER_125_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13118_ _13118_/A _13118_/B vssd1 vssd1 vccd1 vccd1 _13120_/B sky130_fd_sc_hd__nand2_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14098_ _14098_/A _14098_/B vssd1 vssd1 vccd1 vccd1 _14101_/B sky130_fd_sc_hd__nand2_1
XFILLER_113_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_508 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13049_ _13049_/A _13049_/B _13049_/C vssd1 vssd1 vccd1 vccd1 _13061_/B sky130_fd_sc_hd__nand3_1
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_720 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16808_ _16809_/A _16809_/C _15724_/X _16938_/A vssd1 vssd1 vccd1 vccd1 _16808_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_66_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16739_ _16917_/A _16791_/B _16725_/X _16738_/X vssd1 vssd1 vccd1 vccd1 _16739_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_35_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_396 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09211_ _09211_/A _09211_/B _09373_/A vssd1 vssd1 vccd1 vccd1 _09212_/B sky130_fd_sc_hd__nor3_1
XFILLER_14_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09142_ _17419_/A _17417_/A _12127_/C _12127_/D vssd1 vssd1 vccd1 vccd1 _09231_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_148_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09073_ _08985_/A _08985_/B _08985_/C vssd1 vssd1 vccd1 vccd1 _09074_/B sky130_fd_sc_hd__o21ai_1
XFILLER_30_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09975_ _09865_/A _09864_/C _09864_/B vssd1 vssd1 vccd1 vccd1 _09975_/X sky130_fd_sc_hd__a21o_1
XFILLER_103_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08926_ _08917_/X _09053_/A _09012_/A _08910_/Y vssd1 vssd1 vccd1 vccd1 _09012_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_130_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08857_ _17383_/A _11900_/D _09321_/D _17385_/A vssd1 vssd1 vccd1 vccd1 _08859_/A
+ sky130_fd_sc_hd__a22oi_1
XTAP_3605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08788_ _17393_/A _09042_/B _08779_/A _08777_/B vssd1 vssd1 vccd1 vccd1 _08796_/A
+ sky130_fd_sc_hd__a31o_1
XTAP_2915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10750_ _10750_/A _10750_/B _10750_/C vssd1 vssd1 vccd1 vccd1 _10760_/B sky130_fd_sc_hd__nand3_1
XFILLER_13_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1047 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09409_ _09410_/A _09408_/Y _10366_/A _09409_/D vssd1 vssd1 vccd1 vccd1 _09548_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_40_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10681_ _10681_/A _10681_/B vssd1 vssd1 vccd1 vccd1 _10690_/B sky130_fd_sc_hd__xnor2_1
XFILLER_71_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12420_ _12421_/A _12421_/B _12421_/C vssd1 vssd1 vccd1 vccd1 _12588_/A sky130_fd_sc_hd__a21o_1
XFILLER_138_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12351_ _12351_/A _12351_/B _12350_/X vssd1 vssd1 vccd1 vccd1 _12353_/A sky130_fd_sc_hd__or3b_1
XFILLER_126_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11302_ _11302_/A _11302_/B vssd1 vssd1 vccd1 vccd1 _16295_/A sky130_fd_sc_hd__xor2_1
XFILLER_126_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15070_ _14888_/C _14876_/D _14877_/Y _15069_/X vssd1 vssd1 vccd1 vccd1 _15071_/B
+ sky130_fd_sc_hd__o22a_1
X_12282_ _12283_/A _12283_/B vssd1 vssd1 vccd1 vccd1 _12284_/A sky130_fd_sc_hd__and2_1
XFILLER_142_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14021_ _14021_/A _14021_/B vssd1 vssd1 vccd1 vccd1 _14022_/B sky130_fd_sc_hd__or2_1
XFILLER_107_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11233_ _11155_/A _11154_/C _11154_/A vssd1 vssd1 vccd1 vccd1 _11234_/B sky130_fd_sc_hd__o21a_1
XFILLER_134_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11164_ _11164_/A _11164_/B vssd1 vssd1 vccd1 vccd1 _11165_/C sky130_fd_sc_hd__nor2_1
XFILLER_136_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10115_ _10694_/A _10241_/B _14788_/B _10359_/B vssd1 vssd1 vccd1 vccd1 _10116_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_121_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11095_ _11095_/A _11095_/B _11240_/C _11095_/D vssd1 vssd1 vccd1 vccd1 _11098_/A
+ sky130_fd_sc_hd__and4_1
X_15972_ _15972_/A _15972_/B vssd1 vssd1 vccd1 vccd1 _15973_/B sky130_fd_sc_hd__and2_1
XFILLER_1_996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14923_ _15131_/A _14922_/X _15805_/A vssd1 vssd1 vccd1 vccd1 _14923_/Y sky130_fd_sc_hd__a21oi_1
X_10046_ _10046_/A _10046_/B vssd1 vssd1 vccd1 vccd1 _10162_/C sky130_fd_sc_hd__xnor2_1
XFILLER_48_455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14854_ _15709_/A _15709_/B vssd1 vssd1 vccd1 vccd1 _15811_/B sky130_fd_sc_hd__and2_1
XFILLER_90_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13805_ _13805_/A _13805_/B vssd1 vssd1 vccd1 vccd1 _13806_/B sky130_fd_sc_hd__nor2_1
X_17573_ fanout951/X _17573_/D vssd1 vssd1 vccd1 vccd1 _17573_/Q sky130_fd_sc_hd__dfxtp_1
X_11997_ _11998_/A _11998_/B _12197_/B _11998_/D vssd1 vssd1 vccd1 vccd1 _11997_/Y
+ sky130_fd_sc_hd__nor4_1
X_14785_ _15472_/A _15541_/A vssd1 vssd1 vccd1 vccd1 _14785_/X sky130_fd_sc_hd__or2_1
XFILLER_16_341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16524_ _16524_/A _16524_/B vssd1 vssd1 vccd1 vccd1 _16525_/B sky130_fd_sc_hd__and2_1
XFILLER_72_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10948_ _10927_/X _11059_/A _10946_/X _10947_/Y vssd1 vssd1 vccd1 vccd1 _10951_/A
+ sky130_fd_sc_hd__a211o_1
X_13736_ _13736_/A _13849_/A vssd1 vssd1 vccd1 vccd1 _13739_/A sky130_fd_sc_hd__nor2_1
XFILLER_17_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_834 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_396 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16455_ _16455_/A _16455_/B vssd1 vssd1 vccd1 vccd1 _16457_/B sky130_fd_sc_hd__xnor2_1
X_10879_ _10879_/A _10879_/B vssd1 vssd1 vccd1 vccd1 _11114_/B sky130_fd_sc_hd__xnor2_1
X_13667_ _13668_/A _13668_/B vssd1 vssd1 vccd1 vccd1 _13778_/B sky130_fd_sc_hd__nor2_1
XFILLER_32_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_889 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15406_ _15406_/A _15406_/B vssd1 vssd1 vccd1 vccd1 _15408_/C sky130_fd_sc_hd__xor2_1
X_12618_ _12770_/A _12770_/B _12770_/D _12618_/D vssd1 vssd1 vccd1 vccd1 _12619_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_31_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13598_ _13598_/A _13598_/B vssd1 vssd1 vccd1 vccd1 _13600_/B sky130_fd_sc_hd__or2_1
X_16386_ _16911_/A _16386_/B vssd1 vssd1 vccd1 vccd1 _16386_/Y sky130_fd_sc_hd__nand2_1
XFILLER_157_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12549_ _13831_/S _12547_/X _12548_/Y vssd1 vssd1 vccd1 vccd1 _12549_/X sky130_fd_sc_hd__a21o_1
X_15337_ _15337_/A _15337_/B vssd1 vssd1 vccd1 vccd1 _15346_/A sky130_fd_sc_hd__xnor2_1
XFILLER_157_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_1 _17479_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15268_ _15337_/A _15268_/B vssd1 vssd1 vccd1 vccd1 _15281_/A sky130_fd_sc_hd__nand2_1
XFILLER_144_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17007_ _17007_/A _17007_/B vssd1 vssd1 vccd1 vccd1 _17037_/B sky130_fd_sc_hd__xnor2_1
XFILLER_6_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14219_ _14297_/A _14219_/B vssd1 vssd1 vccd1 vccd1 _14221_/C sky130_fd_sc_hd__and2_1
XFILLER_160_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15199_ _14887_/B _15198_/X _14924_/A vssd1 vssd1 vccd1 vccd1 _15199_/Y sky130_fd_sc_hd__a21boi_4
XFILLER_153_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout508 _17518_/Q vssd1 vssd1 vccd1 vccd1 _12592_/A sky130_fd_sc_hd__buf_2
XFILLER_141_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout519 _10638_/B vssd1 vssd1 vccd1 vccd1 _14787_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_141_975 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09760_ _09762_/B _09891_/A _09762_/A vssd1 vssd1 vccd1 vccd1 _09761_/A sky130_fd_sc_hd__a21oi_2
XFILLER_98_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_411 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09691_ _09696_/A _09696_/B vssd1 vssd1 vccd1 vccd1 _09703_/A sky130_fd_sc_hd__nor2_1
XFILLER_67_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09125_ _17417_/A _17306_/A1 _11920_/D _17419_/A vssd1 vssd1 vccd1 vccd1 _09128_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_157_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09056_ _17381_/A _12088_/D _08916_/A _08914_/Y vssd1 vssd1 vccd1 vccd1 _09057_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_108_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_972 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09958_ _09770_/Y _09830_/X _09915_/A _10059_/A vssd1 vssd1 vccd1 vccd1 _09960_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_104_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08909_ _08910_/A _08910_/B _08910_/C vssd1 vssd1 vccd1 vccd1 _09012_/A sky130_fd_sc_hd__a21o_1
XFILLER_58_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09889_ _09765_/X _09887_/Y _09885_/A _09869_/X vssd1 vssd1 vccd1 vccd1 _09912_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_85_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11920_ _17425_/A _17423_/A _12127_/D _11920_/D vssd1 vssd1 vccd1 vccd1 _12179_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_46_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_959 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11851_ _12046_/A _11851_/B vssd1 vssd1 vccd1 vccd1 _11852_/B sky130_fd_sc_hd__nand2_1
XTAP_3479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10802_ _10802_/A _10802_/B vssd1 vssd1 vccd1 vccd1 _10803_/B sky130_fd_sc_hd__nor2_1
XTAP_2767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14570_ _14570_/A _14621_/A _14570_/C vssd1 vssd1 vccd1 vccd1 _14621_/B sky130_fd_sc_hd__nand3_1
XFILLER_13_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11782_ _17476_/D _17477_/D vssd1 vssd1 vccd1 vccd1 _14924_/C sky130_fd_sc_hd__nand2b_2
XTAP_2789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10733_ _10714_/X _10728_/B _10732_/Y _10662_/X vssd1 vssd1 vccd1 vccd1 _10771_/A
+ sky130_fd_sc_hd__a211oi_2
XFILLER_15_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13521_ _13735_/B _13735_/D _13522_/D _13632_/A vssd1 vssd1 vccd1 vccd1 _13524_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_158_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_355 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16240_ _16241_/A _16241_/B _16239_/Y vssd1 vssd1 vccd1 vccd1 _16347_/A sky130_fd_sc_hd__o21ba_1
X_13452_ _13897_/A _13564_/C _13453_/C vssd1 vssd1 vccd1 vccd1 _13454_/A sky130_fd_sc_hd__a21oi_1
X_10664_ _10670_/A _10636_/Y _10651_/Y _10662_/X vssd1 vssd1 vccd1 vccd1 _10665_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_9_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12403_ _12403_/A _12403_/B vssd1 vssd1 vccd1 vccd1 _17579_/D sky130_fd_sc_hd__nand2_1
XFILLER_12_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16171_ _16355_/A _16259_/B vssd1 vssd1 vccd1 vccd1 _16172_/B sky130_fd_sc_hd__nand2_1
XFILLER_127_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13383_ _13504_/B _13382_/X _13261_/A _13263_/A vssd1 vssd1 vccd1 vccd1 _13509_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_139_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10595_ _10595_/A _10595_/B vssd1 vssd1 vccd1 vccd1 _10709_/B sky130_fd_sc_hd__xnor2_1
XFILLER_154_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12334_ _17405_/A _12334_/B _12334_/C vssd1 vssd1 vccd1 vccd1 _12336_/A sky130_fd_sc_hd__and3_1
X_15122_ _15056_/A _10543_/C _11841_/X _15102_/A _15121_/X vssd1 vssd1 vccd1 vccd1
+ _15126_/B sky130_fd_sc_hd__o311a_1
XFILLER_127_758 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_555 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15053_ _11650_/X _11675_/C _11655_/A _15052_/Y vssd1 vssd1 vccd1 vccd1 _15053_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_147_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12265_ _12437_/A _12265_/B _12265_/C vssd1 vssd1 vccd1 vccd1 _12437_/B sky130_fd_sc_hd__nand3_1
X_14004_ _14092_/B _14004_/B vssd1 vssd1 vccd1 vccd1 _14007_/A sky130_fd_sc_hd__nand2_1
XFILLER_107_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11216_ _11216_/A _11216_/B vssd1 vssd1 vccd1 vccd1 _11217_/B sky130_fd_sc_hd__xor2_1
XFILLER_123_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12196_ _12360_/B _12194_/X _11998_/A _11997_/Y vssd1 vssd1 vccd1 vccd1 _12198_/B
+ sky130_fd_sc_hd__a211oi_1
Xoutput71 _17466_/Q vssd1 vssd1 vccd1 vccd1 leds[0] sky130_fd_sc_hd__clkbuf_1
Xoutput82 _17475_/Q vssd1 vssd1 vccd1 vccd1 leds[9] sky130_fd_sc_hd__clkbuf_1
X_11147_ _11148_/A _11148_/B vssd1 vssd1 vccd1 vccd1 _11154_/A sky130_fd_sc_hd__or2_1
XFILLER_123_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput93 _17452_/Q vssd1 vssd1 vccd1 vccd1 o_wb_data[18] sky130_fd_sc_hd__clkbuf_1
XFILLER_95_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11078_ _10895_/A _10864_/Y _10881_/Y _11112_/A vssd1 vssd1 vccd1 vccd1 _11080_/C
+ sky130_fd_sc_hd__a211o_1
X_15955_ _16168_/A _16814_/A vssd1 vssd1 vccd1 vccd1 _15955_/Y sky130_fd_sc_hd__nor2_1
XFILLER_76_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14906_ _15314_/A _14906_/B _15151_/B vssd1 vssd1 vccd1 vccd1 _14906_/X sky130_fd_sc_hd__or3_1
X_10029_ _10029_/A _10029_/B _10029_/C vssd1 vssd1 vccd1 vccd1 _10057_/A sky130_fd_sc_hd__or3_1
XFILLER_37_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15886_ _15884_/Y _15885_/Y _15523_/A vssd1 vssd1 vccd1 vccd1 _15886_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_36_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14837_ _14837_/A _17070_/B vssd1 vssd1 vccd1 vccd1 _14837_/Y sky130_fd_sc_hd__nor2_1
XFILLER_63_255 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17556_ fanout935/X _17556_/D vssd1 vssd1 vccd1 vccd1 _17556_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14768_ _16965_/C _16974_/A vssd1 vssd1 vccd1 vccd1 _16970_/B sky130_fd_sc_hd__or2_1
X_16507_ _16507_/A _16507_/B vssd1 vssd1 vccd1 vccd1 _16509_/C sky130_fd_sc_hd__xnor2_1
X_13719_ _13720_/A _13720_/B vssd1 vssd1 vccd1 vccd1 _13824_/A sky130_fd_sc_hd__nand2_1
X_17487_ fanout942/X _17487_/D vssd1 vssd1 vccd1 vccd1 _17487_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14699_ _14699_/A _14699_/B vssd1 vssd1 vccd1 vccd1 _14701_/B sky130_fd_sc_hd__xor2_1
XFILLER_108_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16438_ _16439_/A _16439_/B vssd1 vssd1 vccd1 vccd1 _16527_/B sky130_fd_sc_hd__nor2_1
XFILLER_31_174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16369_ _16369_/A _16369_/B vssd1 vssd1 vccd1 vccd1 _16372_/A sky130_fd_sc_hd__xor2_2
XFILLER_157_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout305 _14733_/S vssd1 vssd1 vccd1 vccd1 _14757_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_141_761 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout316 _17610_/Q vssd1 vssd1 vccd1 vccd1 _17477_/D sky130_fd_sc_hd__clkbuf_8
XFILLER_98_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout327 _14050_/B vssd1 vssd1 vccd1 vccd1 _14213_/B sky130_fd_sc_hd__clkbuf_4
X_09812_ _09812_/A _09812_/B _09812_/C vssd1 vssd1 vccd1 vccd1 _09813_/C sky130_fd_sc_hd__or3_1
Xfanout338 _13069_/A vssd1 vssd1 vccd1 vccd1 _17100_/C sky130_fd_sc_hd__clkbuf_4
Xfanout349 _17538_/Q vssd1 vssd1 vccd1 vccd1 _09360_/A sky130_fd_sc_hd__buf_2
XFILLER_87_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09743_ _09621_/A _09621_/B _09621_/C vssd1 vssd1 vccd1 vccd1 _09743_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_67_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09674_ _09674_/A _09674_/B _09819_/A vssd1 vssd1 vccd1 vccd1 _09675_/C sky130_fd_sc_hd__nor3_1
XFILLER_82_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09108_ _09108_/A _09108_/B vssd1 vssd1 vccd1 vccd1 _09110_/B sky130_fd_sc_hd__xnor2_1
XFILLER_109_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10380_ _10487_/A _10379_/B _10379_/A vssd1 vssd1 vccd1 vccd1 _10382_/B sky130_fd_sc_hd__o21ba_1
XFILLER_108_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09039_ _09039_/A _09039_/B vssd1 vssd1 vccd1 vccd1 _09047_/A sky130_fd_sc_hd__xnor2_1
XFILLER_105_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12050_ _10016_/D _15898_/A _12050_/S vssd1 vssd1 vccd1 vccd1 _12051_/B sky130_fd_sc_hd__mux2_1
XFILLER_105_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11001_ _10977_/X _11051_/A _10999_/X _11000_/Y vssd1 vssd1 vccd1 vccd1 _11157_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_120_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout850 _14788_/B vssd1 vssd1 vccd1 vccd1 _10963_/C sky130_fd_sc_hd__clkbuf_4
Xfanout861 _10359_/B vssd1 vssd1 vccd1 vccd1 _10703_/B sky130_fd_sc_hd__clkbuf_2
Xfanout872 _10479_/B vssd1 vssd1 vccd1 vccd1 _11005_/B sky130_fd_sc_hd__clkbuf_2
Xfanout883 _11427_/C vssd1 vssd1 vccd1 vccd1 _10805_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_46_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout894 _17480_/Q vssd1 vssd1 vccd1 vccd1 _11006_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_19_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15740_ _15740_/A _15740_/B vssd1 vssd1 vccd1 vccd1 _15741_/B sky130_fd_sc_hd__xor2_2
XFILLER_93_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12952_ _13092_/B _12952_/B vssd1 vssd1 vccd1 vccd1 _12955_/B sky130_fd_sc_hd__nand2_1
XFILLER_45_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11903_ _11903_/A _11903_/B vssd1 vssd1 vccd1 vccd1 _11906_/A sky130_fd_sc_hd__xnor2_1
XTAP_3265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15671_ _15671_/A _15671_/B vssd1 vssd1 vccd1 vccd1 _15673_/B sky130_fd_sc_hd__xor2_1
XFILLER_93_66 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12883_ _12884_/A _12884_/B vssd1 vssd1 vccd1 vccd1 _13033_/B sky130_fd_sc_hd__nand2b_1
XTAP_2531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17410_ input51/X _17422_/A2 _17409_/X _17422_/C1 vssd1 vssd1 vccd1 vccd1 _17533_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_33_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14622_ _14661_/A _14622_/B vssd1 vssd1 vccd1 vccd1 _14624_/B sky130_fd_sc_hd__or2_1
XTAP_2553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11834_ _12320_/D _13067_/D _12050_/S vssd1 vssd1 vccd1 vccd1 _11835_/B sky130_fd_sc_hd__mux2_1
XTAP_2564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_748 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17341_ input50/X _17353_/B _17353_/C vssd1 vssd1 vccd1 vccd1 _17341_/X sky130_fd_sc_hd__or3_1
XTAP_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14553_ _14553_/A _14553_/B vssd1 vssd1 vccd1 vccd1 _14555_/A sky130_fd_sc_hd__nor2_1
X_11765_ _16568_/A _11760_/X _11764_/X vssd1 vssd1 vccd1 vccd1 _16866_/B sky130_fd_sc_hd__a21oi_2
XFILLER_159_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10716_ _10716_/A _10716_/B vssd1 vssd1 vccd1 vccd1 _10722_/A sky130_fd_sc_hd__xnor2_1
X_13504_ _13504_/A _13504_/B vssd1 vssd1 vccd1 vccd1 _13506_/B sky130_fd_sc_hd__or2_1
X_17272_ _17458_/Q _17290_/A2 _17270_/X _17271_/X _17293_/C1 vssd1 vssd1 vccd1 vccd1
+ _17458_/D sky130_fd_sc_hd__o221a_1
X_11696_ _15525_/A _15447_/A _11672_/Y _11624_/Y vssd1 vssd1 vccd1 vccd1 _15614_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_14484_ _14641_/B _14301_/C _14485_/D _14641_/A vssd1 vssd1 vccd1 vccd1 _14486_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_174_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16223_ _16205_/X _16207_/X _16222_/Y _16494_/B1 _14778_/B vssd1 vssd1 vccd1 vccd1
+ _16224_/A sky130_fd_sc_hd__a32o_1
XFILLER_173_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10647_ _10648_/A _10646_/Y _10745_/C _10647_/D vssd1 vssd1 vccd1 vccd1 _10742_/A
+ sky130_fd_sc_hd__and4bb_1
X_13435_ _13435_/A _13586_/A vssd1 vssd1 vccd1 vccd1 _13438_/A sky130_fd_sc_hd__or2_1
XFILLER_127_511 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16154_ _16155_/A _16155_/B vssd1 vssd1 vccd1 vccd1 _16270_/A sky130_fd_sc_hd__nor2_1
XFILLER_127_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13366_ _13366_/A _13366_/B vssd1 vssd1 vccd1 vccd1 _13368_/B sky130_fd_sc_hd__xnor2_1
X_10578_ _10325_/A _10329_/B _10579_/A _10577_/X vssd1 vssd1 vccd1 vccd1 _10579_/B
+ sky130_fd_sc_hd__a211oi_1
X_15105_ _11679_/A _11679_/B _16389_/A vssd1 vssd1 vccd1 vccd1 _15106_/B sky130_fd_sc_hd__o21a_1
XFILLER_155_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_588 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12317_ _12186_/A _12186_/B _12189_/A vssd1 vssd1 vccd1 vccd1 _12357_/A sky130_fd_sc_hd__o21ai_1
X_16085_ _16197_/A _16085_/B vssd1 vssd1 vccd1 vccd1 _16086_/C sky130_fd_sc_hd__and2b_1
X_13297_ _13643_/A _13735_/D _13159_/A _13157_/B vssd1 vssd1 vccd1 vccd1 _13304_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_5_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_227 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12248_ _12429_/B _12248_/B vssd1 vssd1 vccd1 vccd1 _12250_/B sky130_fd_sc_hd__and2b_1
X_15036_ _14949_/Y _14952_/Y _15036_/S vssd1 vssd1 vccd1 vccd1 _15037_/B sky130_fd_sc_hd__mux2_1
XFILLER_142_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12179_ _12179_/A _12179_/B _12179_/C vssd1 vssd1 vccd1 vccd1 _12180_/B sky130_fd_sc_hd__nor3_1
XFILLER_68_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16987_ _17119_/A _16987_/B vssd1 vssd1 vccd1 vccd1 _16989_/B sky130_fd_sc_hd__nand2_1
XFILLER_96_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15938_ _15939_/A _15939_/B vssd1 vssd1 vccd1 vccd1 _16072_/B sky130_fd_sc_hd__and2_1
XFILLER_64_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_840 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15869_ _15414_/B _15746_/X _15750_/X vssd1 vssd1 vccd1 vccd1 _15871_/B sky130_fd_sc_hd__o21ba_1
XFILLER_37_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17608_ fanout949/X _17608_/D vssd1 vssd1 vccd1 vccd1 _17608_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_36_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09390_ _09343_/X _09344_/Y _09387_/A _09388_/Y vssd1 vssd1 vccd1 vccd1 _09393_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_145_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17539_ fanout947/X _17539_/D vssd1 vssd1 vccd1 vccd1 _17539_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_639 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_875 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_823 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout124 _17244_/B vssd1 vssd1 vccd1 vccd1 _17292_/B sky130_fd_sc_hd__buf_2
XFILLER_160_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout135 _15339_/Y vssd1 vssd1 vccd1 vccd1 _15755_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_101_411 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout146 _14973_/Y vssd1 vssd1 vccd1 vccd1 _16165_/A sky130_fd_sc_hd__clkbuf_4
Xfanout157 _17424_/A2 vssd1 vssd1 vccd1 vccd1 _17426_/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_113_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout168 _16497_/D vssd1 vssd1 vccd1 vccd1 _16662_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_101_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout179 _15551_/Y vssd1 vssd1 vccd1 vccd1 _16758_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_41_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09726_ _09730_/C _10421_/D _09587_/A _09585_/Y vssd1 vssd1 vccd1 vccd1 _09727_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_28_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09657_ _09786_/A _09657_/B vssd1 vssd1 vccd1 vccd1 _09658_/B sky130_fd_sc_hd__nor2_1
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09588_ _09589_/B _09589_/A vssd1 vssd1 vccd1 vccd1 _09588_/X sky130_fd_sc_hd__and2b_1
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11550_ _11542_/A _11541_/C _11541_/A vssd1 vssd1 vccd1 vccd1 _11584_/B sky130_fd_sc_hd__o21a_1
XFILLER_51_792 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_280 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10501_ _10501_/A _10501_/B vssd1 vssd1 vccd1 vccd1 _10503_/C sky130_fd_sc_hd__xnor2_1
XFILLER_10_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11481_ _11518_/B _14850_/A _11561_/C _11518_/A vssd1 vssd1 vccd1 vccd1 _11481_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_7_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13220_ _13220_/A _13220_/B _13220_/C vssd1 vssd1 vccd1 vccd1 _13221_/B sky130_fd_sc_hd__nand3_1
X_10432_ _10753_/A _10545_/D _10180_/C vssd1 vssd1 vccd1 vccd1 _10432_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_136_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13151_ _13151_/A _13151_/B vssd1 vssd1 vccd1 vccd1 _13154_/A sky130_fd_sc_hd__xnor2_1
XFILLER_88_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10363_ _10364_/A _10364_/B vssd1 vssd1 vccd1 vccd1 _10374_/B sky130_fd_sc_hd__nor2_1
XFILLER_164_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12102_ _17379_/A _12592_/B _12447_/B _12445_/C vssd1 vssd1 vccd1 vccd1 _12103_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_124_558 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13082_ _13083_/A _13213_/A _13083_/C vssd1 vssd1 vccd1 vccd1 _13084_/A sky130_fd_sc_hd__o21a_1
XFILLER_112_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10294_ _10045_/C _10545_/D _10288_/A _10172_/Y vssd1 vssd1 vccd1 vccd1 _10296_/C
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_105_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16910_ _16910_/A _16910_/B vssd1 vssd1 vccd1 vccd1 _16911_/B sky130_fd_sc_hd__xor2_1
XFILLER_2_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12033_ _08969_/C _12032_/Y _14911_/B vssd1 vssd1 vccd1 vccd1 _12033_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_78_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16841_ _16841_/A _16841_/B vssd1 vssd1 vccd1 vccd1 _16843_/B sky130_fd_sc_hd__xnor2_1
Xfanout680 _08860_/B vssd1 vssd1 vccd1 vccd1 _09926_/B sky130_fd_sc_hd__buf_2
XFILLER_77_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout691 fanout699/X vssd1 vssd1 vccd1 vccd1 _14213_/C sky130_fd_sc_hd__clkbuf_4
X_16772_ _16688_/A _16687_/B _16685_/X vssd1 vssd1 vccd1 vccd1 _16774_/B sky130_fd_sc_hd__a21o_1
X_13984_ _13985_/B _13985_/A vssd1 vssd1 vccd1 vccd1 _14072_/B sky130_fd_sc_hd__and2b_1
XFILLER_46_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15723_ _16315_/B _16747_/A vssd1 vssd1 vccd1 vccd1 _15730_/A sky130_fd_sc_hd__nor2_1
XTAP_3051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12935_ _12935_/A _12935_/B vssd1 vssd1 vccd1 vccd1 _12938_/C sky130_fd_sc_hd__or2_1
XFILLER_18_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15654_ _15743_/A _15654_/B vssd1 vssd1 vccd1 vccd1 _15656_/B sky130_fd_sc_hd__nor2_1
XTAP_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12866_ _14925_/A _12866_/B vssd1 vssd1 vccd1 vccd1 _12866_/Y sky130_fd_sc_hd__nor2_1
XTAP_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14605_ _14606_/B _14606_/A vssd1 vssd1 vccd1 vccd1 _14646_/B sky130_fd_sc_hd__nand2b_1
XTAP_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11817_ _11814_/Y _11816_/Y _12212_/S vssd1 vssd1 vccd1 vccd1 _11818_/B sky130_fd_sc_hd__mux2_1
XTAP_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15585_ _15499_/A _15499_/B _15488_/Y vssd1 vssd1 vccd1 vccd1 _15587_/B sky130_fd_sc_hd__o21ai_1
X_12797_ _12798_/A _12798_/B _12798_/C vssd1 vssd1 vccd1 vccd1 _12799_/A sky130_fd_sc_hd__a21oi_1
XTAP_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17324_ _09030_/C _17360_/A2 _17323_/X _17426_/C1 vssd1 vssd1 vccd1 vccd1 _17491_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_14_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14536_ _14415_/X _14534_/B _14534_/Y _14280_/X vssd1 vssd1 vccd1 vccd1 _14536_/X
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11748_ _16794_/A _11748_/B vssd1 vssd1 vccd1 vccd1 _16727_/B sky130_fd_sc_hd__and2_1
XFILLER_147_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17255_ _17594_/Q _17291_/A2 _17291_/B1 vssd1 vssd1 vccd1 vccd1 _17255_/X sky130_fd_sc_hd__a21o_1
XFILLER_147_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14467_ _14524_/A _14524_/B vssd1 vssd1 vccd1 vccd1 _14469_/B sky130_fd_sc_hd__xnor2_1
X_11679_ _11679_/A _11679_/B vssd1 vssd1 vccd1 vccd1 _15106_/A sky130_fd_sc_hd__nand2_1
X_16206_ _16206_/A _16206_/B vssd1 vssd1 vccd1 vccd1 _16207_/C sky130_fd_sc_hd__nor2_1
X_13418_ _13418_/A _13418_/B vssd1 vssd1 vccd1 vccd1 _13420_/B sky130_fd_sc_hd__and2_1
XFILLER_127_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17186_ input29/X wire215/X vssd1 vssd1 vccd1 vccd1 _17429_/B sky130_fd_sc_hd__nand2_1
X_14398_ _14395_/Y _14396_/X _14316_/A _14332_/X vssd1 vssd1 vccd1 vccd1 _14400_/C
+ sky130_fd_sc_hd__o211ai_1
XFILLER_115_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16137_ _16137_/A _16250_/A vssd1 vssd1 vccd1 vccd1 _16140_/A sky130_fd_sc_hd__or2_1
XFILLER_143_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13349_ _13349_/A _13349_/B vssd1 vssd1 vccd1 vccd1 _13368_/A sky130_fd_sc_hd__xnor2_1
XFILLER_52_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16068_ _16068_/A _16068_/B vssd1 vssd1 vccd1 vccd1 _16070_/B sky130_fd_sc_hd__xor2_1
XFILLER_143_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15019_ _15314_/A _14899_/C _15018_/X _15147_/D vssd1 vssd1 vccd1 vccd1 _15402_/B
+ sky130_fd_sc_hd__o22ai_4
X_08890_ _09020_/A _09020_/B vssd1 vssd1 vccd1 vccd1 _08904_/C sky130_fd_sc_hd__nand2_1
XFILLER_69_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09511_ _09511_/A _09511_/B vssd1 vssd1 vccd1 vccd1 _09522_/A sky130_fd_sc_hd__nor2_1
XFILLER_37_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09442_ _09730_/C _09058_/C _09302_/A _09300_/Y vssd1 vssd1 vccd1 vccd1 _09443_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_80_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_832 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_556 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09373_ _09373_/A _09373_/B vssd1 vssd1 vccd1 vccd1 _09385_/A sky130_fd_sc_hd__nor2_1
XFILLER_40_718 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_497 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_834 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09709_ _09709_/A _09709_/B vssd1 vssd1 vccd1 vccd1 _09717_/A sky130_fd_sc_hd__xnor2_1
X_10981_ _10974_/A _10973_/B _10973_/A vssd1 vssd1 vccd1 vccd1 _10985_/A sky130_fd_sc_hd__o21ba_1
XFILLER_62_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xwb_buttons_leds_965 vssd1 vssd1 vccd1 vccd1 wb_buttons_leds_965/HI led_enb[7] sky130_fd_sc_hd__conb_1
XFILLER_83_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12720_ _12720_/A _12720_/B vssd1 vssd1 vccd1 vccd1 _12727_/A sky130_fd_sc_hd__xor2_1
XFILLER_83_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12651_ _12651_/A _12651_/B vssd1 vssd1 vccd1 vccd1 _12654_/A sky130_fd_sc_hd__nand2_1
XFILLER_31_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11602_ _11568_/A _11568_/C _11568_/B vssd1 vssd1 vccd1 vccd1 _11603_/C sky130_fd_sc_hd__a21oi_1
X_15370_ _11692_/B _11691_/B _11693_/Y vssd1 vssd1 vccd1 vccd1 _15370_/X sky130_fd_sc_hd__a21o_1
X_12582_ _12583_/A _12583_/B vssd1 vssd1 vccd1 vccd1 _12761_/B sky130_fd_sc_hd__and2b_1
XFILLER_12_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14321_ _14387_/A _14383_/B _14321_/C vssd1 vssd1 vccd1 vccd1 _14389_/B sky130_fd_sc_hd__and3_1
X_11533_ _11534_/A _11534_/B vssd1 vssd1 vccd1 vccd1 _11541_/A sky130_fd_sc_hd__or2_1
XFILLER_168_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17040_ _17040_/A _17040_/B vssd1 vssd1 vccd1 vccd1 _17085_/A sky130_fd_sc_hd__nor2_1
X_11464_ _11708_/A _11464_/B vssd1 vssd1 vccd1 vccd1 _11465_/B sky130_fd_sc_hd__or2_1
X_14252_ _14252_/A _14252_/B _14252_/C vssd1 vssd1 vccd1 vccd1 _14253_/B sky130_fd_sc_hd__and3_1
XFILLER_171_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10415_ _10415_/A _10513_/A vssd1 vssd1 vccd1 vccd1 _10423_/A sky130_fd_sc_hd__nor2_1
X_13203_ _13203_/A vssd1 vssd1 vccd1 vccd1 _13332_/B sky130_fd_sc_hd__inv_2
X_11395_ _11395_/A _11395_/B _11435_/A vssd1 vssd1 vccd1 vccd1 _11396_/C sky130_fd_sc_hd__nand3_1
XFILLER_137_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14183_ _14273_/B _14184_/C vssd1 vssd1 vccd1 vccd1 _14185_/B sky130_fd_sc_hd__and2_1
XFILLER_48_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13134_ _13137_/A vssd1 vssd1 vccd1 vccd1 _13134_/Y sky130_fd_sc_hd__inv_2
X_10346_ _10349_/A _10349_/B vssd1 vssd1 vccd1 vccd1 _17105_/A sky130_fd_sc_hd__nor2_1
XFILLER_98_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13065_ _13065_/A _13065_/B _13065_/C vssd1 vssd1 vccd1 vccd1 _13075_/B sky130_fd_sc_hd__nand3_1
XFILLER_151_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10277_ _14788_/A _10993_/D _10167_/A _10165_/Y vssd1 vssd1 vccd1 vccd1 _10278_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_151_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12016_ _12016_/A _12016_/B vssd1 vssd1 vccd1 vccd1 _12377_/A sky130_fd_sc_hd__nand2_1
XFILLER_78_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16824_ _16935_/A _16760_/B _16761_/A _16759_/B vssd1 vssd1 vccd1 vccd1 _16830_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_66_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16755_ _16661_/X _16665_/B _16663_/B vssd1 vssd1 vccd1 vccd1 _16762_/A sky130_fd_sc_hd__o21ai_1
X_13967_ _13967_/A _13967_/B vssd1 vssd1 vccd1 vccd1 _13969_/A sky130_fd_sc_hd__nor2_1
XFILLER_47_873 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15706_ _15705_/A _15705_/B _15705_/C vssd1 vssd1 vccd1 vccd1 _15706_/X sky130_fd_sc_hd__a21o_1
X_12918_ _13065_/A _12918_/B _12918_/C vssd1 vssd1 vccd1 vccd1 _13065_/B sky130_fd_sc_hd__nand3_1
XFILLER_34_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16686_ _16686_/A _16686_/B _16684_/Y vssd1 vssd1 vccd1 vccd1 _16687_/B sky130_fd_sc_hd__or3b_1
XFILLER_34_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13898_ _13898_/A _13898_/B vssd1 vssd1 vccd1 vccd1 _13901_/B sky130_fd_sc_hd__xnor2_1
XFILLER_55_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15637_ _16021_/A _08731_/A _15262_/A vssd1 vssd1 vccd1 vccd1 _15639_/B sky130_fd_sc_hd__a21bo_1
XTAP_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12849_ _13833_/S _12849_/B vssd1 vssd1 vccd1 vccd1 _12849_/X sky130_fd_sc_hd__or2_1
XFILLER_15_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15568_ _15568_/A _15568_/B vssd1 vssd1 vccd1 vccd1 _15570_/A sky130_fd_sc_hd__and2_1
XFILLER_21_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17307_ input63/X _17321_/B _17321_/C vssd1 vssd1 vccd1 vccd1 _17307_/X sky130_fd_sc_hd__or3_1
XFILLER_9_74 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14519_ _14519_/A _14519_/B _14519_/C vssd1 vssd1 vccd1 vccd1 _14519_/X sky130_fd_sc_hd__and3_1
X_15499_ _15499_/A _15499_/B vssd1 vssd1 vccd1 vccd1 _15501_/C sky130_fd_sc_hd__xor2_1
XFILLER_119_127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17238_ _17556_/Q _17292_/B vssd1 vssd1 vccd1 vccd1 _17238_/X sky130_fd_sc_hd__and2_1
XFILLER_174_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17169_ _16304_/A _17167_/X _17168_/Y _17166_/X vssd1 vssd1 vccd1 vccd1 _17169_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_171_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09991_ _10004_/B _10004_/C _10004_/A vssd1 vssd1 vccd1 vccd1 _09991_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_131_826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08942_ _09327_/C _11815_/B vssd1 vssd1 vccd1 vccd1 _08943_/B sky130_fd_sc_hd__nand2_1
XFILLER_9_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_902 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08873_ _08874_/A _08874_/B _08873_/C _08873_/D vssd1 vssd1 vccd1 vccd1 _08873_/X
+ sky130_fd_sc_hd__and4bb_1
XFILLER_96_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_924 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_583 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09425_ _10126_/B _10932_/B vssd1 vssd1 vccd1 vccd1 _16933_/A sky130_fd_sc_hd__nand2_2
XFILLER_25_578 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09356_ _09479_/A _09479_/B vssd1 vssd1 vccd1 vccd1 _09366_/B sky130_fd_sc_hd__nand2b_1
XFILLER_100_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09287_ _09421_/A _09285_/X _17081_/B _16990_/A vssd1 vssd1 vccd1 vccd1 _09289_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_100_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_778 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10200_ _10200_/A _10200_/B vssd1 vssd1 vccd1 vccd1 _10202_/B sky130_fd_sc_hd__nor2_1
XFILLER_107_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11180_ _11180_/A _11180_/B vssd1 vssd1 vccd1 vccd1 _11181_/B sky130_fd_sc_hd__xor2_2
XFILLER_133_130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10131_ _10132_/B _10132_/A vssd1 vssd1 vccd1 vccd1 _10138_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10062_ _10321_/A _10062_/B _10062_/C vssd1 vssd1 vccd1 vccd1 _10198_/A sky130_fd_sc_hd__and3_1
XFILLER_87_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_946 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14870_ _14831_/Y _17151_/B _16485_/A _14869_/X vssd1 vssd1 vccd1 vccd1 _17575_/D
+ sky130_fd_sc_hd__a31o_2
XFILLER_47_136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13821_ _14254_/A _13522_/D _13705_/A _13703_/A vssd1 vssd1 vccd1 vccd1 _13823_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_75_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16540_ _16627_/A vssd1 vssd1 vccd1 vccd1 _16542_/A sky130_fd_sc_hd__inv_2
X_13752_ _13642_/A _13644_/B _13642_/B vssd1 vssd1 vccd1 vccd1 _13754_/B sky130_fd_sc_hd__o21ba_1
X_10964_ _10963_/B _10963_/C _10703_/B _10963_/A vssd1 vssd1 vccd1 vccd1 _10965_/B
+ sky130_fd_sc_hd__a22oi_1
XFILLER_44_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12703_ _12701_/Y _12702_/X _13516_/S vssd1 vssd1 vccd1 vccd1 _12703_/X sky130_fd_sc_hd__mux2_1
X_16471_ _16470_/A _16470_/B _16470_/C vssd1 vssd1 vccd1 vccd1 _16564_/A sky130_fd_sc_hd__a21oi_1
X_13683_ _13683_/A _13683_/B vssd1 vssd1 vccd1 vccd1 _13686_/A sky130_fd_sc_hd__xor2_1
XFILLER_16_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10895_ _10895_/A _11080_/A vssd1 vssd1 vccd1 vccd1 _11082_/B sky130_fd_sc_hd__and2_1
XFILLER_71_695 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15422_ _15422_/A _15422_/B vssd1 vssd1 vccd1 vccd1 _15424_/B sky130_fd_sc_hd__xor2_1
X_12634_ _12518_/A _12518_/B _12516_/Y vssd1 vssd1 vccd1 vccd1 _12675_/A sky130_fd_sc_hd__a21bo_1
XFILLER_169_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15353_ _15750_/A _15397_/A _15279_/A _15276_/Y vssd1 vssd1 vccd1 vccd1 _15355_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_12_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12565_ _12722_/A _12722_/B _13348_/B _12871_/B vssd1 vssd1 vccd1 vccd1 _12566_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_141_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14304_ _14304_/A _14304_/B vssd1 vssd1 vccd1 vccd1 _14306_/B sky130_fd_sc_hd__xnor2_1
X_11516_ _11522_/A _11522_/B vssd1 vssd1 vccd1 vccd1 _11523_/A sky130_fd_sc_hd__nor2_1
XFILLER_11_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15284_ _15285_/A _15285_/B vssd1 vssd1 vccd1 vccd1 _15352_/A sky130_fd_sc_hd__or2_1
XFILLER_157_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12496_ _12496_/A _12496_/B vssd1 vssd1 vccd1 vccd1 _12498_/C sky130_fd_sc_hd__xor2_1
XFILLER_138_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17023_ _17023_/A _17023_/B vssd1 vssd1 vccd1 vccd1 _17024_/B sky130_fd_sc_hd__nand2_1
X_14235_ _14235_/A _14235_/B vssd1 vssd1 vccd1 vccd1 _14236_/B sky130_fd_sc_hd__nand2_1
X_11447_ _11447_/A _11447_/B vssd1 vssd1 vccd1 vccd1 _11448_/B sky130_fd_sc_hd__nand2_1
XFILLER_171_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_480 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11378_ _11553_/B _15238_/A vssd1 vssd1 vccd1 vccd1 _11380_/B sky130_fd_sc_hd__nand2_1
XFILLER_124_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14166_ _14318_/B _14366_/B _14301_/C _14318_/A vssd1 vssd1 vccd1 vccd1 _14170_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_113_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13117_ _13117_/A _13117_/B _13117_/C vssd1 vssd1 vccd1 vccd1 _13118_/B sky130_fd_sc_hd__nand3_1
X_10329_ _10450_/A _10329_/B _10329_/C vssd1 vssd1 vccd1 vccd1 _10451_/A sky130_fd_sc_hd__and3_1
XFILLER_140_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14097_ _14098_/A _14098_/B vssd1 vssd1 vccd1 vccd1 _14188_/B sky130_fd_sc_hd__or2_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13048_ _13049_/A _13049_/B _13049_/C vssd1 vssd1 vccd1 vccd1 _13061_/A sky130_fd_sc_hd__a21o_1
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16807_ _16807_/A _16935_/B vssd1 vssd1 vccd1 vccd1 _16811_/A sky130_fd_sc_hd__nand2_1
XFILLER_26_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14999_ _15100_/A _14999_/B vssd1 vssd1 vccd1 vccd1 _14999_/Y sky130_fd_sc_hd__nand2_1
XFILLER_35_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16738_ _16922_/A _16794_/B _16728_/Y _16737_/X vssd1 vssd1 vccd1 vccd1 _16738_/X
+ sky130_fd_sc_hd__a31o_2
X_16669_ _16667_/A _16938_/D _16670_/A _16814_/A _16813_/B vssd1 vssd1 vccd1 vccd1
+ _16671_/B sky130_fd_sc_hd__o32a_1
XFILLER_50_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09210_ _09211_/B _09373_/A _09211_/A vssd1 vssd1 vccd1 vccd1 _09212_/A sky130_fd_sc_hd__o21a_1
XFILLER_148_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09141_ _17417_/A _12127_/C _12127_/D _17419_/A vssd1 vssd1 vccd1 vccd1 _09143_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_147_200 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09072_ _09071_/A _09259_/A _08930_/X _09018_/Y vssd1 vssd1 vccd1 vccd1 _09119_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_135_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_303 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_280 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09974_ _09885_/A _09885_/B _09885_/C vssd1 vssd1 vccd1 vccd1 _10029_/B sky130_fd_sc_hd__a21oi_1
XFILLER_103_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08925_ _09012_/A _08910_/Y _08917_/X _09053_/A vssd1 vssd1 vccd1 vccd1 _08927_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_69_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08856_ _08856_/A _08856_/B vssd1 vssd1 vccd1 vccd1 _08866_/A sky130_fd_sc_hd__xnor2_1
XTAP_3606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_478 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08787_ _08798_/A _08787_/B _17522_/Q _09319_/D vssd1 vssd1 vccd1 vccd1 _08821_/A
+ sky130_fd_sc_hd__and4b_1
XFILLER_45_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_670 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_448 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09408_ _10236_/B _09843_/C _09985_/D _10236_/A vssd1 vssd1 vccd1 vccd1 _09408_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_80_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10680_ _10673_/A _10673_/B _10674_/Y vssd1 vssd1 vccd1 vccd1 _10690_/A sky130_fd_sc_hd__a21oi_1
XFILLER_41_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09339_ _09339_/A _09344_/B _09339_/C vssd1 vssd1 vccd1 vccd1 _09391_/C sky130_fd_sc_hd__or3_2
XFILLER_138_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12350_ _12517_/A _12350_/B vssd1 vssd1 vccd1 vccd1 _12350_/X sky130_fd_sc_hd__and2_1
X_11301_ _11711_/A _11711_/B vssd1 vssd1 vccd1 vccd1 _11302_/B sky130_fd_sc_hd__and2b_1
XFILLER_126_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12281_ _12281_/A _12281_/B vssd1 vssd1 vccd1 vccd1 _12283_/B sky130_fd_sc_hd__xnor2_1
XFILLER_5_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11232_ _11232_/A _11232_/B vssd1 vssd1 vccd1 vccd1 _11302_/A sky130_fd_sc_hd__xnor2_1
XFILLER_4_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14020_ _14021_/A _14021_/B vssd1 vssd1 vccd1 vccd1 _14113_/B sky130_fd_sc_hd__nand2_1
XFILLER_84_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_910 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11163_ _10545_/C _11841_/B _10756_/A _10754_/Y vssd1 vssd1 vccd1 vccd1 _11165_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_1_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10114_ _10241_/B _14788_/B _10359_/B _10694_/A vssd1 vssd1 vccd1 vccd1 _10116_/A
+ sky130_fd_sc_hd__a22oi_1
X_11094_ _11099_/A _11099_/B vssd1 vssd1 vccd1 vccd1 _11101_/A sky130_fd_sc_hd__nor2_1
X_15971_ _15972_/A _15972_/B vssd1 vssd1 vccd1 vccd1 _16080_/B sky130_fd_sc_hd__nor2_1
XFILLER_121_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14922_ _14920_/X _14921_/X _15254_/S vssd1 vssd1 vccd1 vccd1 _14922_/X sky130_fd_sc_hd__mux2_1
XFILLER_103_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10045_ _10162_/A _10044_/Y _10045_/C _10543_/B vssd1 vssd1 vccd1 vccd1 _10170_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_48_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14853_ _15624_/A _15541_/A _15541_/B vssd1 vssd1 vccd1 vccd1 _15709_/B sky130_fd_sc_hd__and3_1
XFILLER_76_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13804_ _13805_/A _13805_/B vssd1 vssd1 vccd1 vccd1 _13915_/B sky130_fd_sc_hd__and2_1
X_17572_ fanout953/X _17572_/D vssd1 vssd1 vccd1 vccd1 _17572_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14784_ _14784_/A _15624_/A vssd1 vssd1 vccd1 vccd1 _15622_/B sky130_fd_sc_hd__or2_1
X_11996_ _12197_/A _11994_/X _09248_/B _09248_/Y vssd1 vssd1 vccd1 vccd1 _11998_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_72_960 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16523_ _16524_/A _16524_/B vssd1 vssd1 vccd1 vccd1 _16616_/B sky130_fd_sc_hd__nor2_1
XFILLER_16_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13735_ _13735_/A _13735_/B _13846_/B _13735_/D vssd1 vssd1 vccd1 vccd1 _13849_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_32_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10947_ _10946_/A _10946_/B _10946_/C vssd1 vssd1 vccd1 vccd1 _10947_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_91_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_846 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16454_ _16454_/A _16454_/B vssd1 vssd1 vccd1 vccd1 _16455_/B sky130_fd_sc_hd__xor2_1
X_13666_ _14215_/A _13866_/D vssd1 vssd1 vccd1 vccd1 _13668_/B sky130_fd_sc_hd__nand2_1
X_10878_ _10878_/A _11121_/A vssd1 vssd1 vccd1 vccd1 _11114_/A sky130_fd_sc_hd__or2_1
X_15405_ _16315_/C _16262_/A vssd1 vssd1 vccd1 vccd1 _15406_/B sky130_fd_sc_hd__nor2_1
X_12617_ _12770_/B _12770_/D _12618_/D _12770_/A vssd1 vssd1 vccd1 vccd1 _12619_/A
+ sky130_fd_sc_hd__a22oi_1
X_16385_ _16385_/A _16385_/B vssd1 vssd1 vccd1 vccd1 _16386_/B sky130_fd_sc_hd__xor2_2
XFILLER_129_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13597_ _13597_/A _13597_/B vssd1 vssd1 vccd1 vccd1 _13598_/B sky130_fd_sc_hd__nor2_1
XFILLER_8_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15336_ _15337_/A _15337_/B vssd1 vssd1 vccd1 vccd1 _15336_/Y sky130_fd_sc_hd__nand2_1
X_12548_ _13831_/S _12548_/B vssd1 vssd1 vccd1 vccd1 _12548_/Y sky130_fd_sc_hd__nor2_1
XFILLER_117_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15267_ _16127_/A _16536_/A _16533_/A _15726_/A vssd1 vssd1 vccd1 vccd1 _15268_/B
+ sky130_fd_sc_hd__a22o_1
X_12479_ _12481_/A _12481_/B _12481_/C vssd1 vssd1 vccd1 vccd1 _12479_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA_2 _17479_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17006_ _17007_/A _17007_/B vssd1 vssd1 vccd1 vccd1 _17093_/A sky130_fd_sc_hd__or2_1
X_14218_ _14218_/A _14218_/B _14218_/C vssd1 vssd1 vccd1 vccd1 _14219_/B sky130_fd_sc_hd__or3_1
XFILLER_172_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_910 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15198_ _15147_/A _11789_/X _15393_/B vssd1 vssd1 vccd1 vccd1 _15198_/X sky130_fd_sc_hd__a21o_1
X_14149_ _14150_/A _14150_/B _14150_/C vssd1 vssd1 vccd1 vccd1 _14151_/A sky130_fd_sc_hd__o21a_1
Xfanout509 _11370_/A vssd1 vssd1 vccd1 vccd1 _15396_/A sky130_fd_sc_hd__buf_4
XFILLER_113_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_987 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_423 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09690_ _10366_/A _09985_/D _09552_/A _09550_/Y vssd1 vssd1 vccd1 vccd1 _09696_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_6_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_562 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_18 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09124_ _17423_/A _17421_/A _09172_/B _09502_/B vssd1 vssd1 vccd1 vccd1 _09167_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_157_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09055_ _09055_/A _09055_/B _09055_/C vssd1 vssd1 vccd1 vccd1 _09055_/Y sky130_fd_sc_hd__nand3_1
XFILLER_135_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09957_ _09957_/A _09957_/B vssd1 vssd1 vccd1 vccd1 _09960_/B sky130_fd_sc_hd__and2_1
XFILLER_131_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08908_ _08908_/A _08908_/B vssd1 vssd1 vccd1 vccd1 _08910_/C sky130_fd_sc_hd__or2_1
XFILLER_131_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09888_ _09869_/X _09885_/A _09887_/Y _09765_/X vssd1 vssd1 vccd1 vccd1 _09912_/A
+ sky130_fd_sc_hd__a211oi_1
XFILLER_85_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08839_ _08862_/B _08839_/B vssd1 vssd1 vccd1 vccd1 _08845_/A sky130_fd_sc_hd__nor2_1
XFILLER_58_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11850_ _11651_/A _11675_/B _11675_/C vssd1 vssd1 vccd1 vccd1 _11851_/B sky130_fd_sc_hd__o21ai_1
XTAP_2735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10801_ _11115_/A _10963_/C _10800_/C vssd1 vssd1 vccd1 vccd1 _10802_/B sky130_fd_sc_hd__a21oi_1
XTAP_2757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11781_ _12016_/B _11781_/B vssd1 vssd1 vccd1 vccd1 _14837_/A sky130_fd_sc_hd__and2_1
XFILLER_81_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13520_ _14757_/S _14735_/A1 _12548_/B _13519_/Y _14636_/A vssd1 vssd1 vccd1 vccd1
+ _13520_/X sky130_fd_sc_hd__a311o_1
XFILLER_82_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10732_ _10662_/A _10662_/B _10662_/C vssd1 vssd1 vccd1 vccd1 _10732_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_159_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_367 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13451_ _13451_/A _13569_/A vssd1 vssd1 vccd1 vccd1 _13453_/C sky130_fd_sc_hd__nor2_1
XFILLER_51_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10663_ _10651_/Y _10662_/X _10670_/A _10636_/Y vssd1 vssd1 vccd1 vccd1 _10670_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_9_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12402_ _11849_/A _12396_/X _12401_/X _16653_/A vssd1 vssd1 vccd1 vccd1 _12403_/B
+ sky130_fd_sc_hd__a22o_1
X_16170_ _16170_/A _16170_/B vssd1 vssd1 vccd1 vccd1 _16172_/A sky130_fd_sc_hd__nand2_1
X_10594_ _11027_/B _10594_/B vssd1 vssd1 vccd1 vccd1 _10595_/B sky130_fd_sc_hd__nand2_1
X_13382_ _13504_/A _13380_/X _13221_/A _13224_/A vssd1 vssd1 vccd1 vccd1 _13382_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_167_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15121_ _12054_/A _10036_/D _10897_/C _10545_/C vssd1 vssd1 vccd1 vccd1 _15121_/X
+ sky130_fd_sc_hd__a211o_1
X_12333_ _12333_/A _12333_/B vssd1 vssd1 vccd1 vccd1 _12334_/C sky130_fd_sc_hd__xnor2_1
XFILLER_5_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15052_ _11675_/C _11655_/A _11676_/A vssd1 vssd1 vccd1 vccd1 _15052_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_154_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12264_ _12437_/A _12265_/B _12265_/C vssd1 vssd1 vccd1 vccd1 _12266_/A sky130_fd_sc_hd__a21o_1
XFILLER_135_770 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14003_ _14176_/A _14366_/B _14002_/C vssd1 vssd1 vccd1 vccd1 _14004_/B sky130_fd_sc_hd__a21o_1
X_11215_ _11216_/A _11216_/B vssd1 vssd1 vccd1 vccd1 _11215_/Y sky130_fd_sc_hd__nor2_1
X_12195_ _11998_/A _11997_/Y _12360_/B _12194_/X vssd1 vssd1 vccd1 vccd1 _12198_/A
+ sky130_fd_sc_hd__o211a_1
Xoutput72 _17476_/Q vssd1 vssd1 vccd1 vccd1 leds[10] sky130_fd_sc_hd__clkbuf_1
XFILLER_110_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11146_ _11146_/A _11146_/B vssd1 vssd1 vccd1 vccd1 _11148_/B sky130_fd_sc_hd__and2_1
Xoutput83 _17542_/Q vssd1 vssd1 vccd1 vccd1 o_wb_ack sky130_fd_sc_hd__clkbuf_1
XFILLER_95_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput94 _17453_/Q vssd1 vssd1 vccd1 vccd1 o_wb_data[19] sky130_fd_sc_hd__clkbuf_1
XFILLER_96_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11077_ _11077_/A _11110_/A _11077_/C vssd1 vssd1 vccd1 vccd1 _11080_/B sky130_fd_sc_hd__or3_2
X_15954_ _15954_/A _15954_/B vssd1 vssd1 vccd1 vccd1 _15964_/A sky130_fd_sc_hd__and2_1
X_14905_ _15208_/C _15208_/D _14905_/C _14905_/D vssd1 vssd1 vccd1 vccd1 _14905_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_37_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10028_ _10028_/A _10028_/B vssd1 vssd1 vccd1 vccd1 _10029_/C sky130_fd_sc_hd__nor2_1
XFILLER_64_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15885_ _15788_/Y _15790_/X _15787_/X vssd1 vssd1 vccd1 vccd1 _15885_/Y sky130_fd_sc_hd__a21boi_2
X_14836_ _17063_/A _14836_/B _14933_/B vssd1 vssd1 vccd1 vccd1 _14836_/Y sky130_fd_sc_hd__nand3_1
XFILLER_64_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17555_ fanout940/X _17555_/D vssd1 vssd1 vccd1 vccd1 _17555_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14767_ _16965_/C _16974_/A vssd1 vssd1 vccd1 vccd1 _14767_/Y sky130_fd_sc_hd__nor2_1
XFILLER_32_610 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11979_ _17415_/A _12338_/D vssd1 vssd1 vccd1 vccd1 _11980_/B sky130_fd_sc_hd__nand2_1
X_16506_ _16503_/A _16670_/A _16504_/Y _16505_/X vssd1 vssd1 vccd1 vccd1 _16507_/B
+ sky130_fd_sc_hd__o211a_1
X_13718_ _13718_/A _13718_/B vssd1 vssd1 vccd1 vccd1 _13720_/B sky130_fd_sc_hd__nand2_1
X_17486_ fanout948/X _17486_/D vssd1 vssd1 vccd1 vccd1 _17486_/Q sky130_fd_sc_hd__dfxtp_4
X_14698_ _14698_/A _14698_/B vssd1 vssd1 vccd1 vccd1 _14699_/B sky130_fd_sc_hd__nand2_1
XFILLER_108_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16437_ _16437_/A _16437_/B vssd1 vssd1 vccd1 vccd1 _16439_/B sky130_fd_sc_hd__xnor2_1
XFILLER_72_90 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13649_ _13749_/B _13648_/B _13648_/C vssd1 vssd1 vccd1 vccd1 _13650_/B sky130_fd_sc_hd__a21o_1
XFILLER_158_840 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16368_ _16273_/A _16273_/B _16256_/X vssd1 vssd1 vccd1 vccd1 _16369_/B sky130_fd_sc_hd__a21o_1
XFILLER_173_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15319_ _15039_/X _15057_/X _15059_/Y _15061_/Y _15312_/S _15901_/S vssd1 vssd1 vccd1
+ vccd1 _15319_/X sky130_fd_sc_hd__mux4_1
XFILLER_117_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16299_ _16394_/A _16299_/B vssd1 vssd1 vccd1 vccd1 _16301_/A sky130_fd_sc_hd__nand2_1
XFILLER_173_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_386 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout306 _14733_/S vssd1 vssd1 vccd1 vccd1 _13625_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_113_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout317 _17609_/Q vssd1 vssd1 vccd1 vccd1 _17476_/D sky130_fd_sc_hd__buf_6
X_09811_ _09811_/A _09811_/B vssd1 vssd1 vccd1 vccd1 _09813_/B sky130_fd_sc_hd__xor2_1
XFILLER_141_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout328 _08988_/B vssd1 vssd1 vccd1 vccd1 _14050_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_115_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout339 _11922_/A vssd1 vssd1 vccd1 vccd1 _17421_/A sky130_fd_sc_hd__buf_4
XFILLER_87_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09742_ _09812_/B vssd1 vssd1 vccd1 vccd1 _09769_/A sky130_fd_sc_hd__inv_2
XFILLER_100_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09673_ _10559_/A _12340_/B _09386_/B _09384_/X vssd1 vssd1 vccd1 vccd1 _09675_/B
+ sky130_fd_sc_hd__a31oi_1
XFILLER_36_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_383 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09107_ _17421_/A _09362_/D vssd1 vssd1 vccd1 vccd1 _09108_/B sky130_fd_sc_hd__nand2_1
XFILLER_108_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09038_ _09039_/A _09039_/B vssd1 vssd1 vccd1 vccd1 _09055_/A sky130_fd_sc_hd__nand2b_1
XFILLER_136_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11000_ _10999_/A _10999_/B _10999_/C vssd1 vssd1 vccd1 vccd1 _11000_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_105_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout840 _11387_/B vssd1 vssd1 vccd1 vccd1 _10799_/B sky130_fd_sc_hd__buf_4
XFILLER_77_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout851 _14849_/A vssd1 vssd1 vccd1 vccd1 _14788_/B sky130_fd_sc_hd__buf_4
Xfanout862 _12295_/D vssd1 vssd1 vccd1 vccd1 _10359_/B sky130_fd_sc_hd__buf_4
Xfanout873 fanout874/X vssd1 vssd1 vccd1 vccd1 _10479_/B sky130_fd_sc_hd__buf_4
Xfanout884 _11427_/C vssd1 vssd1 vccd1 vccd1 _10594_/B sky130_fd_sc_hd__clkbuf_4
XTAP_3200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout895 _15003_/B vssd1 vssd1 vccd1 vccd1 _09172_/B sky130_fd_sc_hd__clkbuf_4
X_12951_ _13903_/A _13866_/C _12950_/C vssd1 vssd1 vccd1 vccd1 _12952_/B sky130_fd_sc_hd__a21o_1
XTAP_3211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11902_ _17381_/A _11902_/B vssd1 vssd1 vccd1 vccd1 _11903_/B sky130_fd_sc_hd__nand2_1
XFILLER_45_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15670_ _15671_/A _15671_/B vssd1 vssd1 vccd1 vccd1 _15764_/A sky130_fd_sc_hd__nand2_1
XFILLER_46_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12882_ _13040_/B _12882_/B vssd1 vssd1 vccd1 vccd1 _12884_/B sky130_fd_sc_hd__and2b_1
XTAP_3266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14621_ _14621_/A _14621_/B _14621_/C vssd1 vssd1 vccd1 vccd1 _14622_/B sky130_fd_sc_hd__and3_1
XTAP_2543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11833_ _11827_/X _11832_/X _17367_/A vssd1 vssd1 vccd1 vccd1 _11833_/X sky130_fd_sc_hd__mux2_1
XTAP_2554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17340_ _09319_/C _17360_/A2 _17339_/X _17406_/C1 vssd1 vssd1 vccd1 vccd1 _17499_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14552_ _14680_/A _14599_/B _14708_/D _14641_/C vssd1 vssd1 vccd1 vccd1 _14553_/B
+ sky130_fd_sc_hd__and4_1
X_11764_ _16727_/B _16795_/A _11762_/X _11763_/Y vssd1 vssd1 vccd1 vccd1 _11764_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_60_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_142 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13503_ _13503_/A _13503_/B vssd1 vssd1 vccd1 vccd1 _13506_/A sky130_fd_sc_hd__xnor2_1
XTAP_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10715_ _10715_/A _10715_/B _10715_/C vssd1 vssd1 vccd1 vccd1 _10715_/Y sky130_fd_sc_hd__nand3_1
XTAP_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17271_ _17567_/Q _17292_/B vssd1 vssd1 vccd1 vccd1 _17271_/X sky130_fd_sc_hd__and2_1
XFILLER_159_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14483_ _14842_/A1 _14481_/X _14482_/X vssd1 vssd1 vccd1 vccd1 _14483_/Y sky130_fd_sc_hd__a21oi_2
X_11695_ _11691_/Y _11693_/Y _11694_/X _11672_/Y vssd1 vssd1 vccd1 vccd1 _15447_/A
+ sky130_fd_sc_hd__o211a_1
X_16222_ _16212_/Y _16213_/X _16221_/X vssd1 vssd1 vccd1 vccd1 _16222_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_146_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13434_ _13434_/A _13434_/B _13551_/D _13434_/D vssd1 vssd1 vccd1 vccd1 _13586_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_9_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10646_ _10851_/B _10745_/D _10786_/B _11122_/A vssd1 vssd1 vccd1 vccd1 _10646_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_167_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16153_ _16153_/A _16153_/B vssd1 vssd1 vccd1 vccd1 _16155_/B sky130_fd_sc_hd__xor2_1
XFILLER_158_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13365_ _13366_/A _13366_/B vssd1 vssd1 vccd1 vccd1 _13365_/Y sky130_fd_sc_hd__nand2b_1
X_10577_ _10463_/B _10471_/X _10573_/X _10575_/Y vssd1 vssd1 vccd1 vccd1 _10577_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_154_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15104_ _15715_/B _15103_/X _15116_/A vssd1 vssd1 vccd1 vccd1 _15104_/X sky130_fd_sc_hd__mux2_1
XFILLER_170_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12316_ _12316_/A _12316_/B _12316_/C vssd1 vssd1 vccd1 vccd1 _12358_/B sky130_fd_sc_hd__nand3_1
X_16084_ _16084_/A _16084_/B _16082_/X vssd1 vssd1 vccd1 vccd1 _16085_/B sky130_fd_sc_hd__or3b_1
XFILLER_5_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13296_ _13170_/A _13172_/B _13170_/B vssd1 vssd1 vccd1 vccd1 _13306_/A sky130_fd_sc_hd__o21ba_1
XFILLER_154_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15035_ _16011_/C _15034_/Y _15312_/S vssd1 vssd1 vccd1 vccd1 _15627_/B sky130_fd_sc_hd__mux2_1
XFILLER_114_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12247_ _12247_/A _12247_/B vssd1 vssd1 vccd1 vccd1 _12248_/B sky130_fd_sc_hd__nand2_1
XFILLER_68_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12178_ _12179_/A _12179_/B _12179_/C vssd1 vssd1 vccd1 vccd1 _12180_/A sky130_fd_sc_hd__o21a_1
XFILLER_122_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11129_ _11130_/B _11130_/C _11130_/A vssd1 vssd1 vccd1 vccd1 _11139_/A sky130_fd_sc_hd__a21o_1
XFILLER_1_591 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16986_ _16986_/A _16986_/B vssd1 vssd1 vccd1 vccd1 _16991_/B sky130_fd_sc_hd__xnor2_1
XFILLER_49_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15937_ _15937_/A _15937_/B vssd1 vssd1 vccd1 vccd1 _15939_/B sky130_fd_sc_hd__xor2_1
XFILLER_49_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15868_ _15868_/A _15868_/B vssd1 vssd1 vccd1 vccd1 _15871_/A sky130_fd_sc_hd__or2_1
XFILLER_37_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17607_ fanout939/X _17607_/D vssd1 vssd1 vccd1 vccd1 _17607_/Q sky130_fd_sc_hd__dfxtp_4
X_14819_ _16649_/B _16649_/C _16649_/A vssd1 vssd1 vccd1 vccd1 _16730_/A sky130_fd_sc_hd__a21bo_1
XFILLER_91_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_470 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15799_ _15797_/Y _15798_/Y _16111_/A vssd1 vssd1 vccd1 vccd1 _15799_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_51_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17538_ fanout947/X _17538_/D vssd1 vssd1 vccd1 vccd1 _17538_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_51_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_451 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17469_ fanout955/X _17469_/D vssd1 vssd1 vccd1 vccd1 _17469_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_526 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout125 _17244_/B vssd1 vssd1 vccd1 vccd1 _17289_/B sky130_fd_sc_hd__clkbuf_2
Xfanout136 _15199_/Y vssd1 vssd1 vccd1 vccd1 _16536_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_141_592 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout147 _14969_/Y vssd1 vssd1 vccd1 vccd1 _16127_/A sky130_fd_sc_hd__buf_2
XFILLER_59_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_423 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout158 _17371_/B vssd1 vssd1 vccd1 vccd1 _17424_/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_87_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout169 _16987_/B vssd1 vssd1 vccd1 vccd1 _17043_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_41_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09725_ _09725_/A _09725_/B _09725_/C vssd1 vssd1 vccd1 vccd1 _09725_/Y sky130_fd_sc_hd__nand3_1
XFILLER_55_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_690 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09656_ _09656_/A _09656_/B _09656_/C vssd1 vssd1 vccd1 vccd1 _09788_/A sky130_fd_sc_hd__or3_1
XFILLER_82_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09587_ _09587_/A _09727_/A vssd1 vssd1 vccd1 vccd1 _09589_/B sky130_fd_sc_hd__nor2_1
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10500_ _10485_/X _10499_/A _10384_/X _10475_/Y vssd1 vssd1 vccd1 vccd1 _10519_/A
+ sky130_fd_sc_hd__a211oi_4
X_11480_ _11518_/A _11518_/B _14850_/A _15238_/A vssd1 vssd1 vccd1 vccd1 _11484_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_7_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10431_ _10753_/A _10431_/B _14956_/A vssd1 vssd1 vccd1 vccd1 _10434_/A sky130_fd_sc_hd__and3_1
XFILLER_6_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13150_ _13846_/A _14063_/C vssd1 vssd1 vccd1 vccd1 _13151_/B sky130_fd_sc_hd__nand2_1
XFILLER_164_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10362_ _10374_/A _10362_/B vssd1 vssd1 vccd1 vccd1 _10364_/B sky130_fd_sc_hd__or2_1
XFILLER_152_835 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12101_ _11895_/B _12447_/B _12445_/C _17379_/A vssd1 vssd1 vccd1 vccd1 _12103_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_151_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13081_ _13897_/A _13208_/C vssd1 vssd1 vccd1 vccd1 _13083_/C sky130_fd_sc_hd__nand2_1
XFILLER_88_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10293_ _10293_/A _10399_/A vssd1 vssd1 vccd1 vccd1 _10301_/A sky130_fd_sc_hd__nor2_1
XFILLER_2_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12032_ _12050_/S _17134_/B vssd1 vssd1 vccd1 vccd1 _12032_/Y sky130_fd_sc_hd__nor2_1
XFILLER_88_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16840_ _16841_/A _16841_/B vssd1 vssd1 vccd1 vccd1 _16906_/A sky130_fd_sc_hd__nand2b_1
XFILLER_77_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout670 _17503_/Q vssd1 vssd1 vccd1 vccd1 _14865_/B sky130_fd_sc_hd__clkbuf_4
Xfanout681 _17502_/Q vssd1 vssd1 vccd1 vccd1 _08860_/B sky130_fd_sc_hd__buf_2
XFILLER_77_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16771_ _16771_/A _16771_/B vssd1 vssd1 vccd1 vccd1 _16775_/A sky130_fd_sc_hd__and2_1
Xfanout692 fanout699/X vssd1 vssd1 vccd1 vccd1 _13348_/B sky130_fd_sc_hd__buf_2
X_13983_ _13878_/A _13880_/B _13878_/B vssd1 vssd1 vccd1 vccd1 _13985_/B sky130_fd_sc_hd__o21ba_1
XFILLER_77_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15722_ _15206_/A _16977_/A _15721_/X vssd1 vssd1 vccd1 vccd1 _17554_/D sky130_fd_sc_hd__o21a_1
XTAP_3030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12934_ _12933_/A _12933_/B _12933_/C vssd1 vssd1 vccd1 vccd1 _12935_/B sky130_fd_sc_hd__o21a_1
XTAP_3041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15653_ _15742_/A _15742_/B vssd1 vssd1 vccd1 vccd1 _15654_/B sky130_fd_sc_hd__and2_1
XFILLER_160_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12865_ _12390_/X _12393_/B _12865_/S vssd1 vssd1 vccd1 vccd1 _12866_/B sky130_fd_sc_hd__mux2_1
XTAP_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_94 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14604_ _14553_/A _14555_/B _14553_/B vssd1 vssd1 vccd1 vccd1 _14606_/B sky130_fd_sc_hd__o21ba_1
XTAP_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11816_ _14981_/A _14978_/B _11837_/A vssd1 vssd1 vccd1 vccd1 _11816_/Y sky130_fd_sc_hd__o21ai_1
XTAP_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15584_ _15584_/A _15584_/B vssd1 vssd1 vccd1 vccd1 _15685_/B sky130_fd_sc_hd__xnor2_1
XFILLER_18_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12796_ _12796_/A _12796_/B vssd1 vssd1 vccd1 vccd1 _12798_/C sky130_fd_sc_hd__xor2_1
XTAP_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_412 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17323_ input40/X _17359_/B _17359_/C vssd1 vssd1 vccd1 vccd1 _17323_/X sky130_fd_sc_hd__or3_1
XTAP_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14535_ _14414_/A _14475_/A _14533_/B vssd1 vssd1 vccd1 vccd1 _14535_/Y sky130_fd_sc_hd__o21ai_1
XTAP_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11747_ _11758_/A _11747_/B vssd1 vssd1 vccd1 vccd1 _11748_/B sky130_fd_sc_hd__or2_1
XTAP_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17254_ _17452_/Q _17290_/A2 _17252_/X _17253_/X _17293_/C1 vssd1 vssd1 vccd1 vccd1
+ _17452_/D sky130_fd_sc_hd__o221a_1
X_14466_ _14466_/A _14466_/B vssd1 vssd1 vccd1 vccd1 _14524_/B sky130_fd_sc_hd__and2_1
XFILLER_128_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11678_ _11678_/A _11678_/B vssd1 vssd1 vccd1 vccd1 _11679_/B sky130_fd_sc_hd__and2_1
XFILLER_128_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16205_ _16292_/B _16205_/B vssd1 vssd1 vccd1 vccd1 _16205_/X sky130_fd_sc_hd__or2_1
X_13417_ _13417_/A _13417_/B _13417_/C vssd1 vssd1 vccd1 vccd1 _13418_/B sky130_fd_sc_hd__or3_1
X_10629_ _10614_/X _10615_/Y _10623_/X _10627_/X vssd1 vssd1 vccd1 vccd1 _10632_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_127_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17185_ input25/X _17362_/A input1/X _17428_/C vssd1 vssd1 vccd1 vccd1 _17185_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_127_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14397_ _14316_/A _14332_/X _14395_/Y _14396_/X vssd1 vssd1 vccd1 vccd1 _14466_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_128_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16136_ _16136_/A _16136_/B _16136_/C vssd1 vssd1 vccd1 vccd1 _16250_/A sky130_fd_sc_hd__and3_1
XFILLER_128_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13348_ _13578_/A _13348_/B vssd1 vssd1 vccd1 vccd1 _13349_/B sky130_fd_sc_hd__nand2_1
XFILLER_127_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16067_ _15853_/B _15955_/Y _15960_/A _15960_/B vssd1 vssd1 vccd1 vccd1 _16068_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_5_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13279_ _13632_/A _13735_/B _13522_/D _14063_/C vssd1 vssd1 vccd1 vccd1 _13280_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_170_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15018_ _15617_/A _14967_/C _14967_/D _14900_/X _14877_/Y vssd1 vssd1 vccd1 vccd1
+ _15018_/X sky130_fd_sc_hd__o32a_1
XFILLER_97_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16969_ _16969_/A _16969_/B vssd1 vssd1 vccd1 vccd1 _16969_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_49_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09510_ _10560_/A _09843_/C _09382_/C vssd1 vssd1 vccd1 vccd1 _09511_/B sky130_fd_sc_hd__a21oi_1
XFILLER_65_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09441_ _09441_/A _09441_/B _09441_/C vssd1 vssd1 vccd1 vccd1 _09441_/Y sky130_fd_sc_hd__nand3_1
XFILLER_80_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09372_ _17407_/A _09555_/D _09209_/C vssd1 vssd1 vccd1 vccd1 _09373_/B sky130_fd_sc_hd__a21oi_1
XFILLER_33_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_1026 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_966 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09708_ _09709_/A _09709_/B vssd1 vssd1 vccd1 vccd1 _09725_/A sky130_fd_sc_hd__nand2b_1
X_10980_ _10745_/C _10932_/B _10936_/B _10935_/A vssd1 vssd1 vccd1 vccd1 _10987_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_74_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xwb_buttons_leds_966 vssd1 vssd1 vccd1 vccd1 wb_buttons_leds_966/HI led_enb[8] sky130_fd_sc_hd__conb_1
XFILLER_167_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09639_ _09640_/A _09638_/Y _09639_/C _10203_/B vssd1 vssd1 vccd1 vccd1 _09795_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_130_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12650_ _12649_/B _12650_/B vssd1 vssd1 vccd1 vccd1 _12651_/B sky130_fd_sc_hd__nand2b_1
XFILLER_128_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11601_ _11639_/A _11639_/B vssd1 vssd1 vccd1 vccd1 _11603_/B sky130_fd_sc_hd__nand2_1
XFILLER_130_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12581_ _12581_/A _12581_/B vssd1 vssd1 vccd1 vccd1 _12583_/B sky130_fd_sc_hd__xnor2_1
XFILLER_23_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14320_ _14387_/A _14383_/B _14321_/C vssd1 vssd1 vccd1 vccd1 _14324_/A sky130_fd_sc_hd__a21oi_1
X_11532_ _11532_/A _11532_/B _11574_/A vssd1 vssd1 vccd1 vccd1 _11538_/A sky130_fd_sc_hd__nor3b_1
XFILLER_12_966 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14251_ _14252_/A _14252_/B _14252_/C vssd1 vssd1 vccd1 vccd1 _14253_/A sky130_fd_sc_hd__a21oi_1
X_11463_ _11416_/B _11413_/B _11413_/C vssd1 vssd1 vccd1 vccd1 _11464_/B sky130_fd_sc_hd__o21a_1
XFILLER_139_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13202_ _13332_/A _13202_/B _13202_/C vssd1 vssd1 vccd1 vccd1 _13203_/A sky130_fd_sc_hd__and3_1
XFILLER_7_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10414_ _10415_/A _10413_/Y _14788_/A _10745_/D vssd1 vssd1 vccd1 vccd1 _10513_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_125_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14182_ _14254_/A _14181_/B _14181_/C vssd1 vssd1 vccd1 vccd1 _14184_/C sky130_fd_sc_hd__a21o_1
X_11394_ _11453_/A _11394_/B vssd1 vssd1 vccd1 vccd1 _11396_/B sky130_fd_sc_hd__and2_1
XFILLER_99_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_1014 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13133_ _12993_/X _12999_/A _13264_/B _13132_/X vssd1 vssd1 vccd1 vccd1 _13137_/A
+ sky130_fd_sc_hd__a211o_1
X_10345_ _10345_/A _10581_/A vssd1 vssd1 vccd1 vccd1 _10349_/B sky130_fd_sc_hd__nor2_1
XFILLER_3_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13064_ _13065_/A _13065_/B _13065_/C vssd1 vssd1 vccd1 vccd1 _13075_/A sky130_fd_sc_hd__a21o_1
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10276_ _10276_/A _10276_/B vssd1 vssd1 vccd1 vccd1 _10387_/A sky130_fd_sc_hd__xor2_1
XFILLER_78_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12015_ _09679_/A _09826_/A _09679_/B vssd1 vssd1 vccd1 vccd1 _12015_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_39_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16823_ _16897_/A _16823_/B vssd1 vssd1 vccd1 vccd1 _16832_/A sky130_fd_sc_hd__or2_1
XFILLER_93_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16754_ _16680_/X _16684_/B _16682_/B vssd1 vssd1 vccd1 vccd1 _16764_/B sky130_fd_sc_hd__o21a_1
X_13966_ _13966_/A _14050_/B _13966_/C _13966_/D vssd1 vssd1 vccd1 vccd1 _13967_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_111_1042 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12917_ _13065_/A _12918_/B _12918_/C vssd1 vssd1 vccd1 vccd1 _12919_/A sky130_fd_sc_hd__a21o_1
X_15705_ _15705_/A _15705_/B _15705_/C vssd1 vssd1 vccd1 vccd1 _15705_/Y sky130_fd_sc_hd__nand3_1
X_16685_ _16686_/A _16686_/B _16684_/Y vssd1 vssd1 vccd1 vccd1 _16685_/X sky130_fd_sc_hd__o21ba_1
X_13897_ _13897_/A _14485_/D vssd1 vssd1 vccd1 vccd1 _13898_/B sky130_fd_sc_hd__nand2_1
XFILLER_73_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12848_ _12212_/X _12217_/B _12848_/S vssd1 vssd1 vccd1 vccd1 _12849_/B sky130_fd_sc_hd__mux2_1
XTAP_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15636_ _15636_/A vssd1 vssd1 vccd1 vccd1 _17553_/D sky130_fd_sc_hd__inv_2
XFILLER_22_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15567_ _15567_/A _15666_/A vssd1 vssd1 vccd1 vccd1 _15568_/B sky130_fd_sc_hd__nand2_1
X_12779_ _12779_/A _12779_/B vssd1 vssd1 vccd1 vccd1 _12780_/B sky130_fd_sc_hd__nor2_1
XTAP_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17306_ _17306_/A1 _17308_/A2 _17305_/X _17358_/C1 vssd1 vssd1 vccd1 vccd1 _17482_/D
+ sky130_fd_sc_hd__o211a_1
X_14518_ _14518_/A _14518_/B _14518_/C vssd1 vssd1 vccd1 vccd1 _14519_/C sky130_fd_sc_hd__nand3_1
XFILLER_9_86 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15498_ _15498_/A _15498_/B vssd1 vssd1 vccd1 vccd1 _15499_/B sky130_fd_sc_hd__xor2_1
XFILLER_30_774 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17237_ _17588_/Q _17291_/A2 _17291_/B1 vssd1 vssd1 vccd1 vccd1 _17237_/X sky130_fd_sc_hd__a21o_1
X_14449_ _16913_/C _14450_/B vssd1 vssd1 vccd1 vccd1 _14509_/B sky130_fd_sc_hd__nand2_1
XFILLER_162_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17168_ _17167_/A _17167_/B _17167_/C vssd1 vssd1 vccd1 vccd1 _17168_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_116_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16119_ _16112_/B _17162_/A2 _16580_/B1 _16114_/A _17162_/C1 vssd1 vssd1 vccd1 vccd1
+ _16119_/X sky130_fd_sc_hd__a221o_1
XFILLER_127_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17099_ _17099_/A vssd1 vssd1 vccd1 vccd1 _17099_/Y sky130_fd_sc_hd__inv_2
X_09990_ _10106_/A _10106_/B vssd1 vssd1 vccd1 vccd1 _10004_/C sky130_fd_sc_hd__nand2_1
XFILLER_143_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08941_ _08941_/A _08941_/B vssd1 vssd1 vccd1 vccd1 _08943_/A sky130_fd_sc_hd__nor2_1
XFILLER_142_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08872_ _08874_/A _08874_/B _08873_/C _08873_/D vssd1 vssd1 vccd1 vccd1 _08872_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_85_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_936 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09424_ _11790_/A _15898_/A vssd1 vssd1 vccd1 vccd1 _09424_/X sky130_fd_sc_hd__and2_1
XFILLER_52_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09355_ _09355_/A _09355_/B vssd1 vssd1 vccd1 vccd1 _09479_/B sky130_fd_sc_hd__xnor2_1
XFILLER_100_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09286_ _17081_/B _16990_/A _09285_/X vssd1 vssd1 vccd1 vccd1 _09421_/B sky130_fd_sc_hd__o21ai_1
XFILLER_138_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10130_ _10128_/B _10251_/B _10128_/A vssd1 vssd1 vccd1 vccd1 _10132_/B sky130_fd_sc_hd__o21ba_1
XFILLER_79_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10061_ _10061_/A _10061_/B vssd1 vssd1 vccd1 vccd1 _10069_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13820_ _13820_/A _13820_/B vssd1 vssd1 vccd1 vccd1 _13823_/A sky130_fd_sc_hd__xor2_2
XFILLER_47_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13751_ _13751_/A _13751_/B vssd1 vssd1 vccd1 vccd1 _13754_/A sky130_fd_sc_hd__xnor2_1
XFILLER_44_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10963_ _10963_/A _10963_/B _10963_/C _11117_/D vssd1 vssd1 vccd1 vccd1 _10965_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_16_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12702_ _12027_/X _12034_/X _15384_/S vssd1 vssd1 vccd1 vccd1 _12702_/X sky130_fd_sc_hd__mux2_1
X_16470_ _16470_/A _16470_/B _16470_/C vssd1 vssd1 vccd1 vccd1 _16563_/B sky130_fd_sc_hd__and3_1
X_13682_ _13582_/A _13584_/B _13582_/B vssd1 vssd1 vccd1 vccd1 _13683_/B sky130_fd_sc_hd__o21ba_1
X_10894_ _10881_/Y _11112_/A _10895_/A _10864_/Y vssd1 vssd1 vccd1 vccd1 _11080_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_31_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15421_ _15422_/A _15422_/B vssd1 vssd1 vccd1 vccd1 _15507_/A sky130_fd_sc_hd__and2b_1
X_12633_ _12630_/X _12631_/Y _12481_/A _12481_/Y vssd1 vssd1 vccd1 vccd1 _12676_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_169_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15352_ _15352_/A _15352_/B vssd1 vssd1 vccd1 vccd1 _15359_/A sky130_fd_sc_hd__xnor2_1
X_12564_ _12722_/B _13348_/B _12871_/B _12722_/A vssd1 vssd1 vccd1 vccd1 _12566_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_11_251 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14303_ _14554_/A _14366_/B vssd1 vssd1 vccd1 vccd1 _14304_/B sky130_fd_sc_hd__nand2_1
X_11515_ _11520_/C _11518_/C _11484_/B _11481_/Y vssd1 vssd1 vccd1 vccd1 _11522_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_141_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15283_ _15283_/A _15283_/B vssd1 vssd1 vccd1 vccd1 _15285_/B sky130_fd_sc_hd__xnor2_1
X_12495_ _12795_/A _12942_/D vssd1 vssd1 vccd1 vccd1 _12496_/B sky130_fd_sc_hd__nand2_1
X_17022_ _17018_/A _17066_/A _17066_/B _17156_/B vssd1 vssd1 vccd1 vccd1 _17022_/X
+ sky130_fd_sc_hd__a31o_1
X_14234_ _14235_/A _14235_/B vssd1 vssd1 vccd1 vccd1 _14315_/A sky130_fd_sc_hd__or2_1
X_11446_ _11396_/X _11421_/Y _11444_/A _11444_/Y vssd1 vssd1 vccd1 vccd1 _11449_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_50_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14165_ _14165_/A _14165_/B vssd1 vssd1 vccd1 vccd1 _14185_/A sky130_fd_sc_hd__xnor2_1
X_11377_ _11427_/A _11553_/A _11563_/D _11561_/D vssd1 vssd1 vccd1 vccd1 _11380_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_140_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13116_ _13117_/A _13117_/B _13117_/C vssd1 vssd1 vccd1 vccd1 _13118_/A sky130_fd_sc_hd__a21o_1
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10328_ _10329_/B _10329_/C vssd1 vssd1 vccd1 vccd1 _10450_/B sky130_fd_sc_hd__and2_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14096_ _14200_/B _14096_/B vssd1 vssd1 vccd1 vccd1 _14098_/B sky130_fd_sc_hd__or2_1
XFILLER_124_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13047_ _13047_/A _13047_/B vssd1 vssd1 vccd1 vccd1 _13049_/C sky130_fd_sc_hd__nand2_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10259_ _10260_/B _10260_/A vssd1 vssd1 vccd1 vccd1 _10267_/B sky130_fd_sc_hd__nand2b_1
XFILLER_59_91 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_638 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16806_ _16789_/A _16806_/A2 _16805_/X vssd1 vssd1 vccd1 vccd1 _17566_/D sky130_fd_sc_hd__a21oi_1
XFILLER_54_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14998_ _15100_/A _14998_/B vssd1 vssd1 vccd1 vccd1 _14998_/Y sky130_fd_sc_hd__nand2_1
XFILLER_47_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16737_ _16485_/A _16730_/Y _16732_/X _16736_/X vssd1 vssd1 vccd1 vccd1 _16737_/X
+ sky130_fd_sc_hd__a211o_1
X_13949_ _13949_/A _13949_/B vssd1 vssd1 vccd1 vccd1 _13951_/A sky130_fd_sc_hd__nor2_1
XFILLER_81_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16668_ _16670_/A _16670_/B _16670_/C vssd1 vssd1 vccd1 vccd1 _16671_/A sky130_fd_sc_hd__a21oi_1
XFILLER_22_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15619_ _15453_/B _15453_/C _15529_/Y _15449_/Y vssd1 vssd1 vccd1 vccd1 _15620_/B
+ sky130_fd_sc_hd__a211o_1
X_16599_ _16600_/A _16600_/B vssd1 vssd1 vccd1 vccd1 _16601_/A sky130_fd_sc_hd__nand2_1
XFILLER_50_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09140_ _09106_/A _09108_/B _09106_/B vssd1 vssd1 vccd1 vccd1 _09148_/A sky130_fd_sc_hd__o21ba_1
XFILLER_148_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09071_ _09071_/A _09071_/B _09071_/C vssd1 vssd1 vccd1 vccd1 _09259_/A sky130_fd_sc_hd__nor3_1
XFILLER_136_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09973_ _09973_/A _09973_/B vssd1 vssd1 vccd1 vccd1 _10059_/B sky130_fd_sc_hd__and2_1
XFILLER_103_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08924_ _09052_/A _09052_/B vssd1 vssd1 vccd1 vccd1 _09053_/A sky130_fd_sc_hd__and2_1
XFILLER_162_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_711 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08855_ _09321_/C _11895_/C vssd1 vssd1 vccd1 vccd1 _08856_/B sky130_fd_sc_hd__nand2_1
XFILLER_112_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08786_ _08787_/B vssd1 vssd1 vccd1 vccd1 _08786_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_73_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_696 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09407_ _10236_/A _10236_/B _12770_/D _09985_/D vssd1 vssd1 vccd1 vccd1 _09410_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_164_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09338_ _09338_/A _09338_/B vssd1 vssd1 vccd1 vccd1 _09339_/C sky130_fd_sc_hd__xnor2_1
XFILLER_139_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09269_ _09269_/A _09269_/B _09275_/B vssd1 vssd1 vccd1 vccd1 _09290_/B sky130_fd_sc_hd__or3_1
X_11300_ _11299_/B _11415_/A vssd1 vssd1 vccd1 vccd1 _11711_/B sky130_fd_sc_hd__nand2b_1
XFILLER_166_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12280_ _12281_/B _12281_/A vssd1 vssd1 vccd1 vccd1 _12280_/X sky130_fd_sc_hd__and2b_1
XFILLER_5_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11231_ _11229_/A _11199_/X _11229_/B vssd1 vssd1 vccd1 vccd1 _11231_/X sky130_fd_sc_hd__o21a_1
XFILLER_150_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11162_ _11162_/A _11162_/B _11162_/C vssd1 vssd1 vccd1 vccd1 _11168_/B sky130_fd_sc_hd__and3_1
XFILLER_20_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10113_ _10113_/A _10113_/B _10119_/B vssd1 vssd1 vccd1 vccd1 _10133_/B sky130_fd_sc_hd__or3_1
XFILLER_122_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11093_ _11097_/C _17469_/D _10822_/A _10820_/Y vssd1 vssd1 vccd1 vccd1 _11099_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_15970_ _16084_/B _15970_/B vssd1 vssd1 vccd1 vccd1 _15972_/B sky130_fd_sc_hd__or2_1
XFILLER_29_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14921_ _10479_/B _10359_/B _14788_/B _10799_/B _14914_/S _14958_/A vssd1 vssd1 vccd1
+ vccd1 _14921_/X sky130_fd_sc_hd__mux4_1
X_10044_ _10419_/B _17497_/Q _12054_/B _14789_/A vssd1 vssd1 vccd1 vccd1 _10044_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_76_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14852_ _15541_/A _15463_/A _15463_/B vssd1 vssd1 vccd1 vccd1 _15624_/B sky130_fd_sc_hd__and3_1
XFILLER_91_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1042 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13803_ _13803_/A _13803_/B vssd1 vssd1 vccd1 vccd1 _13805_/B sky130_fd_sc_hd__xnor2_1
X_17571_ fanout934/X _17571_/D vssd1 vssd1 vccd1 vccd1 _17571_/Q sky130_fd_sc_hd__dfxtp_1
X_14783_ _15262_/A _15709_/A vssd1 vssd1 vccd1 vccd1 _15707_/B sky130_fd_sc_hd__or2_1
X_11995_ _09248_/B _09248_/Y _12197_/A _11994_/X vssd1 vssd1 vccd1 vccd1 _12197_/B
+ sky130_fd_sc_hd__a211oi_2
XFILLER_63_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16522_ _16522_/A _16522_/B vssd1 vssd1 vccd1 vccd1 _16524_/B sky130_fd_sc_hd__xnor2_1
X_13734_ _13735_/B _13846_/B _13735_/D _13632_/A vssd1 vssd1 vccd1 vccd1 _13736_/A
+ sky130_fd_sc_hd__a22oi_1
X_10946_ _10946_/A _10946_/B _10946_/C vssd1 vssd1 vccd1 vccd1 _10946_/X sky130_fd_sc_hd__and3_1
XFILLER_72_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_82 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16453_ _16453_/A _16453_/B vssd1 vssd1 vccd1 vccd1 _16454_/B sky130_fd_sc_hd__xnor2_1
X_13665_ _13665_/A _13778_/A vssd1 vssd1 vccd1 vccd1 _13668_/A sky130_fd_sc_hd__or2_1
X_10877_ _10878_/A _10876_/Y _11124_/C _10971_/B vssd1 vssd1 vccd1 vccd1 _11121_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_31_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15404_ _15404_/A _15404_/B vssd1 vssd1 vccd1 vccd1 _15406_/A sky130_fd_sc_hd__xnor2_1
X_12616_ _12616_/A _12616_/B vssd1 vssd1 vccd1 vccd1 _12623_/A sky130_fd_sc_hd__or2_1
X_16384_ _16385_/A _16385_/B vssd1 vssd1 vccd1 vccd1 _16384_/Y sky130_fd_sc_hd__nand2_1
XFILLER_31_368 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13596_ _13597_/A _13597_/B vssd1 vssd1 vccd1 vccd1 _13598_/A sky130_fd_sc_hd__and2_1
XFILLER_129_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15335_ _15337_/A _15337_/B vssd1 vssd1 vccd1 vccd1 _15335_/Y sky130_fd_sc_hd__nor2_1
X_12547_ _11810_/X _11818_/B _12848_/S vssd1 vssd1 vccd1 vccd1 _12547_/X sky130_fd_sc_hd__mux2_1
XFILLER_157_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15266_ _15820_/A _16262_/A _15331_/A vssd1 vssd1 vccd1 vccd1 _15337_/A sky130_fd_sc_hd__or3_2
XFILLER_8_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12478_ _12478_/A _12478_/B vssd1 vssd1 vccd1 vccd1 _12481_/C sky130_fd_sc_hd__xor2_1
XFILLER_126_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_3 _17479_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17005_ _16955_/A _16955_/B _16953_/A vssd1 vssd1 vccd1 vccd1 _17007_/B sky130_fd_sc_hd__a21oi_1
X_14217_ _14218_/A _14218_/B _14218_/C vssd1 vssd1 vccd1 vccd1 _14297_/A sky130_fd_sc_hd__o21ai_2
X_11429_ _11506_/B _11427_/C _15402_/A _11427_/A vssd1 vssd1 vccd1 vccd1 _11430_/C
+ sky130_fd_sc_hd__a22oi_1
XFILLER_6_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15197_ _16226_/B _16226_/C vssd1 vssd1 vccd1 vccd1 _15220_/A sky130_fd_sc_hd__nand2_1
XFILLER_125_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_922 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14148_ _14148_/A _14148_/B vssd1 vssd1 vccd1 vccd1 _14150_/C sky130_fd_sc_hd__xnor2_1
XFILLER_112_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14079_ _14318_/B _14301_/C _14080_/C vssd1 vssd1 vccd1 vccd1 _14081_/A sky130_fd_sc_hd__a21oi_1
XFILLER_141_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09123_ _11922_/A _09502_/B vssd1 vssd1 vccd1 vccd1 _09479_/A sky130_fd_sc_hd__nand2_1
XFILLER_163_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09054_ _09055_/A _09055_/B _09055_/C vssd1 vssd1 vccd1 vccd1 _09076_/A sky130_fd_sc_hd__a21o_1
XFILLER_117_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09956_ _09956_/A _09956_/B vssd1 vssd1 vccd1 vccd1 _09957_/B sky130_fd_sc_hd__or2_1
XFILLER_104_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08907_ _08907_/A _08907_/B vssd1 vssd1 vccd1 vccd1 _08908_/B sky130_fd_sc_hd__nor2_1
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09887_ _09765_/A _09765_/B _09765_/C vssd1 vssd1 vccd1 vccd1 _09887_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_97_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08838_ _17381_/A _11900_/D _08835_/Y _08862_/A vssd1 vssd1 vccd1 vccd1 _08839_/B
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_3415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08769_ _17403_/A _17399_/A _09030_/C _09272_/D vssd1 vssd1 vccd1 vccd1 _08773_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_45_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10800_ _11115_/A _10963_/C _10800_/C vssd1 vssd1 vccd1 vccd1 _10802_/A sky130_fd_sc_hd__and3_1
XTAP_2747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11780_ _11781_/B vssd1 vssd1 vccd1 vccd1 _11780_/Y sky130_fd_sc_hd__inv_2
XFILLER_122_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10731_ _10712_/X _10730_/Y _10631_/X _10693_/Y vssd1 vssd1 vccd1 vccd1 _10766_/C
+ sky130_fd_sc_hd__a211o_2
XFILLER_159_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_306 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13450_ _14167_/A _13450_/B _13450_/C _14050_/D vssd1 vssd1 vccd1 vccd1 _13569_/A
+ sky130_fd_sc_hd__and4_1
X_10662_ _10662_/A _10662_/B _10662_/C vssd1 vssd1 vccd1 vccd1 _10662_/X sky130_fd_sc_hd__and3_1
XFILLER_13_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12401_ _12710_/A _12401_/B vssd1 vssd1 vccd1 vccd1 _12401_/X sky130_fd_sc_hd__or2_1
X_13381_ _13221_/A _13224_/A _13504_/A _13380_/X vssd1 vssd1 vccd1 vccd1 _13504_/B
+ sky130_fd_sc_hd__a211oi_1
X_10593_ _10593_/A _10593_/B vssd1 vssd1 vccd1 vccd1 _10595_/A sky130_fd_sc_hd__nand2_1
XFILLER_154_502 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15120_ _15119_/A _15119_/B _17156_/B vssd1 vssd1 vccd1 vccd1 _15120_/X sky130_fd_sc_hd__a21o_1
XFILLER_5_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12332_ _17407_/A _12166_/B _12167_/A _12165_/B vssd1 vssd1 vccd1 vccd1 _12333_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_139_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15051_ _15051_/A _15456_/B _15050_/X vssd1 vssd1 vccd1 vccd1 _15051_/X sky130_fd_sc_hd__or3b_1
X_12263_ _12263_/A _12263_/B vssd1 vssd1 vccd1 vccd1 _12265_/C sky130_fd_sc_hd__xnor2_1
XFILLER_147_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14002_ _14176_/A _14366_/B _14002_/C vssd1 vssd1 vccd1 vccd1 _14092_/B sky130_fd_sc_hd__nand3_1
XFILLER_135_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11214_ _11216_/A _11216_/B vssd1 vssd1 vccd1 vccd1 _11214_/Y sky130_fd_sc_hd__nand2_1
XFILLER_135_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12194_ _12360_/A _12193_/B _12193_/C vssd1 vssd1 vccd1 vccd1 _12194_/X sky130_fd_sc_hd__a21o_1
Xoutput73 _17477_/Q vssd1 vssd1 vccd1 vccd1 leds[11] sky130_fd_sc_hd__clkbuf_1
X_11145_ _11145_/A _11145_/B _11145_/C vssd1 vssd1 vccd1 vccd1 _11153_/B sky130_fd_sc_hd__and3_1
XFILLER_150_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput84 _17434_/Q vssd1 vssd1 vccd1 vccd1 o_wb_data[0] sky130_fd_sc_hd__clkbuf_1
XFILLER_49_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput95 _17435_/Q vssd1 vssd1 vccd1 vccd1 o_wb_data[1] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11076_ _11059_/A _11059_/B _11059_/C vssd1 vssd1 vccd1 vccd1 _11077_/C sky130_fd_sc_hd__a21oi_1
X_15953_ _15953_/A _15953_/B vssd1 vssd1 vccd1 vccd1 _15954_/B sky130_fd_sc_hd__nand2_1
XFILLER_76_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14904_ _08731_/A _15147_/A vssd1 vssd1 vccd1 vccd1 _14905_/D sky130_fd_sc_hd__nand2b_1
X_10027_ _10028_/A _10027_/B _10027_/C _10027_/D vssd1 vssd1 vccd1 vccd1 _10028_/B
+ sky130_fd_sc_hd__and4b_1
X_15884_ _15884_/A _15884_/B vssd1 vssd1 vccd1 vccd1 _15884_/Y sky130_fd_sc_hd__nand2_1
XFILLER_36_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14835_ _17063_/A _14836_/B _14933_/B vssd1 vssd1 vccd1 vccd1 _15108_/A sky130_fd_sc_hd__and3_2
XFILLER_17_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17554_ fanout940/X _17554_/D vssd1 vssd1 vccd1 vccd1 _17554_/Q sky130_fd_sc_hd__dfxtp_1
X_11978_ _11978_/A _11978_/B vssd1 vssd1 vccd1 vccd1 _11980_/A sky130_fd_sc_hd__nor2_1
X_14766_ _14766_/A _17028_/A vssd1 vssd1 vccd1 vccd1 _17023_/B sky130_fd_sc_hd__or2_1
XFILLER_16_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16505_ _16505_/A _16505_/B vssd1 vssd1 vccd1 vccd1 _16505_/X sky130_fd_sc_hd__or2_1
XFILLER_108_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10929_ _11057_/A _11057_/B _11057_/C vssd1 vssd1 vccd1 vccd1 _11059_/A sky130_fd_sc_hd__a21o_1
X_13717_ _13818_/B _13717_/B vssd1 vssd1 vccd1 vccd1 _13720_/A sky130_fd_sc_hd__and2_1
XFILLER_16_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17485_ fanout950/X _17485_/D vssd1 vssd1 vccd1 vccd1 _17485_/Q sky130_fd_sc_hd__dfxtp_1
X_14697_ _14698_/B _14699_/A vssd1 vssd1 vccd1 vccd1 _14729_/A sky130_fd_sc_hd__nor2_1
X_16436_ _16436_/A _16436_/B vssd1 vssd1 vccd1 vccd1 _16437_/B sky130_fd_sc_hd__xnor2_1
XFILLER_158_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13648_ _13749_/B _13648_/B _13648_/C vssd1 vssd1 vccd1 vccd1 _13648_/X sky130_fd_sc_hd__and3_1
XFILLER_32_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_852 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16367_ _16367_/A _16367_/B vssd1 vssd1 vccd1 vccd1 _16369_/A sky130_fd_sc_hd__xor2_2
X_13579_ _13579_/A _13579_/B vssd1 vssd1 vccd1 vccd1 _13597_/A sky130_fd_sc_hd__xnor2_1
XFILLER_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15318_ _15628_/A _16219_/A1 _12710_/B _15315_/X _15317_/X vssd1 vssd1 vccd1 vccd1
+ _15321_/C sky130_fd_sc_hd__o311a_1
XFILLER_145_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16298_ _16298_/A _16571_/B _14777_/A vssd1 vssd1 vccd1 vccd1 _16299_/B sky130_fd_sc_hd__or3b_1
XFILLER_117_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15249_ _15244_/B _14929_/X _15713_/B1 _14906_/B vssd1 vssd1 vccd1 vccd1 _15249_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_114_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_398 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout307 _14733_/S vssd1 vssd1 vccd1 vccd1 _17371_/A sky130_fd_sc_hd__clkbuf_4
X_09810_ _09789_/A _09933_/A _09789_/B _09920_/A vssd1 vssd1 vccd1 vccd1 _09811_/B
+ sky130_fd_sc_hd__o31ai_2
Xfanout318 _14213_/A vssd1 vssd1 vccd1 vccd1 _13966_/A sky130_fd_sc_hd__buf_2
Xfanout329 _08988_/B vssd1 vssd1 vccd1 vccd1 _13434_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_86_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09741_ _09768_/B _09832_/A _09768_/A vssd1 vssd1 vccd1 vccd1 _09812_/B sky130_fd_sc_hd__o21a_1
XFILLER_86_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_850 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09672_ _09674_/B _09819_/A _09674_/A vssd1 vssd1 vccd1 vccd1 _09678_/B sky130_fd_sc_hd__o21a_1
XFILLER_39_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_224 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1013 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09106_ _09106_/A _09106_/B vssd1 vssd1 vccd1 vccd1 _09108_/A sky130_fd_sc_hd__nor2_1
XFILLER_148_395 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09037_ _09037_/A _09037_/B vssd1 vssd1 vccd1 vccd1 _09039_/B sky130_fd_sc_hd__xnor2_1
XFILLER_151_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_730 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout830 _14851_/A vssd1 vssd1 vccd1 vccd1 _14895_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_77_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout841 _11387_/B vssd1 vssd1 vccd1 vccd1 _10962_/B sky130_fd_sc_hd__clkbuf_4
Xfanout852 _17484_/Q vssd1 vssd1 vccd1 vccd1 _14849_/A sky130_fd_sc_hd__buf_4
XFILLER_104_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09939_ _09939_/A _09939_/B vssd1 vssd1 vccd1 vccd1 _09951_/A sky130_fd_sc_hd__nor2_1
XFILLER_133_20 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout863 _17483_/Q vssd1 vssd1 vccd1 vccd1 _12295_/D sky130_fd_sc_hd__clkbuf_4
Xfanout874 _17482_/Q vssd1 vssd1 vccd1 vccd1 fanout874/X sky130_fd_sc_hd__clkbuf_4
XFILLER_86_850 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout885 _17481_/Q vssd1 vssd1 vccd1 vccd1 _11427_/C sky130_fd_sc_hd__buf_2
X_12950_ _13903_/A _13866_/C _12950_/C vssd1 vssd1 vccd1 vccd1 _13092_/B sky130_fd_sc_hd__nand3_1
Xfanout896 _17479_/Q vssd1 vssd1 vccd1 vccd1 _15003_/B sky130_fd_sc_hd__buf_4
XTAP_3201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11901_ _11901_/A _11901_/B vssd1 vssd1 vccd1 vccd1 _11903_/A sky130_fd_sc_hd__nor2_1
XFILLER_85_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12881_ _12881_/A _12881_/B vssd1 vssd1 vccd1 vccd1 _12882_/B sky130_fd_sc_hd__nand2_1
XFILLER_85_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11832_ _11829_/Y _11831_/Y _17365_/A vssd1 vssd1 vccd1 vccd1 _11832_/X sky130_fd_sc_hd__mux2_1
X_14620_ _14621_/A _14621_/B _14621_/C vssd1 vssd1 vccd1 vccd1 _14661_/A sky130_fd_sc_hd__a21oi_1
XTAP_3289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_611 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14551_ _14765_/A _14641_/C _14679_/B vssd1 vssd1 vccd1 vccd1 _14553_/A sky130_fd_sc_hd__a21boi_1
XTAP_2588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11763_ _11750_/A _16794_/A _11750_/B vssd1 vssd1 vccd1 vccd1 _11763_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10714_ _10715_/A _10715_/B _10715_/C vssd1 vssd1 vccd1 vccd1 _10714_/X sky130_fd_sc_hd__a21o_1
XFILLER_42_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13502_ _13347_/B _13349_/B _13347_/A vssd1 vssd1 vccd1 vccd1 _13503_/B sky130_fd_sc_hd__o21ba_1
XTAP_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17270_ _17599_/Q _17282_/A2 _17282_/B1 vssd1 vssd1 vccd1 vccd1 _17270_/X sky130_fd_sc_hd__a21o_1
X_14482_ _13840_/S _12866_/B _14210_/B _14482_/B1 vssd1 vssd1 vccd1 vccd1 _14482_/X
+ sky130_fd_sc_hd__o31a_1
XTAP_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11694_ _11672_/A _11672_/B _11672_/C vssd1 vssd1 vccd1 vccd1 _11694_/X sky130_fd_sc_hd__a21o_1
XFILLER_14_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13433_ _14050_/B _13551_/D _13434_/D _14213_/A vssd1 vssd1 vccd1 vccd1 _13435_/A
+ sky130_fd_sc_hd__a22oi_1
X_16221_ _16221_/A _16221_/B _16215_/X vssd1 vssd1 vccd1 vccd1 _16221_/X sky130_fd_sc_hd__or3b_1
X_10645_ _11122_/A _10851_/B _10745_/D _10786_/B vssd1 vssd1 vccd1 vccd1 _10648_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_127_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16152_ _16152_/A _16812_/A vssd1 vssd1 vccd1 vccd1 _16153_/B sky130_fd_sc_hd__nand2_1
XFILLER_6_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13364_ _13482_/A _13364_/B vssd1 vssd1 vccd1 vccd1 _13366_/B sky130_fd_sc_hd__nor2_1
X_10576_ _10573_/X _10575_/Y _10463_/B _10471_/X vssd1 vssd1 vccd1 vccd1 _10579_/A
+ sky130_fd_sc_hd__a211oi_2
X_12315_ _12316_/A _12316_/B _12316_/C vssd1 vssd1 vccd1 vccd1 _12526_/A sky130_fd_sc_hd__a21o_1
X_15103_ _15100_/Y _15102_/Y _15103_/S vssd1 vssd1 vccd1 vccd1 _15103_/X sky130_fd_sc_hd__mux2_1
X_16083_ _16084_/A _16084_/B _16082_/X vssd1 vssd1 vccd1 vccd1 _16197_/A sky130_fd_sc_hd__o21ba_1
XFILLER_154_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13295_ _13295_/A _13295_/B _13295_/C vssd1 vssd1 vccd1 vccd1 _13308_/B sky130_fd_sc_hd__nand3_1
XFILLER_170_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15034_ _15131_/A _15034_/B vssd1 vssd1 vccd1 vccd1 _15034_/Y sky130_fd_sc_hd__nand2_1
X_12246_ _12247_/A _12247_/B vssd1 vssd1 vccd1 vccd1 _12429_/B sky130_fd_sc_hd__nor2_1
XFILLER_107_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_549 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12177_ _12177_/A _12177_/B vssd1 vssd1 vccd1 vccd1 _12179_/C sky130_fd_sc_hd__xnor2_1
XFILLER_123_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11128_ _11130_/B _11130_/C _11130_/A vssd1 vssd1 vccd1 vccd1 _11128_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16985_ _16986_/A _16986_/B vssd1 vssd1 vccd1 vccd1 _17046_/A sky130_fd_sc_hd__and2b_1
X_11059_ _11059_/A _11059_/B _11059_/C vssd1 vssd1 vccd1 vccd1 _11077_/A sky130_fd_sc_hd__and3_1
X_15936_ _15937_/A _15937_/B vssd1 vssd1 vccd1 vccd1 _16072_/A sky130_fd_sc_hd__and2_1
XFILLER_36_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15867_ _15867_/A _15867_/B vssd1 vssd1 vccd1 vccd1 _15875_/A sky130_fd_sc_hd__and2_1
XFILLER_25_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_950 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17606_ fanout936/X _17606_/D vssd1 vssd1 vccd1 vccd1 _17606_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14818_ _16576_/B _16577_/A _12869_/C vssd1 vssd1 vccd1 vccd1 _16649_/C sky130_fd_sc_hd__a21o_1
XFILLER_24_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15798_ _15705_/B _15705_/C _15705_/A vssd1 vssd1 vccd1 vccd1 _15798_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_17_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17537_ fanout947/X _17537_/D vssd1 vssd1 vccd1 vccd1 _17537_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_33_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14749_ _14750_/A _14750_/B vssd1 vssd1 vccd1 vccd1 _14751_/A sky130_fd_sc_hd__or2_1
XFILLER_32_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17468_ fanout955/X _17468_/D vssd1 vssd1 vccd1 vccd1 _17468_/Q sky130_fd_sc_hd__dfxtp_1
X_16419_ _16419_/A _16419_/B vssd1 vssd1 vccd1 vccd1 _16420_/A sky130_fd_sc_hd__xnor2_1
X_17399_ _17399_/A _17421_/B vssd1 vssd1 vccd1 vccd1 _17399_/X sky130_fd_sc_hd__or2_1
XFILLER_146_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_251 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout126 _17199_/B vssd1 vssd1 vccd1 vccd1 _17244_/B sky130_fd_sc_hd__buf_2
XFILLER_87_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout137 _15199_/Y vssd1 vssd1 vccd1 vccd1 _16355_/A sky130_fd_sc_hd__clkbuf_2
Xfanout148 _14969_/Y vssd1 vssd1 vccd1 vccd1 _15918_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_59_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout159 _17371_/B vssd1 vssd1 vccd1 vccd1 _17377_/B sky130_fd_sc_hd__buf_2
XFILLER_101_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09724_ _09725_/A _09725_/B _09725_/C vssd1 vssd1 vccd1 vccd1 _09724_/X sky130_fd_sc_hd__a21o_2
XFILLER_101_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_820 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09655_ _09655_/A _09784_/A vssd1 vssd1 vccd1 vccd1 _09656_/C sky130_fd_sc_hd__nor2_1
XFILLER_28_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09586_ _09587_/A _09585_/Y _09730_/C _10421_/D vssd1 vssd1 vccd1 vccd1 _09727_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_83_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_647 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10430_ _10430_/A _10657_/B vssd1 vssd1 vccd1 vccd1 _14956_/A sky130_fd_sc_hd__and2_2
XFILLER_164_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10361_ _11027_/A _10479_/B _10594_/B _10591_/A vssd1 vssd1 vccd1 vccd1 _10362_/B
+ sky130_fd_sc_hd__a22oi_1
XFILLER_136_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_387 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12100_ _12097_/X _12268_/B _11891_/A _11891_/Y vssd1 vssd1 vccd1 vccd1 _12122_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_152_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13080_ _13080_/A _13450_/B _13080_/C _13080_/D vssd1 vssd1 vccd1 vccd1 _13213_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_128_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10292_ _10293_/A _10291_/Y _14788_/A _10647_/D vssd1 vssd1 vccd1 vccd1 _10399_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_152_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12031_ _14911_/B _12031_/B vssd1 vssd1 vccd1 vccd1 _12031_/Y sky130_fd_sc_hd__nand2_1
XFILLER_104_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout660 _16974_/A vssd1 vssd1 vccd1 vccd1 _14301_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_144_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout671 _12275_/D vssd1 vssd1 vccd1 vccd1 _11902_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_120_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_872 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16770_ _16770_/A _16770_/B _16770_/C vssd1 vssd1 vccd1 vccd1 _16771_/B sky130_fd_sc_hd__or3_1
Xfanout682 fanout690/X vssd1 vssd1 vccd1 vccd1 _14063_/C sky130_fd_sc_hd__buf_4
X_13982_ _13982_/A _13982_/B vssd1 vssd1 vccd1 vccd1 _13985_/A sky130_fd_sc_hd__xnor2_1
Xfanout693 fanout699/X vssd1 vssd1 vccd1 vccd1 _16722_/A sky130_fd_sc_hd__buf_4
XFILLER_101_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15721_ _17131_/A _15700_/Y _15720_/X vssd1 vssd1 vccd1 vccd1 _15721_/X sky130_fd_sc_hd__a21o_1
XTAP_3031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12933_ _12933_/A _12933_/B _12933_/C vssd1 vssd1 vccd1 vccd1 _12935_/A sky130_fd_sc_hd__nor3_1
XTAP_3042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15652_ _15742_/A _15742_/B vssd1 vssd1 vccd1 vccd1 _15743_/A sky130_fd_sc_hd__nor2_1
XFILLER_18_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12864_ _12864_/A vssd1 vssd1 vccd1 vccd1 _12864_/Y sky130_fd_sc_hd__inv_2
XTAP_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14603_ _14603_/A _14646_/A vssd1 vssd1 vccd1 vccd1 _14606_/A sky130_fd_sc_hd__and2_1
XTAP_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11815_ _12025_/A _11815_/B vssd1 vssd1 vccd1 vccd1 _14978_/B sky130_fd_sc_hd__and2_1
XTAP_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12795_ _12795_/A _13080_/C vssd1 vssd1 vccd1 vccd1 _12796_/B sky130_fd_sc_hd__nand2_1
XTAP_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15583_ _15584_/A _15584_/B vssd1 vssd1 vccd1 vccd1 _15583_/Y sky130_fd_sc_hd__nand2_1
XTAP_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_424 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17322_ _11961_/B _17322_/A2 _17321_/X _17388_/C1 vssd1 vssd1 vccd1 vccd1 _17490_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11746_ _11758_/A _11747_/B vssd1 vssd1 vccd1 vccd1 _16794_/A sky130_fd_sc_hd__nand2_1
X_14534_ _14534_/A _14534_/B vssd1 vssd1 vccd1 vccd1 _14534_/Y sky130_fd_sc_hd__nand2_1
XTAP_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17253_ _17561_/Q _17292_/B vssd1 vssd1 vccd1 vccd1 _17253_/X sky130_fd_sc_hd__and2_1
XFILLER_128_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11677_ _15715_/A _15008_/B _11681_/A _11658_/D vssd1 vssd1 vccd1 vccd1 _11678_/B
+ sky130_fd_sc_hd__a22o_1
X_14465_ _14465_/A _14465_/B vssd1 vssd1 vccd1 vccd1 _14524_/A sky130_fd_sc_hd__nand2_1
XFILLER_169_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16204_ _16098_/A _16101_/Y _16203_/B _15523_/A vssd1 vssd1 vccd1 vccd1 _16205_/B
+ sky130_fd_sc_hd__a31o_1
X_10628_ _10623_/X _10627_/X _10614_/X _10615_/Y vssd1 vssd1 vccd1 vccd1 _10632_/B
+ sky130_fd_sc_hd__o211ai_4
X_13416_ _13417_/A _13417_/B _13417_/C vssd1 vssd1 vccd1 vccd1 _13418_/A sky130_fd_sc_hd__o21ai_1
XFILLER_174_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17184_ input25/X _17428_/C vssd1 vssd1 vccd1 vccd1 _17362_/B sky130_fd_sc_hd__nand2_2
X_14396_ _14396_/A _14396_/B vssd1 vssd1 vccd1 vccd1 _14396_/X sky130_fd_sc_hd__and2_1
XFILLER_139_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16135_ _16315_/C _16662_/D _16234_/C vssd1 vssd1 vccd1 vccd1 _16137_/A sky130_fd_sc_hd__o21a_1
X_13347_ _13347_/A _13347_/B vssd1 vssd1 vccd1 vccd1 _13349_/A sky130_fd_sc_hd__nor2_1
XFILLER_115_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10559_ _10559_/A _11027_/D vssd1 vssd1 vccd1 vccd1 _10669_/A sky130_fd_sc_hd__nand2_1
XFILLER_155_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16066_ _16066_/A _16066_/B vssd1 vssd1 vccd1 vccd1 _16068_/A sky130_fd_sc_hd__xnor2_1
X_13278_ _13735_/B _13522_/D _14063_/C _13632_/A vssd1 vssd1 vccd1 vccd1 _13280_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_142_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12229_ _13831_/S _17164_/B _12229_/C vssd1 vssd1 vccd1 vccd1 _12230_/B sky130_fd_sc_hd__or3_2
X_15017_ _14977_/X _15014_/Y _15016_/Y _16977_/A _11675_/B vssd1 vssd1 vccd1 vccd1
+ _17544_/D sky130_fd_sc_hd__o32a_1
XFILLER_170_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16968_ _16863_/A _16863_/B _16916_/A _16967_/X vssd1 vssd1 vccd1 vccd1 _16969_/B
+ sky130_fd_sc_hd__a31oi_2
XFILLER_111_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15919_ _16025_/A _16662_/C _15917_/Y _15916_/X vssd1 vssd1 vccd1 vccd1 _15921_/A
+ sky130_fd_sc_hd__o31a_1
XFILLER_49_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16899_ _16829_/A _16828_/A _16828_/B _16830_/B _16830_/A vssd1 vssd1 vccd1 vccd1
+ _16900_/C sky130_fd_sc_hd__a32o_1
X_09440_ _09441_/A _09441_/B _09441_/C vssd1 vssd1 vccd1 vccd1 _09440_/X sky130_fd_sc_hd__a21o_2
XFILLER_64_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09371_ _10559_/A _09555_/C vssd1 vssd1 vccd1 vccd1 _09386_/A sky130_fd_sc_hd__nand2_1
XFILLER_33_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_722 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_842 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09707_ _16989_/A _09707_/B vssd1 vssd1 vccd1 vccd1 _09709_/B sky130_fd_sc_hd__xnor2_4
XFILLER_28_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwb_buttons_leds_967 vssd1 vssd1 vccd1 vccd1 wb_buttons_leds_967/HI led_enb[9] sky130_fd_sc_hd__conb_1
XFILLER_28_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09638_ _14770_/A _10067_/B _10446_/B _09797_/A vssd1 vssd1 vccd1 vccd1 _09638_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_169_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09569_ _16933_/A _16982_/B vssd1 vssd1 vccd1 vccd1 _09570_/B sky130_fd_sc_hd__nand2_1
XFILLER_31_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11600_ _11558_/B _11600_/B vssd1 vssd1 vccd1 vccd1 _11639_/B sky130_fd_sc_hd__and2b_1
XFILLER_12_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12580_ _12581_/A _12581_/B vssd1 vssd1 vccd1 vccd1 _12761_/A sky130_fd_sc_hd__and2b_1
XFILLER_142_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11531_ _11496_/B _11493_/B _11493_/C vssd1 vssd1 vccd1 vccd1 _11532_/B sky130_fd_sc_hd__a21oi_1
XFILLER_168_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14250_ _14330_/B _14250_/B vssd1 vssd1 vccd1 vccd1 _14252_/C sky130_fd_sc_hd__nand2_1
X_11462_ _11703_/A _11703_/B vssd1 vssd1 vccd1 vccd1 _11465_/A sky130_fd_sc_hd__or2_1
XFILLER_7_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13201_ _13332_/A _13202_/B _13202_/C vssd1 vssd1 vccd1 vccd1 _13201_/Y sky130_fd_sc_hd__a21oi_1
X_10413_ _14787_/A _10786_/B _10743_/D _14786_/A vssd1 vssd1 vccd1 vccd1 _10413_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_99_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_354 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14181_ _14254_/A _14181_/B _14181_/C vssd1 vssd1 vccd1 vccd1 _14273_/B sky130_fd_sc_hd__nand3_1
XFILLER_99_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11393_ _11393_/A _11393_/B _11393_/C vssd1 vssd1 vccd1 vccd1 _11394_/B sky130_fd_sc_hd__or3_1
XFILLER_137_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13132_ _13264_/A _13130_/Y _12956_/A _12960_/A vssd1 vssd1 vccd1 vccd1 _13132_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_109_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10344_ _10070_/A _10072_/Y _10345_/A _10343_/Y vssd1 vssd1 vccd1 vccd1 _10581_/A
+ sky130_fd_sc_hd__a211oi_1
XFILLER_151_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13063_ _13063_/A _13063_/B vssd1 vssd1 vccd1 vccd1 _13065_/C sky130_fd_sc_hd__nand2_1
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10275_ _10276_/A _10276_/B vssd1 vssd1 vccd1 vccd1 _10275_/X sky130_fd_sc_hd__and2_1
XFILLER_133_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12014_ _12375_/A _12014_/B vssd1 vssd1 vccd1 vccd1 _12374_/A sky130_fd_sc_hd__nor2_1
XFILLER_2_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16822_ _16822_/A _16822_/B vssd1 vssd1 vccd1 vccd1 _16823_/B sky130_fd_sc_hd__and2_1
XFILLER_66_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout490 _09299_/B vssd1 vssd1 vccd1 vccd1 _12275_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_47_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16753_ _16753_/A _16835_/A vssd1 vssd1 vccd1 vccd1 _16767_/A sky130_fd_sc_hd__or2_1
X_13965_ _14213_/B _13966_/C _13966_/D _13966_/A vssd1 vssd1 vccd1 vccd1 _13967_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15704_ _15620_/A _15618_/B _15620_/B _15616_/Y vssd1 vssd1 vccd1 vccd1 _15705_/C
+ sky130_fd_sc_hd__a31o_1
X_12916_ _13072_/B _12916_/B vssd1 vssd1 vccd1 vccd1 _12918_/C sky130_fd_sc_hd__nor2_1
XFILLER_46_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16684_ _16684_/A _16684_/B vssd1 vssd1 vccd1 vccd1 _16684_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_73_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13896_ _13896_/A _13896_/B vssd1 vssd1 vccd1 vccd1 _13898_/A sky130_fd_sc_hd__nor2_1
XFILLER_61_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_396 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15635_ _15624_/A _16401_/C1 _15615_/X _15634_/Y vssd1 vssd1 vccd1 vccd1 _15636_/A
+ sky130_fd_sc_hd__a22o_1
X_12847_ _14421_/S _12847_/B vssd1 vssd1 vccd1 vccd1 _12847_/X sky130_fd_sc_hd__and2_1
XTAP_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15566_ _15932_/A _16619_/A vssd1 vssd1 vccd1 vccd1 _15666_/A sky130_fd_sc_hd__nor2_1
XFILLER_14_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12778_ _12778_/A _12778_/B _12778_/C vssd1 vssd1 vccd1 vccd1 _12779_/B sky130_fd_sc_hd__and3_1
XTAP_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17305_ input62/X _17321_/B _17321_/C vssd1 vssd1 vccd1 vccd1 _17305_/X sky130_fd_sc_hd__or3_1
XFILLER_9_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14517_ _14519_/B vssd1 vssd1 vccd1 vccd1 _14517_/Y sky130_fd_sc_hd__inv_2
XFILLER_147_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11729_ _11731_/B _11729_/B _11729_/C vssd1 vssd1 vccd1 vccd1 _11736_/A sky130_fd_sc_hd__nor3_1
XFILLER_159_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15497_ _15750_/A _16812_/A vssd1 vssd1 vccd1 vccd1 _15498_/B sky130_fd_sc_hd__nand2_1
XFILLER_9_98 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_786 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17236_ _17446_/Q _17275_/A2 _17234_/X _17235_/X _17364_/C1 vssd1 vssd1 vccd1 vccd1
+ _17446_/D sky130_fd_sc_hd__o221a_1
X_14448_ _14383_/A _14450_/B _14383_/B _16913_/C vssd1 vssd1 vccd1 vccd1 _14451_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_174_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17167_ _17167_/A _17167_/B _17167_/C vssd1 vssd1 vccd1 vccd1 _17167_/X sky130_fd_sc_hd__and3_1
X_14379_ _14446_/A _14379_/B vssd1 vssd1 vccd1 vccd1 _14381_/B sky130_fd_sc_hd__nor2_1
XFILLER_142_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16118_ _15175_/A _16116_/X _16117_/X _15808_/A vssd1 vssd1 vccd1 vccd1 _16122_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_171_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17098_ _17100_/C _17134_/C _14867_/A vssd1 vssd1 vccd1 vccd1 _17099_/A sky130_fd_sc_hd__a21boi_1
XFILLER_116_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16049_ _15927_/B _15941_/B _15925_/Y vssd1 vssd1 vccd1 vccd1 _16051_/B sky130_fd_sc_hd__a21oi_1
X_08940_ _17373_/A _09325_/B _09350_/B _11895_/C vssd1 vssd1 vccd1 vccd1 _08941_/B
+ sky130_fd_sc_hd__and4_1
X_08871_ _08868_/X _08869_/Y _08844_/X _08908_/A vssd1 vssd1 vccd1 vccd1 _08873_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_9_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09423_ _09423_/A _09423_/B vssd1 vssd1 vccd1 vccd1 _09433_/A sky130_fd_sc_hd__xnor2_1
XFILLER_25_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_506 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09354_ _09354_/A _09354_/B _09355_/B vssd1 vssd1 vccd1 vccd1 _09366_/A sky130_fd_sc_hd__or3_1
XFILLER_21_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09285_ _08791_/B _12334_/B _12328_/B _08791_/A vssd1 vssd1 vccd1 vccd1 _09285_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_165_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_438 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_611 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_666 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10060_ _10086_/A vssd1 vssd1 vccd1 vccd1 _10060_/Y sky130_fd_sc_hd__inv_2
XFILLER_102_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_552 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10962_ _11097_/C _10962_/B vssd1 vssd1 vccd1 vccd1 _10966_/A sky130_fd_sc_hd__nand2_1
XFILLER_29_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13750_ _13749_/A _13749_/B _13751_/A vssd1 vssd1 vccd1 vccd1 _13861_/A sky130_fd_sc_hd__a21o_1
XFILLER_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_845 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12701_ _13628_/B vssd1 vssd1 vccd1 vccd1 _12701_/Y sky130_fd_sc_hd__clkinv_2
X_10893_ _10893_/A _10893_/B _10893_/C vssd1 vssd1 vccd1 vccd1 _11112_/A sky130_fd_sc_hd__and3_1
X_13681_ _13681_/A _13681_/B vssd1 vssd1 vccd1 vccd1 _13683_/A sky130_fd_sc_hd__nor2_1
XFILLER_44_878 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15420_ _15336_/Y _15346_/B _15335_/Y vssd1 vssd1 vccd1 vccd1 _15422_/B sky130_fd_sc_hd__a21o_1
X_12632_ _12481_/A _12481_/Y _12630_/X _12631_/Y vssd1 vssd1 vccd1 vccd1 _12676_/A
+ sky130_fd_sc_hd__a211oi_2
XFILLER_54_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1022 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12563_ _12563_/A _12730_/A vssd1 vssd1 vccd1 vccd1 _12570_/A sky130_fd_sc_hd__and2_1
XFILLER_34_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15351_ _15352_/A _15352_/B vssd1 vssd1 vccd1 vccd1 _15351_/X sky130_fd_sc_hd__or2_1
X_11514_ _11514_/A _11558_/A _11514_/C vssd1 vssd1 vccd1 vccd1 _11526_/A sky130_fd_sc_hd__or3_1
X_14302_ _14302_/A _14302_/B vssd1 vssd1 vccd1 vccd1 _14304_/A sky130_fd_sc_hd__nor2_1
XFILLER_129_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12494_ _12494_/A _12494_/B vssd1 vssd1 vccd1 vccd1 _12496_/A sky130_fd_sc_hd__nor2_1
X_15282_ _15283_/A _15283_/B vssd1 vssd1 vccd1 vccd1 _15355_/A sky130_fd_sc_hd__nor2_1
XFILLER_8_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17021_ _17018_/A _17066_/A _17066_/B vssd1 vssd1 vccd1 vccd1 _17021_/Y sky130_fd_sc_hd__a21oi_1
X_11445_ _11444_/A _11444_/Y _11396_/X _11421_/Y vssd1 vssd1 vccd1 vccd1 _11453_/B
+ sky130_fd_sc_hd__a211o_1
X_14233_ _14159_/B _14161_/B _14159_/A vssd1 vssd1 vccd1 vccd1 _14235_/B sky130_fd_sc_hd__o21ba_1
XFILLER_137_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14164_ _14165_/A _14165_/B vssd1 vssd1 vccd1 vccd1 _14164_/X sky130_fd_sc_hd__and2b_1
X_11376_ _11376_/A _11376_/B _11376_/C vssd1 vssd1 vccd1 vccd1 _11395_/B sky130_fd_sc_hd__nand3_2
XFILLER_153_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13115_ _13248_/B _13115_/B vssd1 vssd1 vccd1 vccd1 _13117_/C sky130_fd_sc_hd__or2_1
X_10327_ _10560_/B _10594_/B _10326_/C vssd1 vssd1 vccd1 vccd1 _10329_/C sky130_fd_sc_hd__a21o_1
XFILLER_152_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14095_ _14254_/A _14094_/B _14094_/C vssd1 vssd1 vccd1 vccd1 _14096_/B sky130_fd_sc_hd__a21oi_1
XFILLER_113_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13046_ _13046_/A _13046_/B _13046_/C vssd1 vssd1 vccd1 vccd1 _13047_/B sky130_fd_sc_hd__nand3_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10258_ _10372_/A _10257_/B _10257_/A vssd1 vssd1 vccd1 vccd1 _10260_/B sky130_fd_sc_hd__o21ba_1
XFILLER_59_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_915 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10189_ _10207_/A _10161_/X _10188_/A _10188_/Y vssd1 vssd1 vccd1 vccd1 _10192_/B
+ sky130_fd_sc_hd__o211a_1
X_16805_ _08743_/A _16787_/Y _16793_/X _16804_/X vssd1 vssd1 vccd1 vccd1 _16805_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_82_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14997_ _10146_/B _10016_/D _10036_/D _10993_/D _09925_/A _10182_/C vssd1 vssd1 vccd1
+ vccd1 _14999_/B sky130_fd_sc_hd__mux4_1
XFILLER_81_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16736_ _14925_/Y _15313_/Y _16734_/X _16735_/Y vssd1 vssd1 vccd1 vccd1 _16736_/X
+ sky130_fd_sc_hd__a211o_1
X_13948_ _13948_/A _13948_/B _13948_/C _14094_/B vssd1 vssd1 vccd1 vccd1 _13949_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_46_171 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16667_ _16667_/A _16814_/A _16813_/B _16938_/D vssd1 vssd1 vccd1 vccd1 _16670_/C
+ sky130_fd_sc_hd__or4_1
XFILLER_34_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13879_ _14155_/A _14213_/C vssd1 vssd1 vccd1 vccd1 _13880_/B sky130_fd_sc_hd__nand2_1
XFILLER_61_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_664 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15618_ _15616_/Y _15618_/B vssd1 vssd1 vccd1 vccd1 _15621_/A sky130_fd_sc_hd__nand2b_1
X_16598_ _16507_/A _16507_/B _16505_/X vssd1 vssd1 vccd1 vccd1 _16600_/B sky130_fd_sc_hd__a21boi_1
XFILLER_61_185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15549_ _16315_/B _15755_/B vssd1 vssd1 vccd1 vccd1 _15655_/A sky130_fd_sc_hd__nor2_1
X_09070_ _09051_/A _09051_/B _09051_/C vssd1 vssd1 vccd1 vccd1 _09071_/C sky130_fd_sc_hd__a21oi_1
XFILLER_129_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17219_ _17582_/Q _17225_/A2 _17225_/B1 vssd1 vssd1 vccd1 vccd1 _17219_/X sky130_fd_sc_hd__a21o_1
XFILLER_162_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09972_ _09960_/A _09960_/C _09960_/B vssd1 vssd1 vccd1 vccd1 _09972_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_170_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_18 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08923_ _08923_/A _08923_/B vssd1 vssd1 vccd1 vccd1 _09052_/B sky130_fd_sc_hd__xnor2_1
XFILLER_131_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_904 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08854_ _08854_/A _08854_/B vssd1 vssd1 vccd1 vccd1 _08856_/A sky130_fd_sc_hd__nor2_1
XFILLER_85_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_222 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08785_ _08791_/B _09058_/C _09446_/D _17391_/A vssd1 vssd1 vccd1 vccd1 _08787_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_85_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09406_ _09411_/A _09411_/B vssd1 vssd1 vccd1 vccd1 _09417_/A sky130_fd_sc_hd__nor2_1
XFILLER_125_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09337_ _09334_/A _09335_/Y _09344_/A _09316_/X vssd1 vssd1 vccd1 vccd1 _09344_/B
+ sky130_fd_sc_hd__a211oi_2
XFILLER_21_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09268_ _09268_/A _09411_/A vssd1 vssd1 vccd1 vccd1 _09275_/B sky130_fd_sc_hd__nor2_1
XFILLER_154_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09199_ _17407_/A _09555_/C _09198_/C vssd1 vssd1 vccd1 vccd1 _09200_/B sky130_fd_sc_hd__a21o_1
XFILLER_147_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11230_ _11229_/Y _16387_/A vssd1 vssd1 vccd1 vccd1 _11717_/A sky130_fd_sc_hd__and2b_1
XFILLER_119_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11161_ _11162_/A _11162_/B _11162_/C vssd1 vssd1 vccd1 vccd1 _11168_/A sky130_fd_sc_hd__a21oi_2
XFILLER_84_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10112_ _10112_/A _10234_/A vssd1 vssd1 vccd1 vccd1 _10119_/B sky130_fd_sc_hd__nor2_1
XFILLER_122_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11092_ _11092_/A _11092_/B vssd1 vssd1 vccd1 vccd1 _11104_/A sky130_fd_sc_hd__xnor2_1
XFILLER_121_135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14920_ _10062_/B _15003_/B _10111_/D _09981_/D _14914_/S _14958_/A vssd1 vssd1 vccd1
+ vccd1 _14920_/X sky130_fd_sc_hd__mux4_1
X_10043_ _14789_/A _10419_/B _10657_/B _12054_/B vssd1 vssd1 vccd1 vccd1 _10162_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_103_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14851_ _14851_/A _15463_/B vssd1 vssd1 vccd1 vccd1 _15541_/B sky130_fd_sc_hd__and2_1
XFILLER_21_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13802_ _14254_/A _13802_/B vssd1 vssd1 vccd1 vccd1 _13803_/B sky130_fd_sc_hd__nand2_1
XFILLER_29_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17570_ fanout935/X _17570_/D vssd1 vssd1 vccd1 vccd1 _17570_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14782_ _16136_/A _15811_/A vssd1 vssd1 vccd1 vccd1 _15801_/B sky130_fd_sc_hd__or2_1
X_11994_ _12155_/B _11993_/C _11993_/A vssd1 vssd1 vccd1 vccd1 _11994_/X sky130_fd_sc_hd__o21a_1
XFILLER_44_620 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16521_ _16522_/A _16522_/B vssd1 vssd1 vccd1 vccd1 _16625_/B sky130_fd_sc_hd__and2_1
XFILLER_28_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13733_ _14756_/A1 _13731_/Y _13828_/B _13630_/Y vssd1 vssd1 vccd1 vccd1 _17589_/D
+ sky130_fd_sc_hd__a31o_1
X_10945_ _10953_/A _10945_/B vssd1 vssd1 vccd1 vccd1 _10946_/C sky130_fd_sc_hd__and2_1
XFILLER_32_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_664 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16452_ _16453_/B _16453_/A vssd1 vssd1 vccd1 vccd1 _16452_/Y sky130_fd_sc_hd__nand2b_1
X_13664_ _13966_/A _14213_/B _13764_/D _13664_/D vssd1 vssd1 vccd1 vccd1 _13778_/A
+ sky130_fd_sc_hd__and4_1
X_10876_ _11122_/B _10875_/C _10962_/B _10933_/A vssd1 vssd1 vccd1 vccd1 _10876_/Y
+ sky130_fd_sc_hd__a22oi_1
X_15403_ _16127_/A _16533_/A _15484_/A vssd1 vssd1 vccd1 vccd1 _15403_/X sky130_fd_sc_hd__and3_1
X_12615_ _12474_/A _12474_/B _12472_/Y vssd1 vssd1 vccd1 vccd1 _12629_/A sky130_fd_sc_hd__a21bo_1
X_16383_ _16292_/B _16562_/B _16562_/C vssd1 vssd1 vccd1 vccd1 _16385_/B sky130_fd_sc_hd__o21a_1
X_13595_ _13595_/A _13595_/B vssd1 vssd1 vccd1 vccd1 _13597_/B sky130_fd_sc_hd__xnor2_1
XFILLER_84_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15334_ _15334_/A _15334_/B vssd1 vssd1 vccd1 vccd1 _15337_/B sky130_fd_sc_hd__xor2_1
X_12546_ _12845_/S _12700_/B _12546_/C vssd1 vssd1 vccd1 vccd1 _12548_/B sky130_fd_sc_hd__and3_1
XFILLER_118_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15265_ _14899_/X _14968_/X _16446_/A _11675_/B vssd1 vssd1 vccd1 vccd1 _15331_/A
+ sky130_fd_sc_hd__a211o_1
X_12477_ _12477_/A _12477_/B vssd1 vssd1 vccd1 vccd1 _12478_/B sky130_fd_sc_hd__nor2_1
X_17004_ _17090_/A _17004_/B vssd1 vssd1 vccd1 vccd1 _17007_/A sky130_fd_sc_hd__nand2_1
XANTENNA_4 _17493_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14216_ _14216_/A _14216_/B vssd1 vssd1 vccd1 vccd1 _14218_/C sky130_fd_sc_hd__xnor2_1
X_11428_ _11553_/B _11563_/D vssd1 vssd1 vccd1 vccd1 _11430_/B sky130_fd_sc_hd__nand2_1
X_15196_ _17306_/A1 _17162_/C1 _15195_/X vssd1 vssd1 vccd1 vccd1 _17547_/D sky130_fd_sc_hd__a21oi_1
X_11359_ _11359_/A _11359_/B vssd1 vssd1 vccd1 vccd1 _11413_/B sky130_fd_sc_hd__and2_1
X_14147_ _14148_/A _14148_/B vssd1 vssd1 vccd1 vccd1 _14221_/B sky130_fd_sc_hd__and2b_1
XFILLER_113_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14078_ _14188_/A _14078_/B vssd1 vssd1 vccd1 vccd1 _14098_/A sky130_fd_sc_hd__nand2_1
XFILLER_140_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13029_ _13029_/A _13029_/B vssd1 vssd1 vccd1 vccd1 _13031_/B sky130_fd_sc_hd__xnor2_1
XFILLER_6_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_745 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16719_ _16715_/Y _16717_/Y _16718_/Y vssd1 vssd1 vccd1 vccd1 _16719_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_23_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09122_ _09122_/A _09122_/B vssd1 vssd1 vccd1 vccd1 _09256_/A sky130_fd_sc_hd__nor2_1
XFILLER_148_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09053_ _09053_/A _09053_/B vssd1 vssd1 vccd1 vccd1 _09055_/C sky130_fd_sc_hd__or2_1
XFILLER_108_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09955_ _09956_/A _09956_/B vssd1 vssd1 vccd1 vccd1 _09957_/A sky130_fd_sc_hd__nand2_1
XFILLER_106_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08906_ _08905_/A _09051_/A _08832_/Y _08875_/X vssd1 vssd1 vccd1 vccd1 _08930_/A
+ sky130_fd_sc_hd__a211oi_4
XFILLER_98_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09886_ _09914_/B _10029_/A _09914_/A vssd1 vssd1 vccd1 vccd1 _09915_/A sky130_fd_sc_hd__o21a_1
XFILLER_106_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08837_ _08835_/Y _08862_/A _09730_/C _11900_/D vssd1 vssd1 vccd1 vccd1 _08862_/B
+ sky130_fd_sc_hd__and4bb_1
XFILLER_57_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08768_ _08768_/A _08768_/B vssd1 vssd1 vccd1 vccd1 _08780_/A sky130_fd_sc_hd__nor2_1
XTAP_2726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10730_ _11212_/A _11212_/B vssd1 vssd1 vccd1 vccd1 _10730_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_26_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10661_ _10661_/A _10669_/B vssd1 vssd1 vccd1 vccd1 _10662_/C sky130_fd_sc_hd__xnor2_1
XFILLER_9_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12400_ _17164_/A _12400_/B vssd1 vssd1 vccd1 vccd1 _12401_/B sky130_fd_sc_hd__or2_1
XFILLER_167_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13380_ _13500_/B _13378_/X _13252_/Y _13256_/A vssd1 vssd1 vccd1 vccd1 _13380_/X
+ sky130_fd_sc_hd__o211a_1
X_10592_ _10592_/A vssd1 vssd1 vccd1 vccd1 _10593_/B sky130_fd_sc_hd__inv_2
XFILLER_51_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12331_ _12333_/A vssd1 vssd1 vccd1 vccd1 _12331_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_30 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15050_ _14796_/A _14796_/B _14796_/C _14796_/D vssd1 vssd1 vccd1 vccd1 _15050_/X
+ sky130_fd_sc_hd__a22o_1
X_12262_ _12263_/A _12263_/B vssd1 vssd1 vccd1 vccd1 _12454_/B sky130_fd_sc_hd__nand2b_1
XFILLER_135_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11213_ _11181_/A _11181_/B _11182_/Y vssd1 vssd1 vccd1 vccd1 _11216_/B sky130_fd_sc_hd__a21o_1
XFILLER_123_912 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14001_ _14001_/A _14001_/B vssd1 vssd1 vccd1 vccd1 _14002_/C sky130_fd_sc_hd__xor2_1
XFILLER_107_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12193_ _12360_/A _12193_/B _12193_/C vssd1 vssd1 vccd1 vccd1 _12360_/B sky130_fd_sc_hd__nand3_1
XFILLER_107_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11144_ _11144_/A _11237_/A vssd1 vssd1 vccd1 vccd1 _11145_/C sky130_fd_sc_hd__nand2_1
Xoutput74 _17467_/Q vssd1 vssd1 vccd1 vccd1 leds[1] sky130_fd_sc_hd__clkbuf_1
Xoutput85 _17444_/Q vssd1 vssd1 vccd1 vccd1 o_wb_data[10] sky130_fd_sc_hd__clkbuf_1
XFILLER_163_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput96 _17454_/Q vssd1 vssd1 vccd1 vccd1 o_wb_data[20] sky130_fd_sc_hd__clkbuf_1
XFILLER_89_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11075_ _11075_/A _11075_/B _11075_/C vssd1 vssd1 vccd1 vccd1 _11110_/A sky130_fd_sc_hd__or3_1
X_15952_ _15953_/A _15953_/B vssd1 vssd1 vccd1 vccd1 _15954_/A sky130_fd_sc_hd__or2_1
XFILLER_1_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14903_ _14879_/Y _15205_/A _14900_/X _08731_/A _14877_/Y vssd1 vssd1 vccd1 vccd1
+ _14903_/X sky130_fd_sc_hd__a2111o_1
XFILLER_0_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10026_ _09865_/B _09975_/X _09991_/Y _10005_/X vssd1 vssd1 vccd1 vccd1 _10027_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_49_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15883_ _15883_/A _15883_/B _15881_/Y vssd1 vssd1 vccd1 vccd1 _15884_/B sky130_fd_sc_hd__or3b_1
XFILLER_64_726 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14834_ _17477_/D _17476_/D vssd1 vssd1 vccd1 vccd1 _14938_/B sky130_fd_sc_hd__nand2b_1
XFILLER_63_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17553_ fanout940/X _17553_/D vssd1 vssd1 vccd1 vccd1 _17553_/Q sky130_fd_sc_hd__dfxtp_1
X_14765_ _14765_/A _14765_/B vssd1 vssd1 vccd1 vccd1 _14765_/X sky130_fd_sc_hd__or2_1
XFILLER_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11977_ _12804_/A _17417_/A _12174_/D _12129_/B vssd1 vssd1 vccd1 vccd1 _11978_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_44_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16504_ _16503_/Y _16504_/B vssd1 vssd1 vccd1 vccd1 _16504_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_60_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13716_ _13818_/A _13714_/Y _13601_/A _13604_/A vssd1 vssd1 vccd1 vccd1 _13717_/B
+ sky130_fd_sc_hd__a211o_1
X_10928_ _11074_/A _10928_/B vssd1 vssd1 vccd1 vccd1 _11057_/C sky130_fd_sc_hd__xnor2_1
X_17484_ fanout948/X _17484_/D vssd1 vssd1 vccd1 vccd1 _17484_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_44_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14696_ _14698_/A _14699_/A vssd1 vssd1 vccd1 vccd1 _14727_/A sky130_fd_sc_hd__nor2_1
XFILLER_108_1015 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16435_ _16436_/B _16436_/A vssd1 vssd1 vccd1 vccd1 _16435_/X sky130_fd_sc_hd__and2b_1
XFILLER_108_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13647_ _13529_/B _13535_/B _13527_/X vssd1 vssd1 vccd1 vccd1 _13648_/C sky130_fd_sc_hd__a21o_1
XFILLER_32_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10859_ _10859_/A _10859_/B _10859_/C vssd1 vssd1 vccd1 vccd1 _10861_/B sky130_fd_sc_hd__nand3_1
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16366_ _16367_/A _16367_/B vssd1 vssd1 vccd1 vccd1 _16462_/B sky130_fd_sc_hd__nor2_1
XFILLER_9_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13578_ _13578_/A _16859_/A vssd1 vssd1 vccd1 vccd1 _13579_/B sky130_fd_sc_hd__nand2_1
XFILLER_157_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15317_ _11100_/A _14931_/X _15316_/X _16977_/A vssd1 vssd1 vccd1 vccd1 _15317_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_9_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12529_ _12528_/A _12528_/B _12528_/C vssd1 vssd1 vccd1 vccd1 _12530_/B sky130_fd_sc_hd__o21a_1
XFILLER_118_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16297_ _14777_/A _16644_/B _16298_/A vssd1 vssd1 vccd1 vccd1 _16394_/A sky130_fd_sc_hd__a21bo_1
XFILLER_117_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15248_ _15314_/B _15248_/B _15248_/C vssd1 vssd1 vccd1 vccd1 _15257_/B sky130_fd_sc_hd__and3b_1
XFILLER_173_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15179_ _14950_/X _14955_/X _15312_/S vssd1 vssd1 vccd1 vccd1 _15179_/X sky130_fd_sc_hd__mux2_1
XFILLER_153_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout308 _15175_/A vssd1 vssd1 vccd1 vccd1 _14733_/S sky130_fd_sc_hd__buf_2
XFILLER_28_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout319 _14832_/A vssd1 vssd1 vccd1 vccd1 _14213_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_114_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09740_ _09740_/A _09740_/B _09740_/C vssd1 vssd1 vccd1 vccd1 _09832_/A sky130_fd_sc_hd__and3_1
XFILLER_100_116 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
.ends

