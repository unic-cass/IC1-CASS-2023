magic
tech sky130B
magscale 1 2
timestamp 1676037725
use sky130_fd_pr__hvdfl1sd__example_55959141808418  sky130_fd_pr__hvdfl1sd__example_55959141808418_0
timestamp 1676037725
transform -1 0 295 0 -1 682
box 0 0 1 1
use sky130_fd_pr__model__nfet_highvoltage__example_55959141808419  sky130_fd_pr__model__nfet_highvoltage__example_55959141808419_0
timestamp 1676037725
transform 1 0 119 0 -1 284
box -1 0 297 1
use sky130_fd_pr__model__pfet_highvoltage__example_55959141808420  sky130_fd_pr__model__pfet_highvoltage__example_55959141808420_0
timestamp 1676037725
transform -1 0 415 0 -1 682
box -1 0 0 1
use sky130_fd_pr__model__pfet_highvoltage__example_55959141808420  sky130_fd_pr__model__pfet_highvoltage__example_55959141808420_1
timestamp 1676037725
transform 1 0 119 0 -1 682
box -1 0 0 1
use sky130_fd_pr__model__pfet_highvoltage__example_55959141808421  sky130_fd_pr__model__pfet_highvoltage__example_55959141808421_0
timestamp 1676037725
transform 1 0 119 0 1 750
box -1 0 297 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_0
timestamp 1676037725
transform 0 -1 460 -1 0 227
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_1
timestamp 1676037725
transform 0 -1 108 1 0 872
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_2
timestamp 1676037725
transform 0 -1 108 -1 0 227
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_0
timestamp 1676037725
transform 0 -1 390 1 0 316
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_1
timestamp 1676037725
transform 0 -1 212 1 0 316
box 0 0 1 1
<< properties >>
string GDS_END 30058908
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 30056780
<< end >>
