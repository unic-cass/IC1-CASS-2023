magic
tech sky130A
magscale 1 2
timestamp 1676037725
<< pwell >>
rect 761 765 776 783
<< metal1 >>
rect -88 1562 1628 1568
rect -88 1510 -12 1562
rect 40 1510 52 1562
rect 104 1510 116 1562
rect 168 1510 180 1562
rect 232 1510 244 1562
rect 296 1510 308 1562
rect 360 1510 372 1562
rect 424 1510 436 1562
rect 488 1510 500 1562
rect 552 1510 564 1562
rect 616 1510 628 1562
rect 680 1510 692 1562
rect 744 1510 756 1562
rect 808 1510 820 1562
rect 872 1510 884 1562
rect 936 1510 948 1562
rect 1000 1510 1012 1562
rect 1064 1510 1076 1562
rect 1128 1510 1140 1562
rect 1192 1510 1204 1562
rect 1256 1510 1268 1562
rect 1320 1510 1332 1562
rect 1384 1510 1396 1562
rect 1448 1510 1460 1562
rect 1512 1510 1524 1562
rect 1576 1510 1628 1562
rect -88 1504 1628 1510
rect -88 1449 -34 1476
rect -88 1397 -87 1449
rect -35 1397 -34 1449
rect -88 1385 -34 1397
rect -88 1333 -87 1385
rect -35 1333 -34 1385
rect -88 1321 -34 1333
rect -88 1269 -87 1321
rect -35 1269 -34 1321
rect -88 1257 -34 1269
rect -88 1205 -87 1257
rect -35 1205 -34 1257
rect -88 1193 -34 1205
rect -88 1141 -87 1193
rect -35 1141 -34 1193
rect -88 1129 -34 1141
rect -88 1077 -87 1129
rect -35 1077 -34 1129
rect -88 1065 -34 1077
rect -88 1013 -87 1065
rect -35 1013 -34 1065
rect -88 1001 -34 1013
rect -88 949 -87 1001
rect -35 949 -34 1001
rect -88 937 -34 949
rect -88 885 -87 937
rect -35 885 -34 937
rect -88 873 -34 885
rect -88 821 -87 873
rect -35 821 -34 873
rect -88 809 -34 821
rect -88 757 -87 809
rect -35 757 -34 809
rect -88 745 -34 757
rect -88 693 -87 745
rect -35 693 -34 745
rect -88 681 -34 693
rect -88 629 -87 681
rect -35 629 -34 681
rect -88 617 -34 629
rect -88 565 -87 617
rect -35 565 -34 617
rect -88 553 -34 565
rect -88 501 -87 553
rect -35 501 -34 553
rect -88 489 -34 501
rect -88 437 -87 489
rect -35 437 -34 489
rect -88 425 -34 437
rect -88 373 -87 425
rect -35 373 -34 425
rect -88 361 -34 373
rect -88 309 -87 361
rect -35 309 -34 361
rect -88 297 -34 309
rect -88 245 -87 297
rect -35 245 -34 297
rect -88 233 -34 245
rect -88 181 -87 233
rect -35 181 -34 233
rect -88 169 -34 181
rect -88 117 -87 169
rect -35 117 -34 169
rect -88 105 -34 117
rect -88 53 -87 105
rect -35 64 -34 105
rect 0 64 28 1476
rect 56 92 84 1504
rect 112 64 140 1476
rect 168 92 196 1504
rect 224 64 252 1476
rect 280 92 308 1504
rect 336 64 364 1476
rect 392 92 420 1504
rect 448 64 476 1476
rect 504 92 532 1504
rect 560 64 588 1476
rect 616 92 644 1504
rect 672 64 700 1476
rect 728 92 756 1504
rect 784 64 812 1476
rect 840 92 868 1504
rect 896 64 924 1476
rect 952 92 980 1504
rect 1008 64 1036 1476
rect 1064 92 1092 1504
rect 1120 64 1148 1476
rect 1176 92 1204 1504
rect 1232 64 1260 1476
rect 1288 92 1316 1504
rect 1344 64 1372 1476
rect 1400 92 1428 1504
rect 1456 64 1484 1476
rect 1512 92 1540 1504
rect 1574 1494 1628 1504
rect 1574 1442 1575 1494
rect 1627 1442 1628 1494
rect 1574 1430 1628 1442
rect 1574 1378 1575 1430
rect 1627 1378 1628 1430
rect 1574 1366 1628 1378
rect 1574 1314 1575 1366
rect 1627 1314 1628 1366
rect 1574 1302 1628 1314
rect 1574 1250 1575 1302
rect 1627 1250 1628 1302
rect 1574 1238 1628 1250
rect 1574 1186 1575 1238
rect 1627 1186 1628 1238
rect 1574 1174 1628 1186
rect 1574 1122 1575 1174
rect 1627 1122 1628 1174
rect 1574 1110 1628 1122
rect 1574 1058 1575 1110
rect 1627 1058 1628 1110
rect 1574 1046 1628 1058
rect 1574 994 1575 1046
rect 1627 994 1628 1046
rect 1574 982 1628 994
rect 1574 930 1575 982
rect 1627 930 1628 982
rect 1574 918 1628 930
rect 1574 866 1575 918
rect 1627 866 1628 918
rect 1574 854 1628 866
rect 1574 802 1575 854
rect 1627 802 1628 854
rect 1574 790 1628 802
rect 1574 738 1575 790
rect 1627 738 1628 790
rect 1574 726 1628 738
rect 1574 674 1575 726
rect 1627 674 1628 726
rect 1574 662 1628 674
rect 1574 610 1575 662
rect 1627 610 1628 662
rect 1574 598 1628 610
rect 1574 546 1575 598
rect 1627 546 1628 598
rect 1574 534 1628 546
rect 1574 482 1575 534
rect 1627 482 1628 534
rect 1574 470 1628 482
rect 1574 418 1575 470
rect 1627 418 1628 470
rect 1574 406 1628 418
rect 1574 354 1575 406
rect 1627 354 1628 406
rect 1574 342 1628 354
rect 1574 290 1575 342
rect 1627 290 1628 342
rect 1574 278 1628 290
rect 1574 226 1575 278
rect 1627 226 1628 278
rect 1574 214 1628 226
rect 1574 162 1575 214
rect 1627 162 1628 214
rect 1574 150 1628 162
rect 1574 98 1575 150
rect 1627 98 1628 150
rect 1574 92 1628 98
rect -35 58 1628 64
rect -35 53 -12 58
rect -88 6 -12 53
rect 40 6 52 58
rect 104 6 116 58
rect 168 6 180 58
rect 232 6 244 58
rect 296 6 308 58
rect 360 6 372 58
rect 424 6 436 58
rect 488 6 500 58
rect 552 6 564 58
rect 616 6 628 58
rect 680 6 692 58
rect 744 6 756 58
rect 808 6 820 58
rect 872 6 884 58
rect 936 6 948 58
rect 1000 6 1012 58
rect 1064 6 1076 58
rect 1128 6 1140 58
rect 1192 6 1204 58
rect 1256 6 1268 58
rect 1320 6 1332 58
rect 1384 6 1396 58
rect 1448 6 1460 58
rect 1512 6 1524 58
rect 1576 6 1628 58
rect -88 0 1628 6
<< via1 >>
rect -12 1510 40 1562
rect 52 1510 104 1562
rect 116 1510 168 1562
rect 180 1510 232 1562
rect 244 1510 296 1562
rect 308 1510 360 1562
rect 372 1510 424 1562
rect 436 1510 488 1562
rect 500 1510 552 1562
rect 564 1510 616 1562
rect 628 1510 680 1562
rect 692 1510 744 1562
rect 756 1510 808 1562
rect 820 1510 872 1562
rect 884 1510 936 1562
rect 948 1510 1000 1562
rect 1012 1510 1064 1562
rect 1076 1510 1128 1562
rect 1140 1510 1192 1562
rect 1204 1510 1256 1562
rect 1268 1510 1320 1562
rect 1332 1510 1384 1562
rect 1396 1510 1448 1562
rect 1460 1510 1512 1562
rect 1524 1510 1576 1562
rect -87 1397 -35 1449
rect -87 1333 -35 1385
rect -87 1269 -35 1321
rect -87 1205 -35 1257
rect -87 1141 -35 1193
rect -87 1077 -35 1129
rect -87 1013 -35 1065
rect -87 949 -35 1001
rect -87 885 -35 937
rect -87 821 -35 873
rect -87 757 -35 809
rect -87 693 -35 745
rect -87 629 -35 681
rect -87 565 -35 617
rect -87 501 -35 553
rect -87 437 -35 489
rect -87 373 -35 425
rect -87 309 -35 361
rect -87 245 -35 297
rect -87 181 -35 233
rect -87 117 -35 169
rect -87 53 -35 105
rect 1575 1442 1627 1494
rect 1575 1378 1627 1430
rect 1575 1314 1627 1366
rect 1575 1250 1627 1302
rect 1575 1186 1627 1238
rect 1575 1122 1627 1174
rect 1575 1058 1627 1110
rect 1575 994 1627 1046
rect 1575 930 1627 982
rect 1575 866 1627 918
rect 1575 802 1627 854
rect 1575 738 1627 790
rect 1575 674 1627 726
rect 1575 610 1627 662
rect 1575 546 1627 598
rect 1575 482 1627 534
rect 1575 418 1627 470
rect 1575 354 1627 406
rect 1575 290 1627 342
rect 1575 226 1627 278
rect 1575 162 1627 214
rect 1575 98 1627 150
rect -12 6 40 58
rect 52 6 104 58
rect 116 6 168 58
rect 180 6 232 58
rect 244 6 296 58
rect 308 6 360 58
rect 372 6 424 58
rect 436 6 488 58
rect 500 6 552 58
rect 564 6 616 58
rect 628 6 680 58
rect 692 6 744 58
rect 756 6 808 58
rect 820 6 872 58
rect 884 6 936 58
rect 948 6 1000 58
rect 1012 6 1064 58
rect 1076 6 1128 58
rect 1140 6 1192 58
rect 1204 6 1256 58
rect 1268 6 1320 58
rect 1332 6 1384 58
rect 1396 6 1448 58
rect 1460 6 1512 58
rect 1524 6 1576 58
<< metal2 >>
rect -88 1562 1628 1568
rect -88 1510 -12 1562
rect 40 1510 52 1562
rect 104 1510 116 1562
rect 168 1510 180 1562
rect 232 1510 244 1562
rect 296 1510 308 1562
rect 360 1510 372 1562
rect 424 1510 436 1562
rect 488 1510 500 1562
rect 552 1510 564 1562
rect 616 1510 628 1562
rect 680 1510 692 1562
rect 744 1510 756 1562
rect 808 1510 820 1562
rect 872 1510 884 1562
rect 936 1510 948 1562
rect 1000 1510 1012 1562
rect 1064 1510 1076 1562
rect 1128 1510 1140 1562
rect 1192 1510 1204 1562
rect 1256 1510 1268 1562
rect 1320 1510 1332 1562
rect 1384 1510 1396 1562
rect 1448 1510 1460 1562
rect 1512 1510 1524 1562
rect 1576 1510 1628 1562
rect -88 1504 1628 1510
rect -88 1449 -34 1476
rect -88 1397 -87 1449
rect -35 1397 -34 1449
rect -88 1385 -34 1397
rect -88 1333 -87 1385
rect -35 1333 -34 1385
rect -88 1321 -34 1333
rect -88 1269 -87 1321
rect -35 1269 -34 1321
rect -88 1257 -34 1269
rect -88 1205 -87 1257
rect -35 1205 -34 1257
rect -88 1193 -34 1205
rect -88 1141 -87 1193
rect -35 1141 -34 1193
rect -88 1129 -34 1141
rect -88 1077 -87 1129
rect -35 1077 -34 1129
rect -88 1065 -34 1077
rect -88 1013 -87 1065
rect -35 1013 -34 1065
rect -88 1001 -34 1013
rect -88 949 -87 1001
rect -35 949 -34 1001
rect -88 937 -34 949
rect -88 885 -87 937
rect -35 885 -34 937
rect -88 873 -34 885
rect -88 821 -87 873
rect -35 821 -34 873
rect -88 809 -34 821
rect -88 757 -87 809
rect -35 757 -34 809
rect -88 745 -34 757
rect -88 693 -87 745
rect -35 693 -34 745
rect -88 681 -34 693
rect -88 629 -87 681
rect -35 629 -34 681
rect -88 617 -34 629
rect -88 565 -87 617
rect -35 565 -34 617
rect -88 553 -34 565
rect -88 501 -87 553
rect -35 501 -34 553
rect -88 489 -34 501
rect -88 437 -87 489
rect -35 437 -34 489
rect -88 425 -34 437
rect -88 373 -87 425
rect -35 373 -34 425
rect -88 361 -34 373
rect -88 309 -87 361
rect -35 309 -34 361
rect -88 297 -34 309
rect -88 245 -87 297
rect -35 245 -34 297
rect -88 233 -34 245
rect -88 181 -87 233
rect -35 181 -34 233
rect -88 169 -34 181
rect -88 117 -87 169
rect -35 117 -34 169
rect -88 105 -34 117
rect -88 53 -87 105
rect -35 64 -34 105
rect 0 92 28 1504
rect 56 64 84 1476
rect 112 92 140 1504
rect 168 64 196 1476
rect 224 92 252 1504
rect 280 64 308 1476
rect 336 92 364 1504
rect 392 64 420 1476
rect 448 92 476 1504
rect 504 64 532 1476
rect 560 92 588 1504
rect 616 64 644 1476
rect 672 92 700 1504
rect 728 64 756 1476
rect 784 92 812 1504
rect 840 64 868 1476
rect 896 92 924 1504
rect 952 64 980 1476
rect 1008 92 1036 1504
rect 1064 64 1092 1476
rect 1120 92 1148 1504
rect 1176 64 1204 1476
rect 1232 92 1260 1504
rect 1288 64 1316 1476
rect 1344 92 1372 1504
rect 1400 64 1428 1476
rect 1456 92 1484 1504
rect 1574 1494 1628 1504
rect 1512 64 1540 1476
rect 1574 1442 1575 1494
rect 1627 1442 1628 1494
rect 1574 1430 1628 1442
rect 1574 1378 1575 1430
rect 1627 1378 1628 1430
rect 1574 1366 1628 1378
rect 1574 1314 1575 1366
rect 1627 1314 1628 1366
rect 1574 1302 1628 1314
rect 1574 1250 1575 1302
rect 1627 1250 1628 1302
rect 1574 1238 1628 1250
rect 1574 1186 1575 1238
rect 1627 1186 1628 1238
rect 1574 1174 1628 1186
rect 1574 1122 1575 1174
rect 1627 1122 1628 1174
rect 1574 1110 1628 1122
rect 1574 1058 1575 1110
rect 1627 1058 1628 1110
rect 1574 1046 1628 1058
rect 1574 994 1575 1046
rect 1627 994 1628 1046
rect 1574 982 1628 994
rect 1574 930 1575 982
rect 1627 930 1628 982
rect 1574 918 1628 930
rect 1574 866 1575 918
rect 1627 866 1628 918
rect 1574 854 1628 866
rect 1574 802 1575 854
rect 1627 802 1628 854
rect 1574 790 1628 802
rect 1574 738 1575 790
rect 1627 738 1628 790
rect 1574 726 1628 738
rect 1574 674 1575 726
rect 1627 674 1628 726
rect 1574 662 1628 674
rect 1574 610 1575 662
rect 1627 610 1628 662
rect 1574 598 1628 610
rect 1574 546 1575 598
rect 1627 546 1628 598
rect 1574 534 1628 546
rect 1574 482 1575 534
rect 1627 482 1628 534
rect 1574 470 1628 482
rect 1574 418 1575 470
rect 1627 418 1628 470
rect 1574 406 1628 418
rect 1574 354 1575 406
rect 1627 354 1628 406
rect 1574 342 1628 354
rect 1574 290 1575 342
rect 1627 290 1628 342
rect 1574 278 1628 290
rect 1574 226 1575 278
rect 1627 226 1628 278
rect 1574 214 1628 226
rect 1574 162 1575 214
rect 1627 162 1628 214
rect 1574 150 1628 162
rect 1574 98 1575 150
rect 1627 98 1628 150
rect 1574 92 1628 98
rect -35 58 1628 64
rect -35 53 -12 58
rect -88 6 -12 53
rect 40 6 52 58
rect 104 6 116 58
rect 168 6 180 58
rect 232 6 244 58
rect 296 6 308 58
rect 360 6 372 58
rect 424 6 436 58
rect 488 6 500 58
rect 552 6 564 58
rect 616 6 628 58
rect 680 6 692 58
rect 744 6 756 58
rect 808 6 820 58
rect 872 6 884 58
rect 936 6 948 58
rect 1000 6 1012 58
rect 1064 6 1076 58
rect 1128 6 1140 58
rect 1192 6 1204 58
rect 1256 6 1268 58
rect 1320 6 1332 58
rect 1384 6 1396 58
rect 1448 6 1460 58
rect 1512 6 1524 58
rect 1576 6 1628 58
rect -88 0 1628 6
<< labels >>
flabel comment s 735 33 735 33 0 FreeSans 200 0 0 0 For future design recommend using caps in MTM-378
flabel metal2 s 674 1373 697 1400 0 FreeSans 200 0 0 0 C1
port 2 nsew
flabel metal2 s 729 133 754 161 0 FreeSans 200 0 0 0 C0
port 1 nsew
flabel pwell s 761 765 776 783 0 FreeSans 200 0 0 0 SUB
port 3 nsew
<< properties >>
string GDS_END 304028
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 291758
string device primitive
<< end >>
