magic
tech sky130B
magscale 1 2
timestamp 1676037725
<< nwell >>
rect 2539 436 3101 1168
<< pwell >>
rect 1744 -1391 1996 -909
<< mvnmos >>
rect 1770 -1122 1970 -1002
rect 1770 -1298 1970 -1178
<< mvpmos >>
rect 2672 502 2792 1102
rect 2848 502 2968 1102
<< mvndiff >>
rect 1770 -943 1970 -935
rect 1770 -977 1782 -943
rect 1816 -977 1850 -943
rect 1884 -977 1918 -943
rect 1952 -977 1970 -943
rect 1770 -1002 1970 -977
rect 1770 -1133 1970 -1122
rect 1770 -1167 1782 -1133
rect 1816 -1167 1850 -1133
rect 1884 -1167 1918 -1133
rect 1952 -1167 1970 -1133
rect 1770 -1178 1970 -1167
rect 1770 -1323 1970 -1298
rect 1770 -1357 1782 -1323
rect 1816 -1357 1850 -1323
rect 1884 -1357 1918 -1323
rect 1952 -1357 1970 -1323
rect 1770 -1365 1970 -1357
<< mvpdiff >>
rect 2605 1090 2672 1102
rect 2605 1056 2613 1090
rect 2647 1056 2672 1090
rect 2605 1022 2672 1056
rect 2605 988 2613 1022
rect 2647 988 2672 1022
rect 2605 954 2672 988
rect 2605 920 2613 954
rect 2647 920 2672 954
rect 2605 886 2672 920
rect 2605 852 2613 886
rect 2647 852 2672 886
rect 2605 818 2672 852
rect 2605 784 2613 818
rect 2647 784 2672 818
rect 2605 750 2672 784
rect 2605 716 2613 750
rect 2647 716 2672 750
rect 2605 682 2672 716
rect 2605 648 2613 682
rect 2647 648 2672 682
rect 2605 614 2672 648
rect 2605 580 2613 614
rect 2647 580 2672 614
rect 2605 502 2672 580
rect 2792 502 2848 1102
rect 2968 1090 3035 1102
rect 2968 1056 2993 1090
rect 3027 1056 3035 1090
rect 2968 1022 3035 1056
rect 2968 988 2993 1022
rect 3027 988 3035 1022
rect 2968 954 3035 988
rect 2968 920 2993 954
rect 3027 920 3035 954
rect 2968 886 3035 920
rect 2968 852 2993 886
rect 3027 852 3035 886
rect 2968 818 3035 852
rect 2968 784 2993 818
rect 3027 784 3035 818
rect 2968 750 3035 784
rect 2968 716 2993 750
rect 3027 716 3035 750
rect 2968 682 3035 716
rect 2968 648 2993 682
rect 3027 648 3035 682
rect 2968 614 3035 648
rect 2968 580 2993 614
rect 3027 580 3035 614
rect 2968 502 3035 580
<< mvndiffc >>
rect 1782 -977 1816 -943
rect 1850 -977 1884 -943
rect 1918 -977 1952 -943
rect 1782 -1167 1816 -1133
rect 1850 -1167 1884 -1133
rect 1918 -1167 1952 -1133
rect 1782 -1357 1816 -1323
rect 1850 -1357 1884 -1323
rect 1918 -1357 1952 -1323
<< mvpdiffc >>
rect 2613 1056 2647 1090
rect 2613 988 2647 1022
rect 2613 920 2647 954
rect 2613 852 2647 886
rect 2613 784 2647 818
rect 2613 716 2647 750
rect 2613 648 2647 682
rect 2613 580 2647 614
rect 2993 1056 3027 1090
rect 2993 988 3027 1022
rect 2993 920 3027 954
rect 2993 852 3027 886
rect 2993 784 3027 818
rect 2993 716 3027 750
rect 2993 648 3027 682
rect 2993 580 3027 614
<< poly >>
rect 2672 1102 2792 1128
rect 2848 1102 2968 1128
rect 2672 454 2792 502
rect 2672 420 2715 454
rect 2749 420 2792 454
rect 2672 386 2792 420
rect 2672 352 2715 386
rect 2749 352 2792 386
rect 2672 340 2792 352
rect 2848 454 2968 502
rect 2848 420 2891 454
rect 2925 420 2968 454
rect 2848 386 2968 420
rect 2848 352 2891 386
rect 2925 352 2968 386
rect 2848 340 2968 352
rect 2699 336 2765 340
rect 2875 336 2941 340
rect 1744 -1122 1770 -1002
rect 1970 -1047 2140 -1002
rect 1970 -1081 2018 -1047
rect 2052 -1081 2086 -1047
rect 2120 -1081 2140 -1047
rect 1970 -1122 2140 -1081
rect 1744 -1298 1770 -1178
rect 1970 -1229 2140 -1178
rect 1970 -1263 2018 -1229
rect 2052 -1263 2086 -1229
rect 2120 -1263 2140 -1229
rect 1970 -1298 2140 -1263
<< polycont >>
rect 2715 420 2749 454
rect 2715 352 2749 386
rect 2891 420 2925 454
rect 2891 352 2925 386
rect 2018 -1081 2052 -1047
rect 2086 -1081 2120 -1047
rect 2018 -1263 2052 -1229
rect 2086 -1263 2120 -1229
<< locali >>
rect 2613 1090 2647 1125
rect 2613 1022 2647 1053
rect 2613 954 2647 981
rect 2613 886 2647 920
rect 2613 818 2647 852
rect 2613 750 2647 784
rect 2613 682 2647 716
rect 2613 614 2647 648
rect 2613 564 2647 580
rect 2993 1090 3077 1107
rect 3027 1056 3077 1090
rect 2993 1022 3077 1056
rect 3027 988 3077 1022
rect 2993 954 3077 988
rect 3027 920 3077 954
rect 2993 886 3077 920
rect 3027 852 3077 886
rect 2993 818 3077 852
rect 3027 784 3077 818
rect 2993 750 3077 784
rect 3027 716 3077 750
rect 2993 682 3077 716
rect 3027 648 3077 682
rect 2993 614 3077 648
rect 3027 580 3077 614
rect 2993 463 3077 580
rect 2699 420 2715 454
rect 2749 442 2765 454
rect 2699 408 2717 420
rect 2751 408 2765 442
rect 2699 386 2765 408
rect 2699 352 2715 386
rect 2749 370 2765 386
rect 2751 352 2765 370
rect 2875 420 2891 454
rect 2925 442 2941 454
rect 2875 408 2899 420
rect 2933 408 2941 442
rect 2875 386 2941 408
rect 2875 352 2891 386
rect 2925 370 2941 386
rect 2933 352 2941 370
rect 2993 328 3211 463
rect 1766 -977 1782 -943
rect 1816 -977 1850 -943
rect 1884 -977 1918 -943
rect 1956 -977 1968 -943
rect 2002 -1081 2018 -1047
rect 2055 -1081 2086 -1047
rect 2127 -1081 2136 -1047
rect 1766 -1167 1782 -1133
rect 1816 -1167 1850 -1133
rect 1884 -1167 1918 -1133
rect 1952 -1167 1968 -1133
rect 2002 -1263 2018 -1229
rect 2055 -1263 2086 -1229
rect 2127 -1263 2136 -1229
rect 1766 -1357 1782 -1323
rect 1816 -1357 1850 -1323
rect 1884 -1357 1918 -1323
rect 1952 -1357 1968 -1323
<< viali >>
rect 2613 1125 2647 1159
rect 2613 1056 2647 1087
rect 2613 1053 2647 1056
rect 2613 988 2647 1015
rect 2613 981 2647 988
rect 2717 420 2749 442
rect 2749 420 2751 442
rect 2717 408 2751 420
rect 2717 352 2749 370
rect 2749 352 2751 370
rect 2899 420 2925 442
rect 2925 420 2933 442
rect 2899 408 2933 420
rect 2899 352 2925 370
rect 2925 352 2933 370
rect 2717 336 2751 352
rect 2899 336 2933 352
rect 1850 -977 1884 -943
rect 1922 -977 1952 -943
rect 1952 -977 1956 -943
rect 2021 -1081 2052 -1047
rect 2052 -1081 2055 -1047
rect 2093 -1081 2120 -1047
rect 2120 -1081 2127 -1047
rect 2021 -1263 2052 -1229
rect 2052 -1263 2055 -1229
rect 2093 -1263 2120 -1229
rect 2120 -1263 2127 -1229
<< metal1 >>
rect 2571 1159 3078 1172
rect 2571 1125 2613 1159
rect 2647 1125 3078 1159
rect 2571 1087 3078 1125
rect 2571 1053 2613 1087
rect 2647 1053 3078 1087
rect 2571 1015 3078 1053
rect 2571 981 2613 1015
rect 2647 981 3078 1015
rect 2571 969 3078 981
rect 2711 442 2757 454
rect 2711 408 2717 442
rect 2751 408 2757 442
rect 2711 370 2757 408
tri 2675 303 2711 339 se
rect 2711 336 2717 370
rect 2751 336 2757 370
rect 2711 303 2757 336
rect 468 251 474 303
rect 526 251 538 303
rect 590 251 2031 303
rect 2083 251 2095 303
rect 2147 291 2757 303
rect 2147 251 2717 291
tri 2717 251 2757 291 nw
rect 2893 442 2939 454
rect 2893 408 2899 442
rect 2933 408 2939 442
rect 2893 370 2939 408
rect 2893 336 2899 370
rect 2933 336 2939 370
tri 2866 211 2893 238 se
rect 2893 211 2939 336
rect 906 205 1941 211
rect 958 159 1941 205
rect 1993 159 2005 211
rect 2057 210 2939 211
rect 2057 159 2888 210
tri 2888 159 2939 210 nw
rect 906 141 958 153
rect 906 83 958 89
rect 1702 -943 1968 -936
rect 1702 -977 1850 -943
rect 1884 -977 1922 -943
rect 1956 -977 1968 -943
rect 1702 -983 1968 -977
rect 2101 -968 2153 -962
tri 1702 -1021 1740 -983 nw
rect 2101 -1032 2153 -1020
rect 2009 -1047 2101 -1041
rect 2009 -1081 2021 -1047
rect 2055 -1081 2093 -1047
rect 2009 -1084 2101 -1081
rect 2009 -1087 2153 -1084
rect 2101 -1090 2153 -1087
rect 2025 -1223 2031 -1220
rect 2009 -1229 2031 -1223
rect 2083 -1229 2095 -1220
rect 2009 -1263 2021 -1229
rect 2083 -1263 2093 -1229
rect 2009 -1269 2031 -1263
rect 2025 -1272 2031 -1269
rect 2083 -1272 2095 -1263
rect 2147 -1272 2153 -1220
<< via1 >>
rect 474 251 526 303
rect 538 251 590 303
rect 2031 251 2083 303
rect 2095 251 2147 303
rect 906 153 958 205
rect 1941 159 1993 211
rect 2005 159 2057 211
rect 906 89 958 141
rect 2101 -1020 2153 -968
rect 2101 -1047 2153 -1032
rect 2101 -1081 2127 -1047
rect 2127 -1081 2153 -1047
rect 2101 -1084 2153 -1081
rect 2031 -1229 2083 -1220
rect 2095 -1229 2147 -1220
rect 2031 -1263 2055 -1229
rect 2055 -1263 2083 -1229
rect 2095 -1263 2127 -1229
rect 2127 -1263 2147 -1229
rect 2031 -1272 2083 -1263
rect 2095 -1272 2147 -1263
<< metal2 >>
rect 544 303 596 468
rect 468 251 474 303
rect 526 251 538 303
rect 590 251 596 303
rect 2025 251 2031 303
rect 2083 251 2095 303
rect 2147 251 2153 303
rect 906 205 958 211
rect 1935 159 1941 211
rect 1993 159 2005 211
rect 2057 205 2063 211
tri 2063 205 2069 211 sw
rect 2057 159 2069 205
rect 906 141 958 153
rect 906 83 958 89
rect 2017 -1220 2069 159
rect 2101 -968 2153 251
rect 2101 -1032 2153 -1020
rect 2101 -1090 2153 -1084
tri 2069 -1220 2112 -1177 sw
rect 2017 -1272 2031 -1220
rect 2083 -1272 2095 -1220
rect 2147 -1272 2153 -1220
use sky130_fd_pr__model__nfet_highvoltage__example_55959141808139  sky130_fd_pr__model__nfet_highvoltage__example_55959141808139_0
timestamp 1676037725
transform 0 1 1770 -1 0 -1002
box -15 0 311 1
use sky130_fd_pr__model__pfet_highvoltage__example_55959141808141  sky130_fd_pr__model__pfet_highvoltage__example_55959141808141_0
timestamp 1676037725
transform -1 0 2968 0 -1 1102
box -15 0 -14 1
use sky130_fd_pr__model__pfet_highvoltage__example_55959141808141  sky130_fd_pr__model__pfet_highvoltage__example_55959141808141_1
timestamp 1676037725
transform 1 0 2672 0 -1 1102
box -15 0 -14 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_0
timestamp 1676037725
transform 0 -1 2647 -1 0 1159
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_0
timestamp 1676037725
transform 0 -1 2941 -1 0 470
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_1
timestamp 1676037725
transform 0 -1 2765 -1 0 470
box 0 0 1 1
<< properties >>
string GDS_END 32781132
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 32776160
<< end >>
