magic
tech sky130A
magscale 1 2
timestamp 1676037725
<< metal2 >>
rect -7432 33185 -987 33506
rect -7432 32929 -7331 33185
rect -7075 32929 -6807 33185
rect -6551 32929 -6253 33185
rect -5997 32929 -5699 33185
rect -5443 32929 -5175 33185
rect -4919 32929 -4561 33185
rect -4305 32929 -4037 33185
rect -3781 32929 -3483 33185
rect -3227 32929 -2929 33185
rect -2673 32929 -2405 33185
rect -2149 32929 -987 33185
rect -7432 32691 -987 32929
rect -7432 32435 -7331 32691
rect -7075 32435 -6807 32691
rect -6551 32435 -6253 32691
rect -5997 32435 -5699 32691
rect -5443 32435 -5175 32691
rect -4919 32435 -4561 32691
rect -4305 32435 -4037 32691
rect -3781 32435 -3483 32691
rect -3227 32435 -2929 32691
rect -2673 32435 -2405 32691
rect -2149 32435 -987 32691
rect -7432 32077 -987 32435
rect -7432 31821 -7331 32077
rect -7075 31821 -6807 32077
rect -6551 31821 -6253 32077
rect -5997 31821 -5699 32077
rect -5443 31821 -5175 32077
rect -4919 31821 -4561 32077
rect -4305 31821 -4037 32077
rect -3781 31821 -3483 32077
rect -3227 31821 -2929 32077
rect -2673 31821 -2405 32077
rect -2149 31821 -987 32077
rect -7432 31583 -987 31821
rect -7432 31327 -7331 31583
rect -7075 31327 -6807 31583
rect -6551 31327 -6253 31583
rect -5997 31327 -5699 31583
rect -5443 31327 -5175 31583
rect -4919 31327 -4561 31583
rect -4305 31327 -4037 31583
rect -3781 31327 -3483 31583
rect -3227 31327 -2929 31583
rect -2673 31327 -2405 31583
rect -2149 31327 -987 31583
rect -7432 31006 -987 31327
tri -987 31006 1513 33506 sw
tri -2023 28004 979 31006 ne
rect 979 30504 1513 31006
tri 1513 30504 2015 31006 sw
rect 979 30183 7787 30504
rect 979 29927 2504 30183
rect 2760 29927 3028 30183
rect 3284 29927 3582 30183
rect 3838 29927 4136 30183
rect 4392 29927 4660 30183
rect 4916 29927 5274 30183
rect 5530 29927 5798 30183
rect 6054 29927 6352 30183
rect 6608 29927 6906 30183
rect 7162 29927 7430 30183
rect 7686 29927 7787 30183
rect 979 29689 7787 29927
rect 979 29433 2504 29689
rect 2760 29433 3028 29689
rect 3284 29433 3582 29689
rect 3838 29433 4136 29689
rect 4392 29433 4660 29689
rect 4916 29433 5274 29689
rect 5530 29433 5798 29689
rect 6054 29433 6352 29689
rect 6608 29433 6906 29689
rect 7162 29433 7430 29689
rect 7686 29433 7787 29689
rect 979 29075 7787 29433
rect 979 28819 2504 29075
rect 2760 28819 3028 29075
rect 3284 28819 3582 29075
rect 3838 28819 4136 29075
rect 4392 28819 4660 29075
rect 4916 28819 5274 29075
rect 5530 28819 5798 29075
rect 6054 28819 6352 29075
rect 6608 28819 6906 29075
rect 7162 28819 7430 29075
rect 7686 28819 7787 29075
rect 979 28581 7787 28819
rect 979 28325 2504 28581
rect 2760 28325 3028 28581
rect 3284 28325 3582 28581
rect 3838 28325 4136 28581
rect 4392 28325 4660 28581
rect 4916 28325 5274 28581
rect 5530 28325 5798 28581
rect 6054 28325 6352 28581
rect 6608 28325 6906 28581
rect 7162 28325 7430 28581
rect 7686 28325 7787 28581
rect 979 28004 7787 28325
rect -7432 27181 -987 27502
rect -7432 26925 -7331 27181
rect -7075 26925 -6807 27181
rect -6551 26925 -6253 27181
rect -5997 26925 -5699 27181
rect -5443 26925 -5175 27181
rect -4919 26925 -4561 27181
rect -4305 26925 -4037 27181
rect -3781 26925 -3483 27181
rect -3227 26925 -2929 27181
rect -2673 26925 -2405 27181
rect -2149 26925 -987 27181
rect -7432 26687 -987 26925
rect -7432 26431 -7331 26687
rect -7075 26431 -6807 26687
rect -6551 26431 -6253 26687
rect -5997 26431 -5699 26687
rect -5443 26431 -5175 26687
rect -4919 26431 -4561 26687
rect -4305 26431 -4037 26687
rect -3781 26431 -3483 26687
rect -3227 26431 -2929 26687
rect -2673 26431 -2405 26687
rect -2149 26431 -987 26687
rect -7432 26073 -987 26431
rect -7432 25817 -7331 26073
rect -7075 25817 -6807 26073
rect -6551 25817 -6253 26073
rect -5997 25817 -5699 26073
rect -5443 25817 -5175 26073
rect -4919 25817 -4561 26073
rect -4305 25817 -4037 26073
rect -3781 25817 -3483 26073
rect -3227 25817 -2929 26073
rect -2673 25817 -2405 26073
rect -2149 25817 -987 26073
rect -7432 25579 -987 25817
rect -7432 25323 -7331 25579
rect -7075 25323 -6807 25579
rect -6551 25323 -6253 25579
rect -5997 25323 -5699 25579
rect -5443 25323 -5175 25579
rect -4919 25323 -4561 25579
rect -4305 25323 -4037 25579
rect -3781 25323 -3483 25579
rect -3227 25323 -2929 25579
rect -2673 25323 -2405 25579
rect -2149 25323 -987 25579
rect -7432 25002 -987 25323
tri -987 25002 1513 27502 sw
tri -2023 22000 979 25002 ne
rect 979 24500 1513 25002
tri 1513 24500 2015 25002 sw
rect 979 24179 7787 24500
rect 979 23923 2504 24179
rect 2760 23923 3028 24179
rect 3284 23923 3582 24179
rect 3838 23923 4136 24179
rect 4392 23923 4660 24179
rect 4916 23923 5274 24179
rect 5530 23923 5798 24179
rect 6054 23923 6352 24179
rect 6608 23923 6906 24179
rect 7162 23923 7430 24179
rect 7686 23923 7787 24179
rect 979 23685 7787 23923
rect 979 23429 2504 23685
rect 2760 23429 3028 23685
rect 3284 23429 3582 23685
rect 3838 23429 4136 23685
rect 4392 23429 4660 23685
rect 4916 23429 5274 23685
rect 5530 23429 5798 23685
rect 6054 23429 6352 23685
rect 6608 23429 6906 23685
rect 7162 23429 7430 23685
rect 7686 23429 7787 23685
rect 979 23071 7787 23429
rect 979 22815 2504 23071
rect 2760 22815 3028 23071
rect 3284 22815 3582 23071
rect 3838 22815 4136 23071
rect 4392 22815 4660 23071
rect 4916 22815 5274 23071
rect 5530 22815 5798 23071
rect 6054 22815 6352 23071
rect 6608 22815 6906 23071
rect 7162 22815 7430 23071
rect 7686 22815 7787 23071
rect 979 22577 7787 22815
rect 979 22321 2504 22577
rect 2760 22321 3028 22577
rect 3284 22321 3582 22577
rect 3838 22321 4136 22577
rect 4392 22321 4660 22577
rect 4916 22321 5274 22577
rect 5530 22321 5798 22577
rect 6054 22321 6352 22577
rect 6608 22321 6906 22577
rect 7162 22321 7430 22577
rect 7686 22321 7787 22577
rect 979 22000 7787 22321
rect 19408 929 37508 1250
rect 19408 673 19552 929
rect 19808 673 20076 929
rect 20332 673 20630 929
rect 20886 673 37508 929
rect 19408 435 37508 673
rect 19408 179 19552 435
rect 19808 179 20076 435
rect 20332 179 20630 435
rect 20886 179 37508 435
rect 19408 -179 37508 179
rect 19408 -435 19552 -179
rect 19808 -435 20076 -179
rect 20332 -435 20630 -179
rect 20886 -435 37508 -179
rect 19408 -673 37508 -435
rect 19408 -929 19552 -673
rect 19808 -929 20076 -673
rect 20332 -929 20630 -673
rect 20886 -929 37508 -673
rect 19408 -1250 37508 -929
tri -2023 -28004 979 -25002 se
rect 979 -25324 7675 -25002
rect 979 -25580 2393 -25324
rect 2649 -25580 2917 -25324
rect 3173 -25580 3471 -25324
rect 3727 -25580 4025 -25324
rect 4281 -25580 4549 -25324
rect 4805 -25580 5163 -25324
rect 5419 -25580 5687 -25324
rect 5943 -25580 6241 -25324
rect 6497 -25580 6795 -25324
rect 7051 -25580 7319 -25324
rect 7575 -25580 7675 -25324
rect 979 -25818 7675 -25580
rect 979 -26074 2393 -25818
rect 2649 -26074 2917 -25818
rect 3173 -26074 3471 -25818
rect 3727 -26074 4025 -25818
rect 4281 -26074 4549 -25818
rect 4805 -26074 5163 -25818
rect 5419 -26074 5687 -25818
rect 5943 -26074 6241 -25818
rect 6497 -26074 6795 -25818
rect 7051 -26074 7319 -25818
rect 7575 -26074 7675 -25818
rect 979 -26432 7675 -26074
rect 979 -26688 2393 -26432
rect 2649 -26688 2917 -26432
rect 3173 -26688 3471 -26432
rect 3727 -26688 4025 -26432
rect 4281 -26688 4549 -26432
rect 4805 -26688 5163 -26432
rect 5419 -26688 5687 -26432
rect 5943 -26688 6241 -26432
rect 6497 -26688 6795 -26432
rect 7051 -26688 7319 -26432
rect 7575 -26688 7675 -26432
rect 979 -26926 7675 -26688
rect 979 -27182 2393 -26926
rect 2649 -27182 2917 -26926
rect 3173 -27182 3471 -26926
rect 3727 -27182 4025 -26926
rect 4281 -27182 4549 -26926
rect 4805 -27182 5163 -26926
rect 5419 -27182 5687 -26926
rect 5943 -27182 6241 -26926
rect 6497 -27182 6795 -26926
rect 7051 -27182 7319 -26926
rect 7575 -27182 7675 -26926
rect 979 -27502 7675 -27182
rect 979 -28004 1513 -27502
tri 1513 -28004 2015 -27502 nw
rect -7544 -28325 -987 -28004
rect -7544 -28581 -7444 -28325
rect -7188 -28581 -6920 -28325
rect -6664 -28581 -6366 -28325
rect -6110 -28581 -5812 -28325
rect -5556 -28581 -5288 -28325
rect -5032 -28581 -4674 -28325
rect -4418 -28581 -4150 -28325
rect -3894 -28581 -3596 -28325
rect -3340 -28581 -3042 -28325
rect -2786 -28581 -2518 -28325
rect -2262 -28581 -987 -28325
rect -7544 -28819 -987 -28581
rect -7544 -29075 -7444 -28819
rect -7188 -29075 -6920 -28819
rect -6664 -29075 -6366 -28819
rect -6110 -29075 -5812 -28819
rect -5556 -29075 -5288 -28819
rect -5032 -29075 -4674 -28819
rect -4418 -29075 -4150 -28819
rect -3894 -29075 -3596 -28819
rect -3340 -29075 -3042 -28819
rect -2786 -29075 -2518 -28819
rect -2262 -29075 -987 -28819
rect -7544 -29433 -987 -29075
rect -7544 -29689 -7444 -29433
rect -7188 -29689 -6920 -29433
rect -6664 -29689 -6366 -29433
rect -6110 -29689 -5812 -29433
rect -5556 -29689 -5288 -29433
rect -5032 -29689 -4674 -29433
rect -4418 -29689 -4150 -29433
rect -3894 -29689 -3596 -29433
rect -3340 -29689 -3042 -29433
rect -2786 -29689 -2518 -29433
rect -2262 -29689 -987 -29433
rect -7544 -29927 -987 -29689
rect -7544 -30183 -7444 -29927
rect -7188 -30183 -6920 -29927
rect -6664 -30183 -6366 -29927
rect -6110 -30183 -5812 -29927
rect -5556 -30183 -5288 -29927
rect -5032 -30183 -4674 -29927
rect -4418 -30183 -4150 -29927
rect -3894 -30183 -3596 -29927
rect -3340 -30183 -3042 -29927
rect -2786 -30183 -2518 -29927
rect -2262 -30183 -987 -29927
rect -7544 -30504 -987 -30183
tri -987 -30504 1513 -28004 nw
tri -2023 -34008 979 -31006 se
rect 979 -31326 7675 -31006
rect 979 -31582 2393 -31326
rect 2649 -31582 2917 -31326
rect 3173 -31582 3471 -31326
rect 3727 -31582 4025 -31326
rect 4281 -31582 4549 -31326
rect 4805 -31582 5163 -31326
rect 5419 -31582 5687 -31326
rect 5943 -31582 6241 -31326
rect 6497 -31582 6795 -31326
rect 7051 -31582 7319 -31326
rect 7575 -31582 7675 -31326
rect 979 -31820 7675 -31582
rect 979 -32076 2393 -31820
rect 2649 -32076 2917 -31820
rect 3173 -32076 3471 -31820
rect 3727 -32076 4025 -31820
rect 4281 -32076 4549 -31820
rect 4805 -32076 5163 -31820
rect 5419 -32076 5687 -31820
rect 5943 -32076 6241 -31820
rect 6497 -32076 6795 -31820
rect 7051 -32076 7319 -31820
rect 7575 -32076 7675 -31820
rect 979 -32434 7675 -32076
rect 979 -32690 2393 -32434
rect 2649 -32690 2917 -32434
rect 3173 -32690 3471 -32434
rect 3727 -32690 4025 -32434
rect 4281 -32690 4549 -32434
rect 4805 -32690 5163 -32434
rect 5419 -32690 5687 -32434
rect 5943 -32690 6241 -32434
rect 6497 -32690 6795 -32434
rect 7051 -32690 7319 -32434
rect 7575 -32690 7675 -32434
rect 979 -32928 7675 -32690
rect 979 -33184 2393 -32928
rect 2649 -33184 2917 -32928
rect 3173 -33184 3471 -32928
rect 3727 -33184 4025 -32928
rect 4281 -33184 4549 -32928
rect 4805 -33184 5163 -32928
rect 5419 -33184 5687 -32928
rect 5943 -33184 6241 -32928
rect 6497 -33184 6795 -32928
rect 7051 -33184 7319 -32928
rect 7575 -33184 7675 -32928
rect 979 -33506 7675 -33184
rect 979 -34008 1513 -33506
tri 1513 -34008 2015 -33506 nw
rect -7544 -34329 -987 -34008
rect -7544 -34585 -7444 -34329
rect -7188 -34585 -6920 -34329
rect -6664 -34585 -6366 -34329
rect -6110 -34585 -5812 -34329
rect -5556 -34585 -5288 -34329
rect -5032 -34585 -4674 -34329
rect -4418 -34585 -4150 -34329
rect -3894 -34585 -3596 -34329
rect -3340 -34585 -3042 -34329
rect -2786 -34585 -2518 -34329
rect -2262 -34585 -987 -34329
rect -7544 -34823 -987 -34585
rect -7544 -35079 -7444 -34823
rect -7188 -35079 -6920 -34823
rect -6664 -35079 -6366 -34823
rect -6110 -35079 -5812 -34823
rect -5556 -35079 -5288 -34823
rect -5032 -35079 -4674 -34823
rect -4418 -35079 -4150 -34823
rect -3894 -35079 -3596 -34823
rect -3340 -35079 -3042 -34823
rect -2786 -35079 -2518 -34823
rect -2262 -35079 -987 -34823
rect -7544 -35437 -987 -35079
rect -7544 -35693 -7444 -35437
rect -7188 -35693 -6920 -35437
rect -6664 -35693 -6366 -35437
rect -6110 -35693 -5812 -35437
rect -5556 -35693 -5288 -35437
rect -5032 -35693 -4674 -35437
rect -4418 -35693 -4150 -35437
rect -3894 -35693 -3596 -35437
rect -3340 -35693 -3042 -35437
rect -2786 -35693 -2518 -35437
rect -2262 -35693 -987 -35437
rect -7544 -35931 -987 -35693
rect -7544 -36187 -7444 -35931
rect -7188 -36187 -6920 -35931
rect -6664 -36187 -6366 -35931
rect -6110 -36187 -5812 -35931
rect -5556 -36187 -5288 -35931
rect -5032 -36187 -4674 -35931
rect -4418 -36187 -4150 -35931
rect -3894 -36187 -3596 -35931
rect -3340 -36187 -3042 -35931
rect -2786 -36187 -2518 -35931
rect -2262 -36187 -987 -35931
rect -7544 -36508 -987 -36187
tri -987 -36508 1513 -34008 nw
<< via2 >>
rect -7331 32929 -7075 33185
rect -6807 32929 -6551 33185
rect -6253 32929 -5997 33185
rect -5699 32929 -5443 33185
rect -5175 32929 -4919 33185
rect -4561 32929 -4305 33185
rect -4037 32929 -3781 33185
rect -3483 32929 -3227 33185
rect -2929 32929 -2673 33185
rect -2405 32929 -2149 33185
rect -7331 32435 -7075 32691
rect -6807 32435 -6551 32691
rect -6253 32435 -5997 32691
rect -5699 32435 -5443 32691
rect -5175 32435 -4919 32691
rect -4561 32435 -4305 32691
rect -4037 32435 -3781 32691
rect -3483 32435 -3227 32691
rect -2929 32435 -2673 32691
rect -2405 32435 -2149 32691
rect -7331 31821 -7075 32077
rect -6807 31821 -6551 32077
rect -6253 31821 -5997 32077
rect -5699 31821 -5443 32077
rect -5175 31821 -4919 32077
rect -4561 31821 -4305 32077
rect -4037 31821 -3781 32077
rect -3483 31821 -3227 32077
rect -2929 31821 -2673 32077
rect -2405 31821 -2149 32077
rect -7331 31327 -7075 31583
rect -6807 31327 -6551 31583
rect -6253 31327 -5997 31583
rect -5699 31327 -5443 31583
rect -5175 31327 -4919 31583
rect -4561 31327 -4305 31583
rect -4037 31327 -3781 31583
rect -3483 31327 -3227 31583
rect -2929 31327 -2673 31583
rect -2405 31327 -2149 31583
rect 2504 29927 2760 30183
rect 3028 29927 3284 30183
rect 3582 29927 3838 30183
rect 4136 29927 4392 30183
rect 4660 29927 4916 30183
rect 5274 29927 5530 30183
rect 5798 29927 6054 30183
rect 6352 29927 6608 30183
rect 6906 29927 7162 30183
rect 7430 29927 7686 30183
rect 2504 29433 2760 29689
rect 3028 29433 3284 29689
rect 3582 29433 3838 29689
rect 4136 29433 4392 29689
rect 4660 29433 4916 29689
rect 5274 29433 5530 29689
rect 5798 29433 6054 29689
rect 6352 29433 6608 29689
rect 6906 29433 7162 29689
rect 7430 29433 7686 29689
rect 2504 28819 2760 29075
rect 3028 28819 3284 29075
rect 3582 28819 3838 29075
rect 4136 28819 4392 29075
rect 4660 28819 4916 29075
rect 5274 28819 5530 29075
rect 5798 28819 6054 29075
rect 6352 28819 6608 29075
rect 6906 28819 7162 29075
rect 7430 28819 7686 29075
rect 2504 28325 2760 28581
rect 3028 28325 3284 28581
rect 3582 28325 3838 28581
rect 4136 28325 4392 28581
rect 4660 28325 4916 28581
rect 5274 28325 5530 28581
rect 5798 28325 6054 28581
rect 6352 28325 6608 28581
rect 6906 28325 7162 28581
rect 7430 28325 7686 28581
rect -7331 26925 -7075 27181
rect -6807 26925 -6551 27181
rect -6253 26925 -5997 27181
rect -5699 26925 -5443 27181
rect -5175 26925 -4919 27181
rect -4561 26925 -4305 27181
rect -4037 26925 -3781 27181
rect -3483 26925 -3227 27181
rect -2929 26925 -2673 27181
rect -2405 26925 -2149 27181
rect -7331 26431 -7075 26687
rect -6807 26431 -6551 26687
rect -6253 26431 -5997 26687
rect -5699 26431 -5443 26687
rect -5175 26431 -4919 26687
rect -4561 26431 -4305 26687
rect -4037 26431 -3781 26687
rect -3483 26431 -3227 26687
rect -2929 26431 -2673 26687
rect -2405 26431 -2149 26687
rect -7331 25817 -7075 26073
rect -6807 25817 -6551 26073
rect -6253 25817 -5997 26073
rect -5699 25817 -5443 26073
rect -5175 25817 -4919 26073
rect -4561 25817 -4305 26073
rect -4037 25817 -3781 26073
rect -3483 25817 -3227 26073
rect -2929 25817 -2673 26073
rect -2405 25817 -2149 26073
rect -7331 25323 -7075 25579
rect -6807 25323 -6551 25579
rect -6253 25323 -5997 25579
rect -5699 25323 -5443 25579
rect -5175 25323 -4919 25579
rect -4561 25323 -4305 25579
rect -4037 25323 -3781 25579
rect -3483 25323 -3227 25579
rect -2929 25323 -2673 25579
rect -2405 25323 -2149 25579
rect 2504 23923 2760 24179
rect 3028 23923 3284 24179
rect 3582 23923 3838 24179
rect 4136 23923 4392 24179
rect 4660 23923 4916 24179
rect 5274 23923 5530 24179
rect 5798 23923 6054 24179
rect 6352 23923 6608 24179
rect 6906 23923 7162 24179
rect 7430 23923 7686 24179
rect 2504 23429 2760 23685
rect 3028 23429 3284 23685
rect 3582 23429 3838 23685
rect 4136 23429 4392 23685
rect 4660 23429 4916 23685
rect 5274 23429 5530 23685
rect 5798 23429 6054 23685
rect 6352 23429 6608 23685
rect 6906 23429 7162 23685
rect 7430 23429 7686 23685
rect 2504 22815 2760 23071
rect 3028 22815 3284 23071
rect 3582 22815 3838 23071
rect 4136 22815 4392 23071
rect 4660 22815 4916 23071
rect 5274 22815 5530 23071
rect 5798 22815 6054 23071
rect 6352 22815 6608 23071
rect 6906 22815 7162 23071
rect 7430 22815 7686 23071
rect 2504 22321 2760 22577
rect 3028 22321 3284 22577
rect 3582 22321 3838 22577
rect 4136 22321 4392 22577
rect 4660 22321 4916 22577
rect 5274 22321 5530 22577
rect 5798 22321 6054 22577
rect 6352 22321 6608 22577
rect 6906 22321 7162 22577
rect 7430 22321 7686 22577
rect 19552 673 19808 929
rect 20076 673 20332 929
rect 20630 673 20886 929
rect 19552 179 19808 435
rect 20076 179 20332 435
rect 20630 179 20886 435
rect 19552 -435 19808 -179
rect 20076 -435 20332 -179
rect 20630 -435 20886 -179
rect 19552 -929 19808 -673
rect 20076 -929 20332 -673
rect 20630 -929 20886 -673
rect 2393 -25580 2649 -25324
rect 2917 -25580 3173 -25324
rect 3471 -25580 3727 -25324
rect 4025 -25580 4281 -25324
rect 4549 -25580 4805 -25324
rect 5163 -25580 5419 -25324
rect 5687 -25580 5943 -25324
rect 6241 -25580 6497 -25324
rect 6795 -25580 7051 -25324
rect 7319 -25580 7575 -25324
rect 2393 -26074 2649 -25818
rect 2917 -26074 3173 -25818
rect 3471 -26074 3727 -25818
rect 4025 -26074 4281 -25818
rect 4549 -26074 4805 -25818
rect 5163 -26074 5419 -25818
rect 5687 -26074 5943 -25818
rect 6241 -26074 6497 -25818
rect 6795 -26074 7051 -25818
rect 7319 -26074 7575 -25818
rect 2393 -26688 2649 -26432
rect 2917 -26688 3173 -26432
rect 3471 -26688 3727 -26432
rect 4025 -26688 4281 -26432
rect 4549 -26688 4805 -26432
rect 5163 -26688 5419 -26432
rect 5687 -26688 5943 -26432
rect 6241 -26688 6497 -26432
rect 6795 -26688 7051 -26432
rect 7319 -26688 7575 -26432
rect 2393 -27182 2649 -26926
rect 2917 -27182 3173 -26926
rect 3471 -27182 3727 -26926
rect 4025 -27182 4281 -26926
rect 4549 -27182 4805 -26926
rect 5163 -27182 5419 -26926
rect 5687 -27182 5943 -26926
rect 6241 -27182 6497 -26926
rect 6795 -27182 7051 -26926
rect 7319 -27182 7575 -26926
rect -7444 -28581 -7188 -28325
rect -6920 -28581 -6664 -28325
rect -6366 -28581 -6110 -28325
rect -5812 -28581 -5556 -28325
rect -5288 -28581 -5032 -28325
rect -4674 -28581 -4418 -28325
rect -4150 -28581 -3894 -28325
rect -3596 -28581 -3340 -28325
rect -3042 -28581 -2786 -28325
rect -2518 -28581 -2262 -28325
rect -7444 -29075 -7188 -28819
rect -6920 -29075 -6664 -28819
rect -6366 -29075 -6110 -28819
rect -5812 -29075 -5556 -28819
rect -5288 -29075 -5032 -28819
rect -4674 -29075 -4418 -28819
rect -4150 -29075 -3894 -28819
rect -3596 -29075 -3340 -28819
rect -3042 -29075 -2786 -28819
rect -2518 -29075 -2262 -28819
rect -7444 -29689 -7188 -29433
rect -6920 -29689 -6664 -29433
rect -6366 -29689 -6110 -29433
rect -5812 -29689 -5556 -29433
rect -5288 -29689 -5032 -29433
rect -4674 -29689 -4418 -29433
rect -4150 -29689 -3894 -29433
rect -3596 -29689 -3340 -29433
rect -3042 -29689 -2786 -29433
rect -2518 -29689 -2262 -29433
rect -7444 -30183 -7188 -29927
rect -6920 -30183 -6664 -29927
rect -6366 -30183 -6110 -29927
rect -5812 -30183 -5556 -29927
rect -5288 -30183 -5032 -29927
rect -4674 -30183 -4418 -29927
rect -4150 -30183 -3894 -29927
rect -3596 -30183 -3340 -29927
rect -3042 -30183 -2786 -29927
rect -2518 -30183 -2262 -29927
rect 2393 -31582 2649 -31326
rect 2917 -31582 3173 -31326
rect 3471 -31582 3727 -31326
rect 4025 -31582 4281 -31326
rect 4549 -31582 4805 -31326
rect 5163 -31582 5419 -31326
rect 5687 -31582 5943 -31326
rect 6241 -31582 6497 -31326
rect 6795 -31582 7051 -31326
rect 7319 -31582 7575 -31326
rect 2393 -32076 2649 -31820
rect 2917 -32076 3173 -31820
rect 3471 -32076 3727 -31820
rect 4025 -32076 4281 -31820
rect 4549 -32076 4805 -31820
rect 5163 -32076 5419 -31820
rect 5687 -32076 5943 -31820
rect 6241 -32076 6497 -31820
rect 6795 -32076 7051 -31820
rect 7319 -32076 7575 -31820
rect 2393 -32690 2649 -32434
rect 2917 -32690 3173 -32434
rect 3471 -32690 3727 -32434
rect 4025 -32690 4281 -32434
rect 4549 -32690 4805 -32434
rect 5163 -32690 5419 -32434
rect 5687 -32690 5943 -32434
rect 6241 -32690 6497 -32434
rect 6795 -32690 7051 -32434
rect 7319 -32690 7575 -32434
rect 2393 -33184 2649 -32928
rect 2917 -33184 3173 -32928
rect 3471 -33184 3727 -32928
rect 4025 -33184 4281 -32928
rect 4549 -33184 4805 -32928
rect 5163 -33184 5419 -32928
rect 5687 -33184 5943 -32928
rect 6241 -33184 6497 -32928
rect 6795 -33184 7051 -32928
rect 7319 -33184 7575 -32928
rect -7444 -34585 -7188 -34329
rect -6920 -34585 -6664 -34329
rect -6366 -34585 -6110 -34329
rect -5812 -34585 -5556 -34329
rect -5288 -34585 -5032 -34329
rect -4674 -34585 -4418 -34329
rect -4150 -34585 -3894 -34329
rect -3596 -34585 -3340 -34329
rect -3042 -34585 -2786 -34329
rect -2518 -34585 -2262 -34329
rect -7444 -35079 -7188 -34823
rect -6920 -35079 -6664 -34823
rect -6366 -35079 -6110 -34823
rect -5812 -35079 -5556 -34823
rect -5288 -35079 -5032 -34823
rect -4674 -35079 -4418 -34823
rect -4150 -35079 -3894 -34823
rect -3596 -35079 -3340 -34823
rect -3042 -35079 -2786 -34823
rect -2518 -35079 -2262 -34823
rect -7444 -35693 -7188 -35437
rect -6920 -35693 -6664 -35437
rect -6366 -35693 -6110 -35437
rect -5812 -35693 -5556 -35437
rect -5288 -35693 -5032 -35437
rect -4674 -35693 -4418 -35437
rect -4150 -35693 -3894 -35437
rect -3596 -35693 -3340 -35437
rect -3042 -35693 -2786 -35437
rect -2518 -35693 -2262 -35437
rect -7444 -36187 -7188 -35931
rect -6920 -36187 -6664 -35931
rect -6366 -36187 -6110 -35931
rect -5812 -36187 -5556 -35931
rect -5288 -36187 -5032 -35931
rect -4674 -36187 -4418 -35931
rect -4150 -36187 -3894 -35931
rect -3596 -36187 -3340 -35931
rect -3042 -36187 -2786 -35931
rect -2518 -36187 -2262 -35931
<< metal3 >>
tri -18660 32972 -15124 36508 se
rect -15124 36340 15124 36508
tri 15124 36340 15292 36508 sw
rect -15124 34008 15292 36340
rect -15124 33506 -14590 34008
tri -14590 33506 -14088 34008 nw
tri 14088 33506 14590 34008 ne
rect 14590 33506 15292 34008
tri -15124 32972 -14590 33506 nw
tri -14415 32972 -13881 33506 se
rect -13881 33286 -2268 33506
tri -2268 33286 -2048 33506 sw
rect -13881 33185 -2048 33286
rect -13881 32972 -7331 33185
tri -22196 29436 -18660 32972 se
rect -18660 32263 -15833 32972
tri -15833 32263 -15124 32972 nw
tri -15124 32263 -14415 32972 se
rect -14415 32929 -7331 32972
rect -7075 32929 -6807 33185
rect -6551 32929 -6253 33185
rect -5997 32929 -5699 33185
rect -5443 32929 -5175 33185
rect -4919 32929 -4561 33185
rect -4305 32929 -4037 33185
rect -3781 32929 -3483 33185
rect -3227 32929 -2929 33185
rect -2673 32929 -2405 33185
rect -2149 32929 -2048 33185
rect -14415 32691 -2048 32929
rect -14415 32435 -7331 32691
rect -7075 32435 -6807 32691
rect -6551 32435 -6253 32691
rect -5997 32435 -5699 32691
rect -5443 32435 -5175 32691
rect -4919 32435 -4561 32691
rect -4305 32435 -4037 32691
rect -3781 32435 -3483 32691
rect -3227 32435 -2929 32691
rect -2673 32435 -2405 32691
rect -2149 32435 -2048 32691
rect -14415 32263 -2048 32435
rect -18660 31554 -16542 32263
tri -16542 31554 -15833 32263 nw
tri -15833 31554 -15124 32263 se
rect -15124 32077 -2048 32263
rect -15124 31821 -7331 32077
rect -7075 31821 -6807 32077
rect -6551 31821 -6253 32077
rect -5997 31821 -5699 32077
rect -5443 31821 -5175 32077
rect -4919 31821 -4561 32077
rect -4305 31821 -4037 32077
rect -3781 31821 -3483 32077
rect -3227 31821 -2929 32077
rect -2673 31821 -2405 32077
rect -2149 31821 -2048 32077
rect -15124 31583 -2048 31821
rect -15124 31554 -7331 31583
rect -18660 31388 -16708 31554
tri -16708 31388 -16542 31554 nw
tri -15999 31388 -15833 31554 se
rect -15833 31388 -7331 31554
rect -18660 30679 -17417 31388
tri -17417 30679 -16708 31388 nw
tri -16708 30679 -15999 31388 se
rect -15999 31327 -7331 31388
rect -7075 31327 -6807 31583
rect -6551 31327 -6253 31583
rect -5997 31327 -5699 31583
rect -5443 31327 -5175 31583
rect -4919 31327 -4561 31583
rect -4305 31327 -4037 31583
rect -3781 31327 -3483 31583
rect -3227 31327 -2929 31583
rect -2673 31327 -2405 31583
rect -2149 31327 -2048 31583
rect -15999 31226 -2048 31327
rect -15999 31006 -2268 31226
tri -2268 31006 -2048 31226 nw
rect -15999 30679 -13347 31006
rect -18660 29970 -18126 30679
tri -18126 29970 -17417 30679 nw
tri -17417 29970 -16708 30679 se
rect -16708 30504 -13347 30679
tri -13347 30504 -12845 31006 nw
tri -2015 30504 987 33506 se
rect 987 32804 13881 33506
tri 13881 32804 14583 33506 sw
tri 14590 32804 15292 33506 ne
tri 15292 32804 18828 36340 sw
rect 987 32095 14583 32804
tri 14583 32095 15292 32804 sw
tri 15292 32095 16001 32804 ne
rect 16001 32095 18828 32804
rect 987 31561 15292 32095
tri 15292 31561 15826 32095 sw
tri 16001 31561 16535 32095 ne
rect 16535 31561 18828 32095
rect 987 31006 15826 31561
rect 987 30504 1301 31006
rect -16708 29970 -13881 30504
tri -13881 29970 -13347 30504 nw
tri -13171 29970 -12637 30504 se
rect -12637 30284 1301 30504
tri 1301 30284 2023 31006 nw
tri 2403 30284 2623 30504 se
rect 2623 30317 12637 30504
tri 12637 30317 12824 30504 sw
tri 12845 30317 13534 31006 ne
rect 13534 30852 15826 31006
tri 15826 30852 16535 31561 sw
tri 16535 30852 17244 31561 ne
rect 17244 30852 18828 31561
rect 13534 30686 16535 30852
tri 16535 30686 16701 30852 sw
tri 17244 30686 17410 30852 ne
rect 17410 30686 18828 30852
rect 13534 30317 16701 30686
rect 2623 30284 12824 30317
rect -12637 29970 -979 30284
tri -18660 29436 -18126 29970 nw
tri -17951 29436 -17417 29970 se
rect -17417 29436 -14591 29970
tri -25732 25900 -22196 29436 se
rect -22196 28727 -19369 29436
tri -19369 28727 -18660 29436 nw
tri -18660 28727 -17951 29436 se
rect -17951 29260 -14591 29436
tri -14591 29260 -13881 29970 nw
tri -13881 29260 -13171 29970 se
rect -13171 29260 -979 29970
rect -17951 28727 -15301 29260
rect -22196 28018 -20078 28727
tri -20078 28018 -19369 28727 nw
tri -19369 28018 -18660 28727 se
rect -18660 28550 -15301 28727
tri -15301 28550 -14591 29260 nw
tri -14591 28550 -13881 29260 se
rect -13881 28550 -979 29260
rect -18660 28388 -15463 28550
tri -15463 28388 -15301 28550 nw
tri -14753 28388 -14591 28550 se
rect -14591 28388 -979 28550
rect -18660 28018 -16173 28388
rect -22196 27852 -20244 28018
tri -20244 27852 -20078 28018 nw
tri -19535 27852 -19369 28018 se
rect -19369 27852 -16173 28018
rect -22196 27143 -20953 27852
tri -20953 27143 -20244 27852 nw
tri -20244 27143 -19535 27852 se
rect -19535 27678 -16173 27852
tri -16173 27678 -15463 28388 nw
tri -15463 27678 -14753 28388 se
rect -14753 28004 -979 28388
tri -979 28004 1301 30284 nw
rect 2403 30183 12824 30284
rect 2403 29927 2504 30183
rect 2760 29927 3028 30183
rect 3284 29927 3582 30183
rect 3838 29927 4136 30183
rect 4392 29927 4660 30183
rect 4916 29927 5274 30183
rect 5530 29927 5798 30183
rect 6054 29927 6352 30183
rect 6608 29927 6906 30183
rect 7162 29927 7430 30183
rect 7686 29970 12824 30183
tri 12824 29970 13171 30317 sw
tri 13534 29970 13881 30317 ne
rect 13881 29977 16701 30317
tri 16701 29977 17410 30686 sw
tri 17410 29977 18119 30686 ne
rect 18119 29977 18828 30686
rect 13881 29970 17410 29977
rect 7686 29927 13171 29970
rect 2403 29689 13171 29927
rect 2403 29433 2504 29689
rect 2760 29433 3028 29689
rect 3284 29433 3582 29689
rect 3838 29433 4136 29689
rect 4392 29433 4660 29689
rect 4916 29433 5274 29689
rect 5530 29433 5798 29689
rect 6054 29433 6352 29689
rect 6608 29433 6906 29689
rect 7162 29433 7430 29689
rect 7686 29433 13171 29689
rect 2403 29260 13171 29433
tri 13171 29260 13881 29970 sw
tri 13881 29260 14591 29970 ne
rect 14591 29268 17410 29970
tri 17410 29268 18119 29977 sw
tri 18119 29268 18828 29977 ne
tri 18828 29268 22364 32804 sw
rect 14591 29260 18119 29268
rect 2403 29075 13881 29260
rect 2403 28819 2504 29075
rect 2760 28819 3028 29075
rect 3284 28819 3582 29075
rect 3838 28819 4136 29075
rect 4392 28819 4660 29075
rect 4916 28819 5274 29075
rect 5530 28819 5798 29075
rect 6054 28819 6352 29075
rect 6608 28819 6906 29075
rect 7162 28819 7430 29075
rect 7686 28819 13881 29075
rect 2403 28735 13881 28819
tri 13881 28735 14406 29260 sw
tri 14591 28735 15116 29260 ne
rect 15116 28735 18119 29260
rect 2403 28581 14406 28735
rect 2403 28325 2504 28581
rect 2760 28325 3028 28581
rect 3284 28325 3582 28581
rect 3838 28325 4136 28581
rect 4392 28325 4660 28581
rect 4916 28325 5274 28581
rect 5530 28325 5798 28581
rect 6054 28325 6352 28581
rect 6608 28325 6906 28581
rect 7162 28325 7430 28581
rect 7686 28325 14406 28581
rect 2403 28224 14406 28325
tri 2403 28004 2623 28224 ne
rect 2623 28025 14406 28224
tri 14406 28025 15116 28735 sw
tri 15116 28025 15826 28735 ne
rect 15826 28559 18119 28735
tri 18119 28559 18828 29268 sw
tri 18828 28559 19537 29268 ne
rect 19537 28559 22364 29268
rect 15826 28025 18828 28559
tri 18828 28025 19362 28559 sw
tri 19537 28025 20071 28559 ne
rect 20071 28025 22364 28559
rect 2623 28004 15116 28025
rect -14753 27678 -12103 28004
rect -19535 27143 -16883 27678
rect -22196 26434 -21662 27143
tri -21662 26434 -20953 27143 nw
tri -20953 26434 -20244 27143 se
rect -20244 26968 -16883 27143
tri -16883 26968 -16173 27678 nw
tri -16173 26968 -15463 27678 se
rect -15463 27502 -12103 27678
tri -12103 27502 -11601 28004 nw
rect -15463 26968 -12637 27502
tri -12637 26968 -12103 27502 nw
tri -11928 26968 -11394 27502 se
rect -11394 27282 -2268 27502
tri -2268 27282 -2048 27502 sw
rect -11394 27181 -2048 27282
rect -11394 26968 -7331 27181
rect -20244 26434 -17417 26968
tri -17417 26434 -16883 26968 nw
tri -16707 26434 -16173 26968 se
rect -16173 26434 -13346 26968
tri -22196 25900 -21662 26434 nw
tri -21487 25900 -20953 26434 se
rect -20953 25900 -18127 26434
tri -29268 22364 -25732 25900 se
rect -25732 25191 -22905 25900
tri -22905 25191 -22196 25900 nw
tri -22196 25191 -21487 25900 se
rect -21487 25724 -18127 25900
tri -18127 25724 -17417 26434 nw
tri -17417 25724 -16707 26434 se
rect -16707 26259 -13346 26434
tri -13346 26259 -12637 26968 nw
tri -12637 26259 -11928 26968 se
rect -11928 26925 -7331 26968
rect -7075 26925 -6807 27181
rect -6551 26925 -6253 27181
rect -5997 26925 -5699 27181
rect -5443 26925 -5175 27181
rect -4919 26925 -4561 27181
rect -4305 26925 -4037 27181
rect -3781 26925 -3483 27181
rect -3227 26925 -2929 27181
rect -2673 26925 -2405 27181
rect -2149 26925 -2048 27181
rect -11928 26687 -2048 26925
rect -11928 26431 -7331 26687
rect -7075 26431 -6807 26687
rect -6551 26431 -6253 26687
rect -5997 26431 -5699 26687
rect -5443 26431 -5175 26687
rect -4919 26431 -4561 26687
rect -4305 26431 -4037 26687
rect -3781 26431 -3483 26687
rect -3227 26431 -2929 26687
rect -2673 26431 -2405 26687
rect -2149 26431 -2048 26687
rect -11928 26259 -2048 26431
rect -16707 25724 -14055 26259
rect -21487 25191 -18837 25724
rect -25732 24482 -23614 25191
tri -23614 24482 -22905 25191 nw
tri -22905 24482 -22196 25191 se
rect -22196 25014 -18837 25191
tri -18837 25014 -18127 25724 nw
tri -18127 25014 -17417 25724 se
rect -17417 25550 -14055 25724
tri -14055 25550 -13346 26259 nw
tri -13346 25550 -12637 26259 se
rect -12637 26073 -2048 26259
rect -12637 25817 -7331 26073
rect -7075 25817 -6807 26073
rect -6551 25817 -6253 26073
rect -5997 25817 -5699 26073
rect -5443 25817 -5175 26073
rect -4919 25817 -4561 26073
rect -4305 25817 -4037 26073
rect -3781 25817 -3483 26073
rect -3227 25817 -2929 26073
rect -2673 25817 -2405 26073
rect -2149 25817 -2048 26073
rect -12637 25579 -2048 25817
rect -12637 25550 -7331 25579
rect -17417 25384 -14221 25550
tri -14221 25384 -14055 25550 nw
tri -13512 25384 -13346 25550 se
rect -13346 25384 -7331 25550
rect -17417 25014 -14930 25384
rect -22196 24852 -18999 25014
tri -18999 24852 -18837 25014 nw
tri -18289 24852 -18127 25014 se
rect -18127 24852 -14930 25014
rect -22196 24482 -19709 24852
rect -25732 24316 -23780 24482
tri -23780 24316 -23614 24482 nw
tri -23071 24316 -22905 24482 se
rect -22905 24316 -19709 24482
rect -25732 23607 -24489 24316
tri -24489 23607 -23780 24316 nw
tri -23780 23607 -23071 24316 se
rect -23071 24142 -19709 24316
tri -19709 24142 -18999 24852 nw
tri -18999 24142 -18289 24852 se
rect -18289 24675 -14930 24852
tri -14930 24675 -14221 25384 nw
tri -14221 24675 -13512 25384 se
rect -13512 25323 -7331 25384
rect -7075 25323 -6807 25579
rect -6551 25323 -6253 25579
rect -5997 25323 -5699 25579
rect -5443 25323 -5175 25579
rect -4919 25323 -4561 25579
rect -4305 25323 -4037 25579
rect -3781 25323 -3483 25579
rect -3227 25323 -2929 25579
rect -2673 25323 -2405 25579
rect -2149 25323 -2048 25579
rect -13512 25222 -2048 25323
rect -13512 25002 -2268 25222
tri -2268 25002 -2048 25222 nw
rect -13512 24675 -10860 25002
rect -18289 24142 -15639 24675
rect -23071 23607 -20419 24142
rect -25732 22898 -25198 23607
tri -25198 22898 -24489 23607 nw
tri -24489 22898 -23780 23607 se
rect -23780 23432 -20419 23607
tri -20419 23432 -19709 24142 nw
tri -19709 23432 -18999 24142 se
rect -18999 23966 -15639 24142
tri -15639 23966 -14930 24675 nw
tri -14930 23966 -14221 24675 se
rect -14221 24500 -10860 24675
tri -10860 24500 -10358 25002 nw
tri -2015 24500 987 27502 se
rect 987 27490 11394 27502
tri 11394 27490 11406 27502 sw
tri 11601 27490 12115 28004 ne
rect 12115 27490 15116 28004
rect 987 26781 11406 27490
tri 11406 26781 12115 27490 sw
tri 12115 26781 12824 27490 ne
rect 12824 27315 15116 27490
tri 15116 27315 15826 28025 sw
tri 15826 27315 16536 28025 ne
rect 16536 27316 19362 28025
tri 19362 27316 20071 28025 sw
tri 20071 27316 20780 28025 ne
rect 20780 27316 22364 28025
rect 16536 27315 20071 27316
rect 12824 26781 15826 27315
tri 15826 26781 16360 27315 sw
tri 16536 26781 17070 27315 ne
rect 17070 27150 20071 27315
tri 20071 27150 20237 27316 sw
tri 20780 27150 20946 27316 ne
rect 20946 27150 22364 27316
rect 17070 26781 20237 27150
rect 987 26072 12115 26781
tri 12115 26072 12824 26781 sw
tri 12824 26072 13533 26781 ne
rect 13533 26072 16360 26781
rect 987 25538 12824 26072
tri 12824 25538 13358 26072 sw
tri 13533 25538 14067 26072 ne
rect 14067 26071 16360 26072
tri 16360 26071 17070 26781 sw
tri 17070 26071 17780 26781 ne
rect 17780 26441 20237 26781
tri 20237 26441 20946 27150 sw
tri 20946 26441 21655 27150 ne
rect 21655 26441 22364 27150
rect 17780 26071 20946 26441
rect 14067 25909 17070 26071
tri 17070 25909 17232 26071 sw
tri 17780 25909 17942 26071 ne
rect 17942 25909 20946 26071
rect 14067 25538 17232 25909
rect 987 25002 13358 25538
rect 987 24500 1521 25002
tri 1521 24500 2023 25002 nw
rect -14221 23966 -11394 24500
tri -11394 23966 -10860 24500 nw
tri -10684 23966 -10150 24500 se
rect -10150 23966 -979 24500
rect -18999 23432 -16173 23966
tri -16173 23432 -15639 23966 nw
tri -15464 23432 -14930 23966 se
rect -14930 23432 -12104 23966
rect -23780 22898 -20953 23432
tri -20953 22898 -20419 23432 nw
tri -20243 22898 -19709 23432 se
rect -19709 22898 -16882 23432
tri -25732 22364 -25198 22898 nw
tri -25023 22364 -24489 22898 se
rect -24489 22364 -21663 22898
tri -32804 18828 -29268 22364 se
rect -29268 21655 -26441 22364
tri -26441 21655 -25732 22364 nw
tri -25732 21655 -25023 22364 se
rect -25023 22188 -21663 22364
tri -21663 22188 -20953 22898 nw
tri -20953 22188 -20243 22898 se
rect -20243 22723 -16882 22898
tri -16882 22723 -16173 23432 nw
tri -16173 22723 -15464 23432 se
rect -15464 23256 -12104 23432
tri -12104 23256 -11394 23966 nw
tri -11394 23256 -10684 23966 se
rect -10684 23256 -979 23966
rect -15464 22723 -12814 23256
rect -20243 22188 -17591 22723
rect -25023 21655 -22373 22188
rect -29268 20946 -27150 21655
tri -27150 20946 -26441 21655 nw
tri -26441 20946 -25732 21655 se
rect -25732 21478 -22373 21655
tri -22373 21478 -21663 22188 nw
tri -21663 21478 -20953 22188 se
rect -20953 22014 -17591 22188
tri -17591 22014 -16882 22723 nw
tri -16882 22014 -16173 22723 se
rect -16173 22546 -12814 22723
tri -12814 22546 -12104 23256 nw
tri -12104 22546 -11394 23256 se
rect -11394 22546 -979 23256
rect -16173 22384 -12976 22546
tri -12976 22384 -12814 22546 nw
tri -12266 22384 -12104 22546 se
rect -12104 22384 -979 22546
rect -16173 22014 -13686 22384
rect -20953 21848 -17757 22014
tri -17757 21848 -17591 22014 nw
tri -17048 21848 -16882 22014 se
rect -16882 21848 -13686 22014
rect -20953 21478 -18466 21848
rect -25732 21316 -22535 21478
tri -22535 21316 -22373 21478 nw
tri -21825 21316 -21663 21478 se
rect -21663 21316 -18466 21478
rect -25732 20946 -23245 21316
rect -29268 20780 -27316 20946
tri -27316 20780 -27150 20946 nw
tri -26607 20780 -26441 20946 se
rect -26441 20780 -23245 20946
rect -29268 20071 -28025 20780
tri -28025 20071 -27316 20780 nw
tri -27316 20071 -26607 20780 se
rect -26607 20606 -23245 20780
tri -23245 20606 -22535 21316 nw
tri -22535 20606 -21825 21316 se
rect -21825 21139 -18466 21316
tri -18466 21139 -17757 21848 nw
tri -17757 21139 -17048 21848 se
rect -17048 21674 -13686 21848
tri -13686 21674 -12976 22384 nw
tri -12976 21674 -12266 22384 se
rect -12266 22000 -979 22384
tri -979 22000 1521 24500 nw
tri 2403 24280 2623 24500 se
rect 2623 24294 10150 24500
tri 10150 24294 10356 24500 sw
tri 10358 24294 11066 25002 ne
rect 11066 24829 13358 25002
tri 13358 24829 14067 25538 sw
tri 14067 24829 14776 25538 ne
rect 14776 25199 17232 25538
tri 17232 25199 17942 25909 sw
tri 17942 25199 18652 25909 ne
rect 18652 25732 20946 25909
tri 20946 25732 21655 26441 sw
tri 21655 25732 22364 26441 ne
tri 22364 25732 25900 29268 sw
rect 18652 25199 21655 25732
rect 14776 24829 17942 25199
rect 11066 24663 14067 24829
tri 14067 24663 14233 24829 sw
tri 14776 24663 14942 24829 ne
rect 14942 24663 17942 24829
rect 11066 24294 14233 24663
rect 2623 24280 10356 24294
rect 2403 24179 10356 24280
rect 2403 23923 2504 24179
rect 2760 23923 3028 24179
rect 3284 23923 3582 24179
rect 3838 23923 4136 24179
rect 4392 23923 4660 24179
rect 4916 23923 5274 24179
rect 5530 23923 5798 24179
rect 6054 23923 6352 24179
rect 6608 23923 6906 24179
rect 7162 23923 7430 24179
rect 7686 23966 10356 24179
tri 10356 23966 10684 24294 sw
tri 11066 23966 11394 24294 ne
rect 11394 23966 14233 24294
rect 7686 23923 10684 23966
rect 2403 23685 10684 23923
rect 2403 23429 2504 23685
rect 2760 23429 3028 23685
rect 3284 23429 3582 23685
rect 3838 23429 4136 23685
rect 4392 23429 4660 23685
rect 4916 23429 5274 23685
rect 5530 23429 5798 23685
rect 6054 23429 6352 23685
rect 6608 23429 6906 23685
rect 7162 23429 7430 23685
rect 7686 23429 10684 23685
rect 2403 23256 10684 23429
tri 10684 23256 11394 23966 sw
tri 11394 23256 12104 23966 ne
rect 12104 23954 14233 23966
tri 14233 23954 14942 24663 sw
tri 14942 23954 15651 24663 ne
rect 15651 24489 17942 24663
tri 17942 24489 18652 25199 sw
tri 18652 24489 19362 25199 ne
rect 19362 25023 21655 25199
tri 21655 25023 22364 25732 sw
tri 22364 25023 23073 25732 ne
rect 23073 25023 25900 25732
rect 19362 24489 22364 25023
tri 22364 24489 22898 25023 sw
tri 23073 24489 23607 25023 ne
rect 23607 24489 25900 25023
rect 15651 23954 18652 24489
rect 12104 23256 14942 23954
rect 2403 23071 11394 23256
rect 2403 22815 2504 23071
rect 2760 22815 3028 23071
rect 3284 22815 3582 23071
rect 3838 22815 4136 23071
rect 4392 22815 4660 23071
rect 4916 22815 5274 23071
rect 5530 22815 5798 23071
rect 6054 22815 6352 23071
rect 6608 22815 6906 23071
rect 7162 22815 7430 23071
rect 7686 22815 11394 23071
rect 2403 22712 11394 22815
tri 11394 22712 11938 23256 sw
tri 12104 22712 12648 23256 ne
rect 12648 23245 14942 23256
tri 14942 23245 15651 23954 sw
tri 15651 23245 16360 23954 ne
rect 16360 23779 18652 23954
tri 18652 23779 19362 24489 sw
tri 19362 23779 20072 24489 ne
rect 20072 23780 22898 24489
tri 22898 23780 23607 24489 sw
tri 23607 23780 24316 24489 ne
rect 24316 23780 25900 24489
rect 20072 23779 23607 23780
rect 16360 23245 19362 23779
tri 19362 23245 19896 23779 sw
tri 20072 23245 20606 23779 ne
rect 20606 23614 23607 23779
tri 23607 23614 23773 23780 sw
tri 24316 23614 24482 23780 ne
rect 24482 23614 25900 23780
rect 20606 23245 23773 23614
rect 12648 22712 15651 23245
rect 2403 22577 11938 22712
rect 2403 22321 2504 22577
rect 2760 22321 3028 22577
rect 3284 22321 3582 22577
rect 3838 22321 4136 22577
rect 4392 22321 4660 22577
rect 4916 22321 5274 22577
rect 5530 22321 5798 22577
rect 6054 22321 6352 22577
rect 6608 22321 6906 22577
rect 7162 22321 7430 22577
rect 7686 22321 11938 22577
rect 2403 22220 11938 22321
tri 2403 22000 2623 22220 ne
rect 2623 22002 11938 22220
tri 11938 22002 12648 22712 sw
tri 12648 22002 13358 22712 ne
rect 13358 22536 15651 22712
tri 15651 22536 16360 23245 sw
tri 16360 22536 17069 23245 ne
rect 17069 22536 19896 23245
rect 13358 22002 16360 22536
tri 16360 22002 16894 22536 sw
tri 17069 22002 17603 22536 ne
rect 17603 22535 19896 22536
tri 19896 22535 20606 23245 sw
tri 20606 22535 21316 23245 ne
rect 21316 22905 23773 23245
tri 23773 22905 24482 23614 sw
tri 24482 22905 25191 23614 ne
rect 25191 22905 25900 23614
rect 21316 22535 24482 22905
rect 17603 22373 20606 22535
tri 20606 22373 20768 22535 sw
tri 21316 22373 21478 22535 ne
rect 21478 22373 24482 22535
rect 17603 22002 20768 22373
rect 2623 22000 12648 22002
rect -12266 21674 -10150 22000
rect -17048 21139 -14396 21674
rect -21825 20606 -19175 21139
rect -26607 20071 -23955 20606
rect -29268 19362 -28734 20071
tri -28734 19362 -28025 20071 nw
tri -28025 19362 -27316 20071 se
rect -27316 19896 -23955 20071
tri -23955 19896 -23245 20606 nw
tri -23245 19896 -22535 20606 se
rect -22535 20430 -19175 20606
tri -19175 20430 -18466 21139 nw
tri -18466 20430 -17757 21139 se
rect -17757 20964 -14396 21139
tri -14396 20964 -13686 21674 nw
tri -13686 20964 -12976 21674 se
rect -12976 20964 -10150 21674
tri -10150 20964 -9114 22000 nw
rect -17757 20430 -14930 20964
tri -14930 20430 -14396 20964 nw
tri -14220 20430 -13686 20964 se
rect -13686 20430 -10684 20964
tri -10684 20430 -10150 20964 nw
tri 9114 20758 10356 22000 ne
rect 10356 21292 12648 22000
tri 12648 21292 13358 22002 sw
tri 13358 21292 14068 22002 ne
rect 14068 21293 16894 22002
tri 16894 21293 17603 22002 sw
tri 17603 21293 18312 22002 ne
rect 18312 21663 20768 22002
tri 20768 21663 21478 22373 sw
tri 21478 21663 22188 22373 ne
rect 22188 22196 24482 22373
tri 24482 22196 25191 22905 sw
tri 25191 22196 25900 22905 ne
tri 25900 22196 29436 25732 sw
rect 22188 21663 25191 22196
rect 18312 21293 21478 21663
rect 14068 21292 17603 21293
rect 10356 20758 13358 21292
tri 13358 20758 13892 21292 sw
tri 14068 20758 14602 21292 ne
rect 14602 21127 17603 21292
tri 17603 21127 17769 21293 sw
tri 18312 21127 18478 21293 ne
rect 18478 21127 21478 21293
rect 14602 20758 17769 21127
rect -22535 19896 -19709 20430
tri -19709 19896 -19175 20430 nw
tri -19000 19896 -18466 20430 se
rect -18466 19896 -15640 20430
rect -27316 19362 -24489 19896
tri -24489 19362 -23955 19896 nw
tri -23779 19362 -23245 19896 se
rect -23245 19362 -20418 19896
tri -29268 18828 -28734 19362 nw
tri -28559 18828 -28025 19362 se
rect -28025 18828 -25199 19362
tri -36340 15292 -32804 18828 se
rect -32804 18119 -29977 18828
tri -29977 18119 -29268 18828 nw
tri -29268 18119 -28559 18828 se
rect -28559 18652 -25199 18828
tri -25199 18652 -24489 19362 nw
tri -24489 18652 -23779 19362 se
rect -23779 19187 -20418 19362
tri -20418 19187 -19709 19896 nw
tri -19709 19187 -19000 19896 se
rect -19000 19720 -15640 19896
tri -15640 19720 -14930 20430 nw
tri -14930 19720 -14220 20430 se
rect -14220 19720 -13686 20430
rect -19000 19187 -16350 19720
rect -23779 18652 -21127 19187
rect -28559 18119 -25909 18652
rect -32804 17410 -30686 18119
tri -30686 17410 -29977 18119 nw
tri -29977 17410 -29268 18119 se
rect -29268 17942 -25909 18119
tri -25909 17942 -25199 18652 nw
tri -25199 17942 -24489 18652 se
rect -24489 18478 -21127 18652
tri -21127 18478 -20418 19187 nw
tri -20418 18478 -19709 19187 se
rect -19709 19010 -16350 19187
tri -16350 19010 -15640 19720 nw
tri -15640 19010 -14930 19720 se
rect -14930 19010 -13686 19720
rect -19709 18848 -16512 19010
tri -16512 18848 -16350 19010 nw
tri -15802 18848 -15640 19010 se
rect -15640 18848 -13686 19010
rect -19709 18478 -17222 18848
rect -24489 18312 -21293 18478
tri -21293 18312 -21127 18478 nw
tri -20584 18312 -20418 18478 se
rect -20418 18312 -17222 18478
rect -24489 17942 -22002 18312
rect -29268 17780 -26071 17942
tri -26071 17780 -25909 17942 nw
tri -25361 17780 -25199 17942 se
rect -25199 17780 -22002 17942
rect -29268 17410 -26781 17780
rect -32804 17244 -30852 17410
tri -30852 17244 -30686 17410 nw
tri -30143 17244 -29977 17410 se
rect -29977 17244 -26781 17410
rect -32804 16535 -31561 17244
tri -31561 16535 -30852 17244 nw
tri -30852 16535 -30143 17244 se
rect -30143 17070 -26781 17244
tri -26781 17070 -26071 17780 nw
tri -26071 17070 -25361 17780 se
rect -25361 17603 -22002 17780
tri -22002 17603 -21293 18312 nw
tri -21293 17603 -20584 18312 se
rect -20584 18138 -17222 18312
tri -17222 18138 -16512 18848 nw
tri -16512 18138 -15802 18848 se
rect -15802 18138 -13686 18848
rect -20584 17603 -17932 18138
rect -25361 17070 -22711 17603
rect -30143 16535 -27491 17070
rect -32804 15826 -32270 16535
tri -32270 15826 -31561 16535 nw
tri -31561 15826 -30852 16535 se
rect -30852 16360 -27491 16535
tri -27491 16360 -26781 17070 nw
tri -26781 16360 -26071 17070 se
rect -26071 16894 -22711 17070
tri -22711 16894 -22002 17603 nw
tri -22002 16894 -21293 17603 se
rect -21293 17428 -17932 17603
tri -17932 17428 -17222 18138 nw
tri -17222 17428 -16512 18138 se
rect -16512 17428 -13686 18138
tri -13686 17428 -10684 20430 nw
tri 10356 18466 12648 20758 ne
rect 12648 20048 13892 20758
tri 13892 20048 14602 20758 sw
tri 14602 20048 15312 20758 ne
rect 15312 20418 17769 20758
tri 17769 20418 18478 21127 sw
tri 18478 20418 19187 21127 ne
rect 19187 20953 21478 21127
tri 21478 20953 22188 21663 sw
tri 22188 20953 22898 21663 ne
rect 22898 21487 25191 21663
tri 25191 21487 25900 22196 sw
tri 25900 21487 26609 22196 ne
rect 26609 21487 29436 22196
rect 22898 20953 25900 21487
tri 25900 20953 26434 21487 sw
tri 26609 20953 27143 21487 ne
rect 27143 20953 29436 21487
rect 19187 20418 22188 20953
rect 15312 20048 18478 20418
rect 12648 19886 14602 20048
tri 14602 19886 14764 20048 sw
tri 15312 19886 15474 20048 ne
rect 15474 19886 18478 20048
rect 12648 19176 14764 19886
tri 14764 19176 15474 19886 sw
tri 15474 19176 16184 19886 ne
rect 16184 19709 18478 19886
tri 18478 19709 19187 20418 sw
tri 19187 19709 19896 20418 ne
rect 19896 20243 22188 20418
tri 22188 20243 22898 20953 sw
tri 22898 20243 23608 20953 ne
rect 23608 20244 26434 20953
tri 26434 20244 27143 20953 sw
tri 27143 20244 27852 20953 ne
rect 27852 20244 29436 20953
rect 23608 20243 27143 20244
rect 19896 19709 22898 20243
tri 22898 19709 23432 20243 sw
tri 23608 19709 24142 20243 ne
rect 24142 20078 27143 20243
tri 27143 20078 27309 20244 sw
tri 27852 20078 28018 20244 ne
rect 28018 20078 29436 20244
rect 24142 19709 27309 20078
rect 16184 19176 19187 19709
rect 12648 18466 15474 19176
tri 15474 18466 16184 19176 sw
tri 16184 18466 16894 19176 ne
rect 16894 19000 19187 19176
tri 19187 19000 19896 19709 sw
tri 19896 19000 20605 19709 ne
rect 20605 19000 23432 19709
rect 16894 18466 19896 19000
tri 19896 18466 20430 19000 sw
tri 20605 18466 21139 19000 ne
rect 21139 18999 23432 19000
tri 23432 18999 24142 19709 sw
tri 24142 18999 24852 19709 ne
rect 24852 19369 27309 19709
tri 27309 19369 28018 20078 sw
tri 28018 19369 28727 20078 ne
rect 28727 19369 29436 20078
rect 24852 18999 28018 19369
rect 21139 18837 24142 18999
tri 24142 18837 24304 18999 sw
tri 24852 18837 25014 18999 ne
rect 25014 18837 28018 18999
rect 21139 18466 24304 18837
rect -21293 16894 -18466 17428
tri -18466 16894 -17932 17428 nw
tri -17756 16894 -17222 17428 se
rect -17222 16894 -14220 17428
tri -14220 16894 -13686 17428 nw
tri 12648 17222 13892 18466 ne
rect 13892 17756 16184 18466
tri 16184 17756 16894 18466 sw
tri 16894 17756 17604 18466 ne
rect 17604 17757 20430 18466
tri 20430 17757 21139 18466 sw
tri 21139 17757 21848 18466 ne
rect 21848 18127 24304 18466
tri 24304 18127 25014 18837 sw
tri 25014 18127 25724 18837 ne
rect 25724 18660 28018 18837
tri 28018 18660 28727 19369 sw
tri 28727 18660 29436 19369 ne
tri 29436 18660 32972 22196 sw
rect 25724 18127 28727 18660
rect 21848 17757 25014 18127
rect 17604 17756 21139 17757
rect 13892 17222 16894 17756
tri 16894 17222 17428 17756 sw
tri 17604 17222 18138 17756 ne
rect 18138 17591 21139 17756
tri 21139 17591 21305 17757 sw
tri 21848 17591 22014 17757 ne
rect 22014 17591 25014 17757
rect 18138 17222 21305 17591
rect -26071 16360 -23245 16894
tri -23245 16360 -22711 16894 nw
tri -22536 16360 -22002 16894 se
rect -22002 16360 -19176 16894
rect -30852 15826 -28025 16360
tri -28025 15826 -27491 16360 nw
tri -27315 15826 -26781 16360 se
rect -26781 15826 -23954 16360
tri -32804 15292 -32270 15826 nw
tri -32095 15292 -31561 15826 se
rect -31561 15292 -28735 15826
tri -36508 15124 -36340 15292 se
rect -36340 15124 -32972 15292
tri -32972 15124 -32804 15292 nw
tri -32263 15124 -32095 15292 se
rect -32095 15124 -28735 15292
rect -36508 14415 -33681 15124
tri -33681 14415 -32972 15124 nw
tri -32972 14415 -32263 15124 se
rect -32263 15116 -28735 15124
tri -28735 15116 -28025 15826 nw
tri -28025 15116 -27315 15826 se
rect -27315 15651 -23954 15826
tri -23954 15651 -23245 16360 nw
tri -23245 15651 -22536 16360 se
rect -22536 16184 -19176 16360
tri -19176 16184 -18466 16894 nw
tri -18466 16184 -17756 16894 se
rect -17756 16184 -17222 16894
rect -22536 15651 -19886 16184
rect -27315 15116 -24663 15651
rect -32263 14591 -29260 15116
tri -29260 14591 -28735 15116 nw
tri -28550 14591 -28025 15116 se
rect -28025 14942 -24663 15116
tri -24663 14942 -23954 15651 nw
tri -23954 14942 -23245 15651 se
rect -23245 15474 -19886 15651
tri -19886 15474 -19176 16184 nw
tri -19176 15474 -18466 16184 se
rect -18466 15474 -17222 16184
rect -23245 15312 -20048 15474
tri -20048 15312 -19886 15474 nw
tri -19338 15312 -19176 15474 se
rect -19176 15312 -17222 15474
rect -23245 14942 -20758 15312
rect -28025 14776 -24829 14942
tri -24829 14776 -24663 14942 nw
tri -24120 14776 -23954 14942 se
rect -23954 14776 -20758 14942
rect -28025 14591 -25538 14776
rect -32263 14415 -29970 14591
rect -36508 -14415 -34008 14415
tri -34008 14088 -33681 14415 nw
tri -33506 13881 -32972 14415 se
rect -32972 13881 -29970 14415
tri -29970 13881 -29260 14591 nw
tri -29260 13881 -28550 14591 se
rect -28550 14067 -25538 14591
tri -25538 14067 -24829 14776 nw
tri -24829 14067 -24120 14776 se
rect -24120 14602 -20758 14776
tri -20758 14602 -20048 15312 nw
tri -20048 14602 -19338 15312 se
rect -19338 14602 -17222 15312
rect -24120 14067 -21468 14602
rect -28550 13881 -26247 14067
rect -33506 13171 -30680 13881
tri -30680 13171 -29970 13881 nw
tri -29970 13171 -29260 13881 se
rect -29260 13358 -26247 13881
tri -26247 13358 -25538 14067 nw
tri -25538 13358 -24829 14067 se
rect -24829 13892 -21468 14067
tri -21468 13892 -20758 14602 nw
tri -20758 13892 -20048 14602 se
rect -20048 13892 -17222 14602
tri -17222 13892 -14220 16894 nw
tri 13892 14930 16184 17222 ne
rect 16184 16512 17428 17222
tri 17428 16512 18138 17222 sw
tri 18138 16512 18848 17222 ne
rect 18848 16882 21305 17222
tri 21305 16882 22014 17591 sw
tri 22014 16882 22723 17591 ne
rect 22723 17417 25014 17591
tri 25014 17417 25724 18127 sw
tri 25724 17417 26434 18127 ne
rect 26434 17951 28727 18127
tri 28727 17951 29436 18660 sw
tri 29436 17951 30145 18660 ne
rect 30145 17951 32972 18660
rect 26434 17417 29436 17951
tri 29436 17417 29970 17951 sw
tri 30145 17417 30679 17951 ne
rect 30679 17417 32972 17951
rect 22723 16882 25724 17417
rect 18848 16512 22014 16882
rect 16184 16350 18138 16512
tri 18138 16350 18300 16512 sw
tri 18848 16350 19010 16512 ne
rect 19010 16350 22014 16512
rect 16184 15640 18300 16350
tri 18300 15640 19010 16350 sw
tri 19010 15640 19720 16350 ne
rect 19720 16173 22014 16350
tri 22014 16173 22723 16882 sw
tri 22723 16173 23432 16882 ne
rect 23432 16707 25724 16882
tri 25724 16707 26434 17417 sw
tri 26434 16707 27144 17417 ne
rect 27144 16708 29970 17417
tri 29970 16708 30679 17417 sw
tri 30679 16708 31388 17417 ne
rect 31388 16708 32972 17417
rect 27144 16707 30679 16708
rect 23432 16173 26434 16707
tri 26434 16173 26968 16707 sw
tri 27144 16173 27678 16707 ne
rect 27678 16542 30679 16707
tri 30679 16542 30845 16708 sw
tri 31388 16542 31554 16708 ne
rect 31554 16542 32972 16708
rect 27678 16173 30845 16542
rect 19720 15640 22723 16173
rect 16184 14930 19010 15640
tri 19010 14930 19720 15640 sw
tri 19720 14930 20430 15640 ne
rect 20430 15464 22723 15640
tri 22723 15464 23432 16173 sw
tri 23432 15464 24141 16173 ne
rect 24141 15464 26968 16173
rect 20430 14930 23432 15464
tri 23432 14930 23966 15464 sw
tri 24141 14930 24675 15464 ne
rect 24675 15463 26968 15464
tri 26968 15463 27678 16173 sw
tri 27678 15463 28388 16173 ne
rect 28388 15833 30845 16173
tri 30845 15833 31554 16542 sw
tri 31554 15833 32263 16542 ne
rect 32263 15833 32972 16542
rect 28388 15463 31554 15833
rect 24675 15301 27678 15463
tri 27678 15301 27840 15463 sw
tri 28388 15301 28550 15463 ne
rect 28550 15301 31554 15463
rect 24675 14930 27840 15301
rect -24829 13358 -22002 13892
tri -22002 13358 -21468 13892 nw
tri -21292 13358 -20758 13892 se
rect -20758 13358 -17756 13892
tri -17756 13358 -17222 13892 nw
tri 16184 13686 17428 14930 ne
rect 17428 14220 19720 14930
tri 19720 14220 20430 14930 sw
tri 20430 14220 21140 14930 ne
rect 21140 14221 23966 14930
tri 23966 14221 24675 14930 sw
tri 24675 14221 25384 14930 ne
rect 25384 14591 27840 14930
tri 27840 14591 28550 15301 sw
tri 28550 14591 29260 15301 ne
rect 29260 15124 31554 15301
tri 31554 15124 32263 15833 sw
tri 32263 15124 32972 15833 ne
tri 32972 15124 36508 18660 sw
rect 29260 14591 32263 15124
rect 25384 14221 28550 14591
rect 21140 14220 24675 14221
rect 17428 13686 20430 14220
tri 20430 13686 20964 14220 sw
tri 21140 13686 21674 14220 ne
rect 21674 14055 24675 14220
tri 24675 14055 24841 14221 sw
tri 25384 14055 25550 14221 ne
rect 25550 14055 28550 14221
rect 21674 13686 24841 14055
rect -29260 13171 -26781 13358
rect -33506 -13171 -31006 13171
tri -31006 12845 -30680 13171 nw
tri -30504 12637 -29970 13171 se
rect -29970 12824 -26781 13171
tri -26781 12824 -26247 13358 nw
tri -26072 12824 -25538 13358 se
rect -25538 12824 -22712 13358
rect -29970 12637 -26968 12824
tri -26968 12637 -26781 12824 nw
tri -26259 12637 -26072 12824 se
rect -26072 12648 -22712 12824
tri -22712 12648 -22002 13358 nw
tri -22002 12648 -21292 13358 se
rect -21292 12648 -20758 13358
rect -26072 12637 -23256 12648
rect -30504 11928 -27677 12637
tri -27677 11928 -26968 12637 nw
tri -26968 11928 -26259 12637 se
rect -26259 12104 -23256 12637
tri -23256 12104 -22712 12648 nw
tri -22546 12104 -22002 12648 se
rect -22002 12104 -20758 12648
rect -26259 11928 -23966 12104
rect -30504 -11928 -28004 11928
tri -28004 11601 -27677 11928 nw
tri -27502 11394 -26968 11928 se
rect -26968 11394 -23966 11928
tri -23966 11394 -23256 12104 nw
tri -23256 11394 -22546 12104 se
rect -22546 11394 -20758 12104
rect -27502 10684 -24676 11394
tri -24676 10684 -23966 11394 nw
tri -23966 10684 -23256 11394 se
rect -23256 10684 -20758 11394
rect -27502 -10684 -25002 10684
tri -25002 10358 -24676 10684 nw
tri -24500 10150 -23966 10684 se
rect -23966 10356 -20758 10684
tri -20758 10356 -17756 13358 nw
tri 17428 11394 19720 13686 ne
rect 19720 12976 20964 13686
tri 20964 12976 21674 13686 sw
tri 21674 12976 22384 13686 ne
rect 22384 13346 24841 13686
tri 24841 13346 25550 14055 sw
tri 25550 13346 26259 14055 ne
rect 26259 13881 28550 14055
tri 28550 13881 29260 14591 sw
tri 29260 13881 29970 14591 ne
rect 29970 14415 32263 14591
tri 32263 14415 32972 15124 sw
tri 32972 14415 33681 15124 ne
rect 33681 14415 36508 15124
rect 29970 13881 32972 14415
tri 32972 13881 33506 14415 sw
tri 33681 14088 34008 14415 ne
rect 26259 13346 29260 13881
rect 22384 12976 25550 13346
rect 19720 12814 21674 12976
tri 21674 12814 21836 12976 sw
tri 22384 12814 22546 12976 ne
rect 22546 12814 25550 12976
rect 19720 12104 21836 12814
tri 21836 12104 22546 12814 sw
tri 22546 12104 23256 12814 ne
rect 23256 12637 25550 12814
tri 25550 12637 26259 13346 sw
tri 26259 12637 26968 13346 ne
rect 26968 13171 29260 13346
tri 29260 13171 29970 13881 sw
tri 29970 13171 30680 13881 ne
rect 30680 13171 33506 13881
rect 26968 12637 29970 13171
tri 29970 12637 30504 13171 sw
tri 30680 12845 31006 13171 ne
rect 23256 12104 26259 12637
rect 19720 11394 22546 12104
tri 22546 11394 23256 12104 sw
tri 23256 11394 23966 12104 ne
rect 23966 11928 26259 12104
tri 26259 11928 26968 12637 sw
tri 26968 11928 27677 12637 ne
rect 27677 11928 30504 12637
rect 23966 11394 26968 11928
tri 26968 11394 27502 11928 sw
tri 27677 11601 28004 11928 ne
rect -23966 10150 -22000 10356
rect -24500 1250 -22000 10150
tri -22000 9114 -20758 10356 nw
tri 19720 9114 22000 11394 ne
rect 22000 10684 23256 11394
tri 23256 10684 23966 11394 sw
tri 23966 10684 24676 11394 ne
rect 24676 10684 27502 11394
rect 22000 10150 23966 10684
tri 23966 10150 24500 10684 sw
tri 24676 10358 25002 10684 ne
rect -24500 929 21000 1250
rect -24500 673 19552 929
rect 19808 673 20076 929
rect 20332 673 20630 929
rect 20886 673 21000 929
rect -24500 435 21000 673
rect -24500 179 19552 435
rect 19808 179 20076 435
rect 20332 179 20630 435
rect 20886 179 21000 435
rect -24500 -179 21000 179
rect -24500 -435 19552 -179
rect 19808 -435 20076 -179
rect 20332 -435 20630 -179
rect 20886 -435 21000 -179
rect -24500 -673 21000 -435
rect -24500 -929 19552 -673
rect 19808 -929 20076 -673
rect 20332 -929 20630 -673
rect 20886 -929 21000 -673
rect -24500 -1250 21000 -929
rect -24500 -10150 -22000 -1250
tri -22000 -10150 -20964 -9114 sw
tri -25002 -10684 -24676 -10358 sw
tri -24500 -10684 -23966 -10150 ne
rect -23966 -10684 -20964 -10150
rect -27502 -11394 -24676 -10684
tri -24676 -11394 -23966 -10684 sw
tri -23966 -11394 -23256 -10684 ne
rect -23256 -11394 -20964 -10684
tri -28004 -11928 -27677 -11601 sw
tri -27502 -11928 -26968 -11394 ne
rect -26968 -11928 -23966 -11394
rect -30504 -12637 -27677 -11928
tri -27677 -12637 -26968 -11928 sw
tri -26968 -12637 -26259 -11928 ne
rect -26259 -12104 -23966 -11928
tri -23966 -12104 -23256 -11394 sw
tri -23256 -12104 -22546 -11394 ne
rect -22546 -12104 -20964 -11394
rect -26259 -12637 -23256 -12104
tri -31006 -13171 -30680 -12845 sw
tri -30504 -13171 -29970 -12637 ne
rect -29970 -13171 -26968 -12637
rect -33506 -13881 -30680 -13171
tri -30680 -13881 -29970 -13171 sw
tri -29970 -13881 -29260 -13171 ne
rect -29260 -13346 -26968 -13171
tri -26968 -13346 -26259 -12637 sw
tri -26259 -13346 -25550 -12637 ne
rect -25550 -12814 -23256 -12637
tri -23256 -12814 -22546 -12104 sw
tri -22546 -12814 -21836 -12104 ne
rect -21836 -12814 -20964 -12104
rect -25550 -12976 -22546 -12814
tri -22546 -12976 -22384 -12814 sw
tri -21836 -12976 -21674 -12814 ne
rect -21674 -12976 -20964 -12814
rect -25550 -13346 -22384 -12976
rect -29260 -13881 -26259 -13346
tri -34008 -14415 -33681 -14088 sw
tri -33506 -14415 -32972 -13881 ne
rect -32972 -14415 -29970 -13881
rect -36508 -15124 -33681 -14415
tri -33681 -15124 -32972 -14415 sw
tri -32972 -15124 -32263 -14415 ne
rect -32263 -14591 -29970 -14415
tri -29970 -14591 -29260 -13881 sw
tri -29260 -14591 -28550 -13881 ne
rect -28550 -14055 -26259 -13881
tri -26259 -14055 -25550 -13346 sw
tri -25550 -14055 -24841 -13346 ne
rect -24841 -13686 -22384 -13346
tri -22384 -13686 -21674 -12976 sw
tri -21674 -13686 -20964 -12976 ne
tri -20964 -13686 -17428 -10150 sw
tri 20758 -10356 22000 -9114 se
rect 22000 -10150 24500 10150
rect 22000 -10356 23966 -10150
rect -24841 -14055 -21674 -13686
rect -28550 -14221 -25550 -14055
tri -25550 -14221 -25384 -14055 sw
tri -24841 -14221 -24675 -14055 ne
rect -24675 -14220 -21674 -14055
tri -21674 -14220 -21140 -13686 sw
tri -20964 -14220 -20430 -13686 ne
rect -20430 -14220 -17428 -13686
rect -24675 -14221 -21140 -14220
rect -28550 -14591 -25384 -14221
rect -32263 -15124 -29260 -14591
tri -36508 -18660 -32972 -15124 ne
tri -32972 -15833 -32263 -15124 sw
tri -32263 -15833 -31554 -15124 ne
rect -31554 -15301 -29260 -15124
tri -29260 -15301 -28550 -14591 sw
tri -28550 -15301 -27840 -14591 ne
rect -27840 -14930 -25384 -14591
tri -25384 -14930 -24675 -14221 sw
tri -24675 -14930 -23966 -14221 ne
rect -23966 -14930 -21140 -14221
tri -21140 -14930 -20430 -14220 sw
tri -20430 -14930 -19720 -14220 ne
rect -19720 -14930 -17428 -14220
rect -27840 -15301 -24675 -14930
rect -31554 -15463 -28550 -15301
tri -28550 -15463 -28388 -15301 sw
tri -27840 -15463 -27678 -15301 ne
rect -27678 -15463 -24675 -15301
rect -31554 -15833 -28388 -15463
rect -32972 -16542 -32263 -15833
tri -32263 -16542 -31554 -15833 sw
tri -31554 -16542 -30845 -15833 ne
rect -30845 -16173 -28388 -15833
tri -28388 -16173 -27678 -15463 sw
tri -27678 -16173 -26968 -15463 ne
rect -26968 -15464 -24675 -15463
tri -24675 -15464 -24141 -14930 sw
tri -23966 -15464 -23432 -14930 ne
rect -23432 -15464 -20430 -14930
rect -26968 -16173 -24141 -15464
tri -24141 -16173 -23432 -15464 sw
tri -23432 -16173 -22723 -15464 ne
rect -22723 -15640 -20430 -15464
tri -20430 -15640 -19720 -14930 sw
tri -19720 -15640 -19010 -14930 ne
rect -19010 -15640 -17428 -14930
rect -22723 -16173 -19720 -15640
rect -30845 -16542 -27678 -16173
rect -32972 -16708 -31554 -16542
tri -31554 -16708 -31388 -16542 sw
tri -30845 -16708 -30679 -16542 ne
rect -30679 -16707 -27678 -16542
tri -27678 -16707 -27144 -16173 sw
tri -26968 -16707 -26434 -16173 ne
rect -26434 -16707 -23432 -16173
rect -30679 -16708 -27144 -16707
rect -32972 -17417 -31388 -16708
tri -31388 -17417 -30679 -16708 sw
tri -30679 -17417 -29970 -16708 ne
rect -29970 -17417 -27144 -16708
tri -27144 -17417 -26434 -16707 sw
tri -26434 -17417 -25724 -16707 ne
rect -25724 -16882 -23432 -16707
tri -23432 -16882 -22723 -16173 sw
tri -22723 -16882 -22014 -16173 ne
rect -22014 -16350 -19720 -16173
tri -19720 -16350 -19010 -15640 sw
tri -19010 -16350 -18300 -15640 ne
rect -18300 -16350 -17428 -15640
rect -22014 -16512 -19010 -16350
tri -19010 -16512 -18848 -16350 sw
tri -18300 -16512 -18138 -16350 ne
rect -18138 -16512 -17428 -16350
rect -22014 -16882 -18848 -16512
rect -25724 -17417 -22723 -16882
rect -32972 -17951 -30679 -17417
tri -30679 -17951 -30145 -17417 sw
tri -29970 -17951 -29436 -17417 ne
rect -29436 -17951 -26434 -17417
rect -32972 -18660 -30145 -17951
tri -30145 -18660 -29436 -17951 sw
tri -29436 -18660 -28727 -17951 ne
rect -28727 -18127 -26434 -17951
tri -26434 -18127 -25724 -17417 sw
tri -25724 -18127 -25014 -17417 ne
rect -25014 -17591 -22723 -17417
tri -22723 -17591 -22014 -16882 sw
tri -22014 -17591 -21305 -16882 ne
rect -21305 -17222 -18848 -16882
tri -18848 -17222 -18138 -16512 sw
tri -18138 -17222 -17428 -16512 ne
tri -17428 -17222 -13892 -13686 sw
tri 17222 -13892 20758 -10356 se
rect 20758 -10684 23966 -10356
tri 23966 -10684 24500 -10150 nw
tri 24676 -10684 25002 -10358 se
rect 25002 -10684 27502 10684
rect 20758 -11394 23256 -10684
tri 23256 -11394 23966 -10684 nw
tri 23966 -11394 24676 -10684 se
rect 24676 -11394 27502 -10684
rect 20758 -12104 22546 -11394
tri 22546 -12104 23256 -11394 nw
tri 23256 -12104 23966 -11394 se
rect 23966 -11928 26968 -11394
tri 26968 -11928 27502 -11394 nw
tri 27677 -11928 28004 -11601 se
rect 28004 -11928 30504 11928
rect 23966 -12104 26259 -11928
rect 20758 -12648 22002 -12104
tri 22002 -12648 22546 -12104 nw
tri 22712 -12648 23256 -12104 se
rect 23256 -12637 26259 -12104
tri 26259 -12637 26968 -11928 nw
tri 26968 -12637 27677 -11928 se
rect 27677 -12637 30504 -11928
rect 23256 -12648 26072 -12637
rect 20758 -13358 21292 -12648
tri 21292 -13358 22002 -12648 nw
tri 22002 -13358 22712 -12648 se
rect 22712 -12824 26072 -12648
tri 26072 -12824 26259 -12637 nw
tri 26781 -12824 26968 -12637 se
rect 26968 -12824 29970 -12637
rect 22712 -13358 25363 -12824
tri 20758 -13892 21292 -13358 nw
tri 21468 -13892 22002 -13358 se
rect 22002 -13533 25363 -13358
tri 25363 -13533 26072 -12824 nw
tri 26072 -13533 26781 -12824 se
rect 26781 -13171 29970 -12824
tri 29970 -13171 30504 -12637 nw
tri 30680 -13171 31006 -12845 se
rect 31006 -13171 33506 13171
rect 34008 5500 36508 14415
rect 34008 3000 37508 5500
rect 26781 -13533 29260 -13171
rect 22002 -13881 25015 -13533
tri 25015 -13881 25363 -13533 nw
tri 25724 -13881 26072 -13533 se
rect 26072 -13881 29260 -13533
tri 29260 -13881 29970 -13171 nw
tri 29970 -13881 30680 -13171 se
rect 30680 -13881 33506 -13171
rect 22002 -13892 24306 -13881
rect -21305 -17591 -18138 -17222
rect -25014 -17757 -22014 -17591
tri -22014 -17757 -21848 -17591 sw
tri -21305 -17757 -21139 -17591 ne
rect -21139 -17756 -18138 -17591
tri -18138 -17756 -17604 -17222 sw
tri -17428 -17756 -16894 -17222 ne
rect -16894 -17756 -13892 -17222
rect -21139 -17757 -17604 -17756
rect -25014 -18127 -21848 -17757
rect -28727 -18660 -25724 -18127
tri -32972 -22196 -29436 -18660 ne
tri -29436 -19369 -28727 -18660 sw
tri -28727 -19369 -28018 -18660 ne
rect -28018 -18837 -25724 -18660
tri -25724 -18837 -25014 -18127 sw
tri -25014 -18837 -24304 -18127 ne
rect -24304 -18466 -21848 -18127
tri -21848 -18466 -21139 -17757 sw
tri -21139 -18466 -20430 -17757 ne
rect -20430 -18466 -17604 -17757
tri -17604 -18466 -16894 -17756 sw
tri -16894 -18466 -16184 -17756 ne
rect -16184 -18466 -13892 -17756
rect -24304 -18837 -21139 -18466
rect -28018 -18999 -25014 -18837
tri -25014 -18999 -24852 -18837 sw
tri -24304 -18999 -24142 -18837 ne
rect -24142 -18999 -21139 -18837
rect -28018 -19369 -24852 -18999
rect -29436 -20078 -28727 -19369
tri -28727 -20078 -28018 -19369 sw
tri -28018 -20078 -27309 -19369 ne
rect -27309 -19709 -24852 -19369
tri -24852 -19709 -24142 -18999 sw
tri -24142 -19709 -23432 -18999 ne
rect -23432 -19000 -21139 -18999
tri -21139 -19000 -20605 -18466 sw
tri -20430 -19000 -19896 -18466 ne
rect -19896 -19000 -16894 -18466
rect -23432 -19709 -20605 -19000
tri -20605 -19709 -19896 -19000 sw
tri -19896 -19709 -19187 -19000 ne
rect -19187 -19176 -16894 -19000
tri -16894 -19176 -16184 -18466 sw
tri -16184 -19176 -15474 -18466 ne
rect -15474 -19176 -13892 -18466
rect -19187 -19709 -16184 -19176
rect -27309 -20078 -24142 -19709
rect -29436 -20244 -28018 -20078
tri -28018 -20244 -27852 -20078 sw
tri -27309 -20244 -27143 -20078 ne
rect -27143 -20243 -24142 -20078
tri -24142 -20243 -23608 -19709 sw
tri -23432 -20243 -22898 -19709 ne
rect -22898 -20243 -19896 -19709
rect -27143 -20244 -23608 -20243
rect -29436 -20953 -27852 -20244
tri -27852 -20953 -27143 -20244 sw
tri -27143 -20953 -26434 -20244 ne
rect -26434 -20953 -23608 -20244
tri -23608 -20953 -22898 -20243 sw
tri -22898 -20953 -22188 -20243 ne
rect -22188 -20418 -19896 -20243
tri -19896 -20418 -19187 -19709 sw
tri -19187 -20418 -18478 -19709 ne
rect -18478 -19886 -16184 -19709
tri -16184 -19886 -15474 -19176 sw
tri -15474 -19886 -14764 -19176 ne
rect -14764 -19886 -13892 -19176
rect -18478 -20048 -15474 -19886
tri -15474 -20048 -15312 -19886 sw
tri -14764 -20048 -14602 -19886 ne
rect -14602 -20048 -13892 -19886
rect -18478 -20418 -15312 -20048
rect -22188 -20953 -19187 -20418
rect -29436 -21487 -27143 -20953
tri -27143 -21487 -26609 -20953 sw
tri -26434 -21487 -25900 -20953 ne
rect -25900 -21487 -22898 -20953
rect -29436 -22196 -26609 -21487
tri -26609 -22196 -25900 -21487 sw
tri -25900 -22196 -25191 -21487 ne
rect -25191 -21663 -22898 -21487
tri -22898 -21663 -22188 -20953 sw
tri -22188 -21663 -21478 -20953 ne
rect -21478 -21127 -19187 -20953
tri -19187 -21127 -18478 -20418 sw
tri -18478 -21127 -17769 -20418 ne
rect -17769 -20758 -15312 -20418
tri -15312 -20758 -14602 -20048 sw
tri -14602 -20758 -13892 -20048 ne
tri -13892 -20758 -10356 -17222 sw
tri 13686 -17428 17222 -13892 se
rect 17222 -14602 20048 -13892
tri 20048 -14602 20758 -13892 nw
tri 20758 -14602 21468 -13892 se
rect 21468 -14590 24306 -13892
tri 24306 -14590 25015 -13881 nw
tri 25015 -14590 25724 -13881 se
rect 25724 -14590 28550 -13881
rect 21468 -14602 23954 -14590
rect 17222 -15312 19338 -14602
tri 19338 -15312 20048 -14602 nw
tri 20048 -15312 20758 -14602 se
rect 20758 -14942 23954 -14602
tri 23954 -14942 24306 -14590 nw
tri 24663 -14942 25015 -14590 se
rect 25015 -14591 28550 -14590
tri 28550 -14591 29260 -13881 nw
tri 29260 -14591 29970 -13881 se
rect 29970 -14415 32972 -13881
tri 32972 -14415 33506 -13881 nw
rect 34008 -5500 37508 -3000
tri 33681 -14415 34008 -14088 se
rect 34008 -14415 36508 -5500
rect 29970 -14591 32263 -14415
rect 25015 -14942 28025 -14591
rect 20758 -15312 23245 -14942
rect 17222 -15474 19176 -15312
tri 19176 -15474 19338 -15312 nw
tri 19886 -15474 20048 -15312 se
rect 20048 -15474 23245 -15312
rect 17222 -16184 18466 -15474
tri 18466 -16184 19176 -15474 nw
tri 19176 -16184 19886 -15474 se
rect 19886 -15651 23245 -15474
tri 23245 -15651 23954 -14942 nw
tri 23954 -15651 24663 -14942 se
rect 24663 -15116 28025 -14942
tri 28025 -15116 28550 -14591 nw
rect 24663 -15651 27315 -15116
rect 19886 -16184 22536 -15651
rect 17222 -16894 17756 -16184
tri 17756 -16894 18466 -16184 nw
tri 18466 -16894 19176 -16184 se
rect 19176 -16360 22536 -16184
tri 22536 -16360 23245 -15651 nw
tri 23245 -16360 23954 -15651 se
rect 23954 -15826 27315 -15651
tri 27315 -15826 28025 -15116 nw
tri 28727 -15124 29260 -14591 se
rect 29260 -15124 32263 -14591
tri 32263 -15124 32972 -14415 nw
tri 32972 -15124 33681 -14415 se
rect 33681 -15124 36508 -14415
tri 28025 -15826 28727 -15124 se
rect 28727 -15826 31561 -15124
tri 31561 -15826 32263 -15124 nw
tri 32804 -15292 32972 -15124 se
rect 32972 -15292 36340 -15124
tri 36340 -15292 36508 -15124 nw
tri 32270 -15826 32804 -15292 se
rect 23954 -16360 26781 -15826
tri 26781 -16360 27315 -15826 nw
tri 27491 -16360 28025 -15826 se
rect 28025 -16360 30852 -15826
rect 19176 -16894 22002 -16360
tri 22002 -16894 22536 -16360 nw
tri 22711 -16894 23245 -16360 se
rect 23245 -16894 26071 -16360
tri 17222 -17428 17756 -16894 nw
tri 17932 -17428 18466 -16894 se
rect 18466 -17428 21293 -16894
rect -17769 -21127 -14602 -20758
rect -21478 -21293 -18478 -21127
tri -18478 -21293 -18312 -21127 sw
tri -17769 -21293 -17603 -21127 ne
rect -17603 -21292 -14602 -21127
tri -14602 -21292 -14068 -20758 sw
tri -13892 -21292 -13358 -20758 ne
rect -13358 -21292 -10356 -20758
rect -17603 -21293 -14068 -21292
rect -21478 -21663 -18312 -21293
rect -25191 -22196 -22188 -21663
tri -29436 -25732 -25900 -22196 ne
tri -25900 -22905 -25191 -22196 sw
tri -25191 -22905 -24482 -22196 ne
rect -24482 -22373 -22188 -22196
tri -22188 -22373 -21478 -21663 sw
tri -21478 -22373 -20768 -21663 ne
rect -20768 -22002 -18312 -21663
tri -18312 -22002 -17603 -21293 sw
tri -17603 -22002 -16894 -21293 ne
rect -16894 -22002 -14068 -21293
tri -14068 -22002 -13358 -21292 sw
tri -13358 -22002 -12648 -21292 ne
rect -12648 -22000 -10356 -21292
tri -10356 -22000 -9114 -20758 sw
tri 10150 -20964 13686 -17428 se
rect 13686 -18138 16512 -17428
tri 16512 -18138 17222 -17428 nw
tri 17222 -18138 17932 -17428 se
rect 17932 -17603 21293 -17428
tri 21293 -17603 22002 -16894 nw
tri 22002 -17603 22711 -16894 se
rect 22711 -17070 26071 -16894
tri 26071 -17070 26781 -16360 nw
tri 26781 -17070 27491 -16360 se
rect 27491 -16535 30852 -16360
tri 30852 -16535 31561 -15826 nw
tri 31561 -16535 32270 -15826 se
rect 32270 -16535 32804 -15826
rect 27491 -17070 30143 -16535
rect 22711 -17603 25361 -17070
rect 17932 -18138 20584 -17603
rect 13686 -18848 15802 -18138
tri 15802 -18848 16512 -18138 nw
tri 16512 -18848 17222 -18138 se
rect 17222 -18312 20584 -18138
tri 20584 -18312 21293 -17603 nw
tri 21293 -18312 22002 -17603 se
rect 22002 -17780 25361 -17603
tri 25361 -17780 26071 -17070 nw
tri 26071 -17780 26781 -17070 se
rect 26781 -17244 30143 -17070
tri 30143 -17244 30852 -16535 nw
tri 30852 -17244 31561 -16535 se
rect 31561 -17244 32804 -16535
rect 26781 -17410 29977 -17244
tri 29977 -17410 30143 -17244 nw
tri 30686 -17410 30852 -17244 se
rect 30852 -17410 32804 -17244
rect 26781 -17780 29268 -17410
rect 22002 -17942 25199 -17780
tri 25199 -17942 25361 -17780 nw
tri 25909 -17942 26071 -17780 se
rect 26071 -17942 29268 -17780
rect 22002 -18312 24489 -17942
rect 17222 -18478 20418 -18312
tri 20418 -18478 20584 -18312 nw
tri 21127 -18478 21293 -18312 se
rect 21293 -18478 24489 -18312
rect 17222 -18848 19709 -18478
rect 13686 -19010 15640 -18848
tri 15640 -19010 15802 -18848 nw
tri 16350 -19010 16512 -18848 se
rect 16512 -19010 19709 -18848
rect 13686 -19720 14930 -19010
tri 14930 -19720 15640 -19010 nw
tri 15640 -19720 16350 -19010 se
rect 16350 -19187 19709 -19010
tri 19709 -19187 20418 -18478 nw
tri 20418 -19187 21127 -18478 se
rect 21127 -18652 24489 -18478
tri 24489 -18652 25199 -17942 nw
tri 25199 -18652 25909 -17942 se
rect 25909 -18119 29268 -17942
tri 29268 -18119 29977 -17410 nw
tri 29977 -18119 30686 -17410 se
rect 30686 -18119 32804 -17410
rect 25909 -18652 28559 -18119
rect 21127 -19187 23779 -18652
rect 16350 -19720 19000 -19187
rect 13686 -20430 14220 -19720
tri 14220 -20430 14930 -19720 nw
tri 14930 -20430 15640 -19720 se
rect 15640 -19896 19000 -19720
tri 19000 -19896 19709 -19187 nw
tri 19709 -19896 20418 -19187 se
rect 20418 -19362 23779 -19187
tri 23779 -19362 24489 -18652 nw
tri 24489 -19362 25199 -18652 se
rect 25199 -18828 28559 -18652
tri 28559 -18828 29268 -18119 nw
tri 29268 -18828 29977 -18119 se
rect 29977 -18828 32804 -18119
tri 32804 -18828 36340 -15292 nw
rect 25199 -19362 28025 -18828
tri 28025 -19362 28559 -18828 nw
tri 28734 -19362 29268 -18828 se
rect 20418 -19896 23245 -19362
tri 23245 -19896 23779 -19362 nw
tri 23955 -19896 24489 -19362 se
rect 24489 -19896 27316 -19362
rect 15640 -20430 18466 -19896
tri 18466 -20430 19000 -19896 nw
tri 19175 -20430 19709 -19896 se
rect 19709 -20430 22535 -19896
tri 13686 -20964 14220 -20430 nw
tri 14396 -20964 14930 -20430 se
rect 14930 -20964 17757 -20430
tri 9114 -22000 10150 -20964 se
rect 10150 -21674 12976 -20964
tri 12976 -21674 13686 -20964 nw
tri 13686 -21674 14396 -20964 se
rect 14396 -21139 17757 -20964
tri 17757 -21139 18466 -20430 nw
tri 18466 -21139 19175 -20430 se
rect 19175 -20606 22535 -20430
tri 22535 -20606 23245 -19896 nw
tri 23245 -20606 23955 -19896 se
rect 23955 -20071 27316 -19896
tri 27316 -20071 28025 -19362 nw
tri 28025 -20071 28734 -19362 se
rect 28734 -20071 29268 -19362
rect 23955 -20606 26607 -20071
rect 19175 -21139 21825 -20606
rect 14396 -21674 17048 -21139
rect 10150 -22000 12266 -21674
rect -12648 -22002 12266 -22000
rect -20768 -22373 -17603 -22002
rect -24482 -22535 -21478 -22373
tri -21478 -22535 -21316 -22373 sw
tri -20768 -22535 -20606 -22373 ne
rect -20606 -22535 -17603 -22373
rect -24482 -22905 -21316 -22535
rect -25900 -23614 -25191 -22905
tri -25191 -23614 -24482 -22905 sw
tri -24482 -23614 -23773 -22905 ne
rect -23773 -23245 -21316 -22905
tri -21316 -23245 -20606 -22535 sw
tri -20606 -23245 -19896 -22535 ne
rect -19896 -22536 -17603 -22535
tri -17603 -22536 -17069 -22002 sw
tri -16894 -22536 -16360 -22002 ne
rect -16360 -22536 -13358 -22002
rect -19896 -23245 -17069 -22536
tri -17069 -23245 -16360 -22536 sw
tri -16360 -23245 -15651 -22536 ne
rect -15651 -22712 -13358 -22536
tri -13358 -22712 -12648 -22002 sw
tri -12648 -22712 -11938 -22002 ne
rect -11938 -22384 12266 -22002
tri 12266 -22384 12976 -21674 nw
tri 12976 -22384 13686 -21674 se
rect 13686 -21848 17048 -21674
tri 17048 -21848 17757 -21139 nw
tri 17757 -21848 18466 -21139 se
rect 18466 -21316 21825 -21139
tri 21825 -21316 22535 -20606 nw
tri 22535 -21316 23245 -20606 se
rect 23245 -20780 26607 -20606
tri 26607 -20780 27316 -20071 nw
tri 27316 -20780 28025 -20071 se
rect 28025 -20780 29268 -20071
rect 23245 -20946 26441 -20780
tri 26441 -20946 26607 -20780 nw
tri 27150 -20946 27316 -20780 se
rect 27316 -20946 29268 -20780
rect 23245 -21316 25732 -20946
rect 18466 -21478 21663 -21316
tri 21663 -21478 21825 -21316 nw
tri 22373 -21478 22535 -21316 se
rect 22535 -21478 25732 -21316
rect 18466 -21848 20953 -21478
rect 13686 -22014 16882 -21848
tri 16882 -22014 17048 -21848 nw
tri 17591 -22014 17757 -21848 se
rect 17757 -22014 20953 -21848
rect 13686 -22384 16173 -22014
rect -11938 -22546 12104 -22384
tri 12104 -22546 12266 -22384 nw
tri 12814 -22546 12976 -22384 se
rect 12976 -22546 16173 -22384
rect -11938 -22712 11394 -22546
rect -15651 -23245 -12648 -22712
rect -23773 -23614 -20606 -23245
rect -25900 -23780 -24482 -23614
tri -24482 -23780 -24316 -23614 sw
tri -23773 -23780 -23607 -23614 ne
rect -23607 -23779 -20606 -23614
tri -20606 -23779 -20072 -23245 sw
tri -19896 -23779 -19362 -23245 ne
rect -19362 -23779 -16360 -23245
rect -23607 -23780 -20072 -23779
rect -25900 -24489 -24316 -23780
tri -24316 -24489 -23607 -23780 sw
tri -23607 -24489 -22898 -23780 ne
rect -22898 -24489 -20072 -23780
tri -20072 -24489 -19362 -23779 sw
tri -19362 -24489 -18652 -23779 ne
rect -18652 -23954 -16360 -23779
tri -16360 -23954 -15651 -23245 sw
tri -15651 -23954 -14942 -23245 ne
rect -14942 -23256 -12648 -23245
tri -12648 -23256 -12104 -22712 sw
tri -11938 -23256 -11394 -22712 ne
rect -11394 -23256 11394 -22712
tri 11394 -23256 12104 -22546 nw
tri 12104 -23256 12814 -22546 se
rect 12814 -22723 16173 -22546
tri 16173 -22723 16882 -22014 nw
tri 16882 -22723 17591 -22014 se
rect 17591 -22188 20953 -22014
tri 20953 -22188 21663 -21478 nw
tri 21663 -22188 22373 -21478 se
rect 22373 -21655 25732 -21478
tri 25732 -21655 26441 -20946 nw
tri 26441 -21655 27150 -20946 se
rect 27150 -21655 29268 -20946
rect 22373 -22188 25023 -21655
rect 17591 -22723 20243 -22188
rect 12814 -23256 15464 -22723
rect -14942 -23954 -12104 -23256
rect -18652 -24489 -15651 -23954
rect -25900 -25023 -23607 -24489
tri -23607 -25023 -23073 -24489 sw
tri -22898 -25023 -22364 -24489 ne
rect -22364 -25023 -19362 -24489
rect -25900 -25732 -23073 -25023
tri -23073 -25732 -22364 -25023 sw
tri -22364 -25732 -21655 -25023 ne
rect -21655 -25199 -19362 -25023
tri -19362 -25199 -18652 -24489 sw
tri -18652 -25199 -17942 -24489 ne
rect -17942 -24663 -15651 -24489
tri -15651 -24663 -14942 -23954 sw
tri -14942 -24663 -14233 -23954 ne
rect -14233 -23966 -12104 -23954
tri -12104 -23966 -11394 -23256 sw
tri -11394 -23966 -10684 -23256 ne
rect -10684 -23966 10684 -23256
tri 10684 -23966 11394 -23256 nw
tri 11394 -23966 12104 -23256 se
rect 12104 -23432 15464 -23256
tri 15464 -23432 16173 -22723 nw
tri 16173 -23432 16882 -22723 se
rect 16882 -22898 20243 -22723
tri 20243 -22898 20953 -22188 nw
tri 20953 -22898 21663 -22188 se
rect 21663 -22364 25023 -22188
tri 25023 -22364 25732 -21655 nw
tri 25732 -22364 26441 -21655 se
rect 26441 -22364 29268 -21655
tri 29268 -22364 32804 -18828 nw
rect 21663 -22898 24489 -22364
tri 24489 -22898 25023 -22364 nw
tri 25198 -22898 25732 -22364 se
rect 16882 -23432 19709 -22898
tri 19709 -23432 20243 -22898 nw
tri 20419 -23432 20953 -22898 se
rect 20953 -23432 23780 -22898
rect 12104 -23966 14930 -23432
tri 14930 -23966 15464 -23432 nw
tri 15639 -23966 16173 -23432 se
rect 16173 -23966 18999 -23432
rect -14233 -24500 -11394 -23966
tri -11394 -24500 -10860 -23966 sw
tri -10684 -24500 -10150 -23966 ne
rect -10150 -24500 10150 -23966
tri 10150 -24500 10684 -23966 nw
tri 10860 -24500 11394 -23966 se
rect 11394 -24500 14221 -23966
rect -14233 -24663 -10860 -24500
rect -17942 -24829 -14942 -24663
tri -14942 -24829 -14776 -24663 sw
tri -14233 -24829 -14067 -24663 ne
rect -14067 -24829 -10860 -24663
rect -17942 -25199 -14776 -24829
rect -21655 -25732 -18652 -25199
tri -25900 -29268 -22364 -25732 ne
tri -22364 -26441 -21655 -25732 sw
tri -21655 -26441 -20946 -25732 ne
rect -20946 -25909 -18652 -25732
tri -18652 -25909 -17942 -25199 sw
tri -17942 -25909 -17232 -25199 ne
rect -17232 -25538 -14776 -25199
tri -14776 -25538 -14067 -24829 sw
tri -14067 -25538 -13358 -24829 ne
rect -13358 -25002 -10860 -24829
tri -10860 -25002 -10358 -24500 sw
tri 10358 -25002 10860 -24500 se
rect 10860 -24675 14221 -24500
tri 14221 -24675 14930 -23966 nw
tri 14930 -24675 15639 -23966 se
rect 15639 -24142 18999 -23966
tri 18999 -24142 19709 -23432 nw
tri 19709 -24142 20419 -23432 se
rect 20419 -23607 23780 -23432
tri 23780 -23607 24489 -22898 nw
tri 24489 -23607 25198 -22898 se
rect 25198 -23607 25732 -22898
rect 20419 -24142 23071 -23607
rect 15639 -24675 18289 -24142
rect 10860 -25002 13512 -24675
rect -13358 -25538 -979 -25002
rect -17232 -25909 -14067 -25538
rect -20946 -26071 -17942 -25909
tri -17942 -26071 -17780 -25909 sw
tri -17232 -26071 -17070 -25909 ne
rect -17070 -26071 -14067 -25909
rect -20946 -26441 -17780 -26071
rect -22364 -27150 -21655 -26441
tri -21655 -27150 -20946 -26441 sw
tri -20946 -27150 -20237 -26441 ne
rect -20237 -26781 -17780 -26441
tri -17780 -26781 -17070 -26071 sw
tri -17070 -26781 -16360 -26071 ne
rect -16360 -26072 -14067 -26071
tri -14067 -26072 -13533 -25538 sw
tri -13358 -26072 -12824 -25538 ne
rect -12824 -26072 -979 -25538
rect -16360 -26781 -13533 -26072
tri -13533 -26781 -12824 -26072 sw
tri -12824 -26781 -12115 -26072 ne
rect -12115 -26781 -979 -26072
rect -20237 -27150 -17070 -26781
rect -22364 -27316 -20946 -27150
tri -20946 -27316 -20780 -27150 sw
tri -20237 -27316 -20071 -27150 ne
rect -20071 -27315 -17070 -27150
tri -17070 -27315 -16536 -26781 sw
tri -16360 -27315 -15826 -26781 ne
rect -15826 -27315 -12824 -26781
rect -20071 -27316 -16536 -27315
rect -22364 -28025 -20780 -27316
tri -20780 -28025 -20071 -27316 sw
tri -20071 -28025 -19362 -27316 ne
rect -19362 -28025 -16536 -27316
tri -16536 -28025 -15826 -27315 sw
tri -15826 -28025 -15116 -27315 ne
rect -15116 -27490 -12824 -27315
tri -12824 -27490 -12115 -26781 sw
tri -12115 -27490 -11406 -26781 ne
rect -11406 -27490 -979 -26781
rect -15116 -27502 -12115 -27490
tri -12115 -27502 -12103 -27490 sw
tri -11406 -27502 -11394 -27490 ne
rect -11394 -27502 -979 -27490
tri -979 -27502 1521 -25002 sw
tri 2291 -25222 2511 -25002 se
rect 2511 -25222 13512 -25002
rect 2291 -25324 13512 -25222
rect 2291 -25580 2393 -25324
rect 2649 -25580 2917 -25324
rect 3173 -25580 3471 -25324
rect 3727 -25580 4025 -25324
rect 4281 -25580 4549 -25324
rect 4805 -25580 5163 -25324
rect 5419 -25580 5687 -25324
rect 5943 -25580 6241 -25324
rect 6497 -25580 6795 -25324
rect 7051 -25580 7319 -25324
rect 7575 -25384 13512 -25324
tri 13512 -25384 14221 -24675 nw
tri 14221 -25384 14930 -24675 se
rect 14930 -24852 18289 -24675
tri 18289 -24852 18999 -24142 nw
tri 18999 -24852 19709 -24142 se
rect 19709 -24316 23071 -24142
tri 23071 -24316 23780 -23607 nw
tri 23780 -24316 24489 -23607 se
rect 24489 -24316 25732 -23607
rect 19709 -24482 22905 -24316
tri 22905 -24482 23071 -24316 nw
tri 23614 -24482 23780 -24316 se
rect 23780 -24482 25732 -24316
rect 19709 -24852 22196 -24482
rect 14930 -25014 18127 -24852
tri 18127 -25014 18289 -24852 nw
tri 18837 -25014 18999 -24852 se
rect 18999 -25014 22196 -24852
rect 14930 -25384 17417 -25014
rect 7575 -25550 13346 -25384
tri 13346 -25550 13512 -25384 nw
tri 14055 -25550 14221 -25384 se
rect 14221 -25550 17417 -25384
rect 7575 -25580 12637 -25550
rect 2291 -25818 12637 -25580
rect 2291 -26074 2393 -25818
rect 2649 -26074 2917 -25818
rect 3173 -26074 3471 -25818
rect 3727 -26074 4025 -25818
rect 4281 -26074 4549 -25818
rect 4805 -26074 5163 -25818
rect 5419 -26074 5687 -25818
rect 5943 -26074 6241 -25818
rect 6497 -26074 6795 -25818
rect 7051 -26074 7319 -25818
rect 7575 -26074 12637 -25818
rect 2291 -26259 12637 -26074
tri 12637 -26259 13346 -25550 nw
tri 13346 -26259 14055 -25550 se
rect 14055 -25724 17417 -25550
tri 17417 -25724 18127 -25014 nw
tri 18127 -25724 18837 -25014 se
rect 18837 -25191 22196 -25014
tri 22196 -25191 22905 -24482 nw
tri 22905 -25191 23614 -24482 se
rect 23614 -25191 25732 -24482
rect 18837 -25724 21487 -25191
rect 14055 -26259 16707 -25724
rect 2291 -26432 11928 -26259
rect 2291 -26688 2393 -26432
rect 2649 -26688 2917 -26432
rect 3173 -26688 3471 -26432
rect 3727 -26688 4025 -26432
rect 4281 -26688 4549 -26432
rect 4805 -26688 5163 -26432
rect 5419 -26688 5687 -26432
rect 5943 -26688 6241 -26432
rect 6497 -26688 6795 -26432
rect 7051 -26688 7319 -26432
rect 7575 -26688 11928 -26432
rect 2291 -26926 11928 -26688
rect 2291 -27182 2393 -26926
rect 2649 -27182 2917 -26926
rect 3173 -27182 3471 -26926
rect 3727 -27182 4025 -26926
rect 4281 -27182 4549 -26926
rect 4805 -27182 5163 -26926
rect 5419 -27182 5687 -26926
rect 5943 -27182 6241 -26926
rect 6497 -27182 6795 -26926
rect 7051 -27182 7319 -26926
rect 7575 -26968 11928 -26926
tri 11928 -26968 12637 -26259 nw
tri 12637 -26968 13346 -26259 se
rect 13346 -26434 16707 -26259
tri 16707 -26434 17417 -25724 nw
tri 17417 -26434 18127 -25724 se
rect 18127 -25900 21487 -25724
tri 21487 -25900 22196 -25191 nw
tri 22196 -25900 22905 -25191 se
rect 22905 -25900 25732 -25191
tri 25732 -25900 29268 -22364 nw
rect 18127 -26434 20953 -25900
tri 20953 -26434 21487 -25900 nw
tri 21662 -26434 22196 -25900 se
rect 13346 -26968 16173 -26434
tri 16173 -26968 16707 -26434 nw
tri 16883 -26968 17417 -26434 se
rect 17417 -26968 20244 -26434
rect 7575 -27182 11394 -26968
rect 2291 -27282 11394 -27182
tri 2291 -27502 2511 -27282 ne
rect 2511 -27502 11394 -27282
tri 11394 -27502 11928 -26968 nw
tri 12103 -27502 12637 -26968 se
rect 12637 -27502 15463 -26968
rect -15116 -28004 -12103 -27502
tri -12103 -28004 -11601 -27502 sw
rect -15116 -28025 -2380 -28004
rect -22364 -28559 -20071 -28025
tri -20071 -28559 -19537 -28025 sw
tri -19362 -28559 -18828 -28025 ne
rect -18828 -28559 -15826 -28025
rect -22364 -29268 -19537 -28559
tri -19537 -29268 -18828 -28559 sw
tri -18828 -29268 -18119 -28559 ne
rect -18119 -28735 -15826 -28559
tri -15826 -28735 -15116 -28025 sw
tri -15116 -28735 -14406 -28025 ne
rect -14406 -28224 -2380 -28025
tri -2380 -28224 -2160 -28004 sw
rect -14406 -28325 -2160 -28224
rect -14406 -28581 -7444 -28325
rect -7188 -28581 -6920 -28325
rect -6664 -28581 -6366 -28325
rect -6110 -28581 -5812 -28325
rect -5556 -28581 -5288 -28325
rect -5032 -28581 -4674 -28325
rect -4418 -28581 -4150 -28325
rect -3894 -28581 -3596 -28325
rect -3340 -28581 -3042 -28325
rect -2786 -28581 -2518 -28325
rect -2262 -28581 -2160 -28325
rect -14406 -28735 -2160 -28581
rect -18119 -29260 -15116 -28735
tri -15116 -29260 -14591 -28735 sw
tri -14406 -29260 -13881 -28735 ne
rect -13881 -28819 -2160 -28735
rect -13881 -29075 -7444 -28819
rect -7188 -29075 -6920 -28819
rect -6664 -29075 -6366 -28819
rect -6110 -29075 -5812 -28819
rect -5556 -29075 -5288 -28819
rect -5032 -29075 -4674 -28819
rect -4418 -29075 -4150 -28819
rect -3894 -29075 -3596 -28819
rect -3340 -29075 -3042 -28819
rect -2786 -29075 -2518 -28819
rect -2262 -29075 -2160 -28819
rect -13881 -29260 -2160 -29075
rect -18119 -29268 -14591 -29260
tri -22364 -32804 -18828 -29268 ne
tri -18828 -29977 -18119 -29268 sw
tri -18119 -29977 -17410 -29268 ne
rect -17410 -29970 -14591 -29268
tri -14591 -29970 -13881 -29260 sw
tri -13881 -29970 -13171 -29260 ne
rect -13171 -29433 -2160 -29260
rect -13171 -29689 -7444 -29433
rect -7188 -29689 -6920 -29433
rect -6664 -29689 -6366 -29433
rect -6110 -29689 -5812 -29433
rect -5556 -29689 -5288 -29433
rect -5032 -29689 -4674 -29433
rect -4418 -29689 -4150 -29433
rect -3894 -29689 -3596 -29433
rect -3340 -29689 -3042 -29433
rect -2786 -29689 -2518 -29433
rect -2262 -29689 -2160 -29433
rect -13171 -29927 -2160 -29689
rect -13171 -29970 -7444 -29927
rect -17410 -29977 -13881 -29970
rect -18828 -30686 -18119 -29977
tri -18119 -30686 -17410 -29977 sw
tri -17410 -30686 -16701 -29977 ne
rect -16701 -30504 -13881 -29977
tri -13881 -30504 -13347 -29970 sw
tri -13171 -30504 -12637 -29970 ne
rect -12637 -30183 -7444 -29970
rect -7188 -30183 -6920 -29927
rect -6664 -30183 -6366 -29927
rect -6110 -30183 -5812 -29927
rect -5556 -30183 -5288 -29927
rect -5032 -30183 -4674 -29927
rect -4418 -30183 -4150 -29927
rect -3894 -30183 -3596 -29927
rect -3340 -30183 -3042 -29927
rect -2786 -30183 -2518 -29927
rect -2262 -30183 -2160 -29927
rect -12637 -30284 -2160 -30183
rect -12637 -30504 -2380 -30284
tri -2380 -30504 -2160 -30284 nw
tri -2015 -30504 987 -27502 ne
rect 987 -28004 1521 -27502
tri 1521 -28004 2023 -27502 sw
tri 11601 -28004 12103 -27502 se
rect 12103 -27678 15463 -27502
tri 15463 -27678 16173 -26968 nw
tri 16173 -27678 16883 -26968 se
rect 16883 -27143 20244 -26968
tri 20244 -27143 20953 -26434 nw
tri 20953 -27143 21662 -26434 se
rect 21662 -27143 22196 -26434
rect 16883 -27678 19535 -27143
rect 12103 -28004 14753 -27678
rect 987 -28388 14753 -28004
tri 14753 -28388 15463 -27678 nw
tri 15463 -28388 16173 -27678 se
rect 16173 -27852 19535 -27678
tri 19535 -27852 20244 -27143 nw
tri 20244 -27852 20953 -27143 se
rect 20953 -27852 22196 -27143
rect 16173 -28018 19369 -27852
tri 19369 -28018 19535 -27852 nw
tri 20078 -28018 20244 -27852 se
rect 20244 -28018 22196 -27852
rect 16173 -28388 18660 -28018
rect 987 -28550 14591 -28388
tri 14591 -28550 14753 -28388 nw
tri 15301 -28550 15463 -28388 se
rect 15463 -28550 18660 -28388
rect 987 -29260 13881 -28550
tri 13881 -29260 14591 -28550 nw
tri 14591 -29260 15301 -28550 se
rect 15301 -28727 18660 -28550
tri 18660 -28727 19369 -28018 nw
tri 19369 -28727 20078 -28018 se
rect 20078 -28727 22196 -28018
rect 15301 -29260 17951 -28727
rect 987 -29970 13171 -29260
tri 13171 -29970 13881 -29260 nw
tri 13881 -29970 14591 -29260 se
rect 14591 -29436 17951 -29260
tri 17951 -29436 18660 -28727 nw
tri 18660 -29436 19369 -28727 se
rect 19369 -29436 22196 -28727
tri 22196 -29436 25732 -25900 nw
rect 14591 -29970 17417 -29436
tri 17417 -29970 17951 -29436 nw
tri 18126 -29970 18660 -29436 se
rect 987 -30504 12637 -29970
tri 12637 -30504 13171 -29970 nw
tri 13347 -30504 13881 -29970 se
rect 13881 -30504 16708 -29970
rect -16701 -30686 -13347 -30504
rect -18828 -30852 -17410 -30686
tri -17410 -30852 -17244 -30686 sw
tri -16701 -30852 -16535 -30686 ne
rect -16535 -30852 -13347 -30686
rect -18828 -31561 -17244 -30852
tri -17244 -31561 -16535 -30852 sw
tri -16535 -31561 -15826 -30852 ne
rect -15826 -31006 -13347 -30852
tri -13347 -31006 -12845 -30504 sw
tri 12845 -31006 13347 -30504 se
rect 13347 -30679 16708 -30504
tri 16708 -30679 17417 -29970 nw
tri 17417 -30679 18126 -29970 se
rect 18126 -30679 18660 -29970
rect 13347 -31006 15999 -30679
rect -15826 -31561 -979 -31006
rect -18828 -32095 -16535 -31561
tri -16535 -32095 -16001 -31561 sw
tri -15826 -32095 -15292 -31561 ne
rect -15292 -32095 -979 -31561
rect -18828 -32804 -16001 -32095
tri -16001 -32804 -15292 -32095 sw
tri -15292 -32804 -14583 -32095 ne
rect -14583 -32804 -979 -32095
tri -18828 -36340 -15292 -32804 ne
tri -15292 -33506 -14590 -32804 sw
tri -14583 -33506 -13881 -32804 ne
rect -13881 -33506 -979 -32804
tri -979 -33506 1521 -31006 sw
tri 2291 -31226 2511 -31006 se
rect 2511 -31226 15999 -31006
rect 2291 -31326 15999 -31226
rect 2291 -31582 2393 -31326
rect 2649 -31582 2917 -31326
rect 3173 -31582 3471 -31326
rect 3727 -31582 4025 -31326
rect 4281 -31582 4549 -31326
rect 4805 -31582 5163 -31326
rect 5419 -31582 5687 -31326
rect 5943 -31582 6241 -31326
rect 6497 -31582 6795 -31326
rect 7051 -31582 7319 -31326
rect 7575 -31388 15999 -31326
tri 15999 -31388 16708 -30679 nw
tri 16708 -31388 17417 -30679 se
rect 17417 -31388 18660 -30679
rect 7575 -31554 15833 -31388
tri 15833 -31554 15999 -31388 nw
tri 16542 -31554 16708 -31388 se
rect 16708 -31554 18660 -31388
rect 7575 -31582 15124 -31554
rect 2291 -31820 15124 -31582
rect 2291 -32076 2393 -31820
rect 2649 -32076 2917 -31820
rect 3173 -32076 3471 -31820
rect 3727 -32076 4025 -31820
rect 4281 -32076 4549 -31820
rect 4805 -32076 5163 -31820
rect 5419 -32076 5687 -31820
rect 5943 -32076 6241 -31820
rect 6497 -32076 6795 -31820
rect 7051 -32076 7319 -31820
rect 7575 -32076 15124 -31820
rect 2291 -32263 15124 -32076
tri 15124 -32263 15833 -31554 nw
tri 15833 -32263 16542 -31554 se
rect 16542 -32263 18660 -31554
rect 2291 -32434 14415 -32263
rect 2291 -32690 2393 -32434
rect 2649 -32690 2917 -32434
rect 3173 -32690 3471 -32434
rect 3727 -32690 4025 -32434
rect 4281 -32690 4549 -32434
rect 4805 -32690 5163 -32434
rect 5419 -32690 5687 -32434
rect 5943 -32690 6241 -32434
rect 6497 -32690 6795 -32434
rect 7051 -32690 7319 -32434
rect 7575 -32690 14415 -32434
rect 2291 -32928 14415 -32690
rect 2291 -33184 2393 -32928
rect 2649 -33184 2917 -32928
rect 3173 -33184 3471 -32928
rect 3727 -33184 4025 -32928
rect 4281 -33184 4549 -32928
rect 4805 -33184 5163 -32928
rect 5419 -33184 5687 -32928
rect 5943 -33184 6241 -32928
rect 6497 -33184 6795 -32928
rect 7051 -33184 7319 -32928
rect 7575 -32972 14415 -32928
tri 14415 -32972 15124 -32263 nw
tri 15124 -32972 15833 -32263 se
rect 15833 -32972 18660 -32263
tri 18660 -32972 22196 -29436 nw
rect 7575 -33184 13881 -32972
rect 2291 -33286 13881 -33184
tri 2291 -33506 2511 -33286 ne
rect 2511 -33506 13881 -33286
tri 13881 -33506 14415 -32972 nw
tri 14590 -33506 15124 -32972 se
rect -15292 -34008 -14590 -33506
tri -14590 -34008 -14088 -33506 sw
rect -15292 -34228 -2380 -34008
tri -2380 -34228 -2160 -34008 sw
rect -15292 -34329 -2160 -34228
rect -15292 -34585 -7444 -34329
rect -7188 -34585 -6920 -34329
rect -6664 -34585 -6366 -34329
rect -6110 -34585 -5812 -34329
rect -5556 -34585 -5288 -34329
rect -5032 -34585 -4674 -34329
rect -4418 -34585 -4150 -34329
rect -3894 -34585 -3596 -34329
rect -3340 -34585 -3042 -34329
rect -2786 -34585 -2518 -34329
rect -2262 -34585 -2160 -34329
rect -15292 -34823 -2160 -34585
rect -15292 -35079 -7444 -34823
rect -7188 -35079 -6920 -34823
rect -6664 -35079 -6366 -34823
rect -6110 -35079 -5812 -34823
rect -5556 -35079 -5288 -34823
rect -5032 -35079 -4674 -34823
rect -4418 -35079 -4150 -34823
rect -3894 -35079 -3596 -34823
rect -3340 -35079 -3042 -34823
rect -2786 -35079 -2518 -34823
rect -2262 -35079 -2160 -34823
rect -15292 -35437 -2160 -35079
rect -15292 -35693 -7444 -35437
rect -7188 -35693 -6920 -35437
rect -6664 -35693 -6366 -35437
rect -6110 -35693 -5812 -35437
rect -5556 -35693 -5288 -35437
rect -5032 -35693 -4674 -35437
rect -4418 -35693 -4150 -35437
rect -3894 -35693 -3596 -35437
rect -3340 -35693 -3042 -35437
rect -2786 -35693 -2518 -35437
rect -2262 -35693 -2160 -35437
rect -15292 -35931 -2160 -35693
rect -15292 -36187 -7444 -35931
rect -7188 -36187 -6920 -35931
rect -6664 -36187 -6366 -35931
rect -6110 -36187 -5812 -35931
rect -5556 -36187 -5288 -35931
rect -5032 -36187 -4674 -35931
rect -4418 -36187 -4150 -35931
rect -3894 -36187 -3596 -35931
rect -3340 -36187 -3042 -35931
rect -2786 -36187 -2518 -35931
rect -2262 -36187 -2160 -35931
rect -15292 -36288 -2160 -36187
rect -15292 -36340 -2380 -36288
tri -15292 -36508 -15124 -36340 ne
rect -15124 -36508 -2380 -36340
tri -2380 -36508 -2160 -36288 nw
tri -2015 -36508 987 -33506 ne
rect 987 -34008 1521 -33506
tri 1521 -34008 2023 -33506 sw
tri 14088 -34008 14590 -33506 se
rect 14590 -34008 15124 -33506
rect 987 -36508 15124 -34008
tri 15124 -36508 18660 -32972 nw
<< comment >>
tri -15125 15126 -6267 36508 ne
rect -6267 15125 6266 36508
tri 6266 15125 15125 36508 nw
tri -36508 6266 -15125 15125 sw
tri -6267 6266 -2596 15125 ne
rect -2596 6266 2596 15125
tri 2596 6266 6266 15125 nw
tri 15125 6266 36508 15125 se
rect -36508 1075 -15125 6266
tri -15125 1075 -2596 6266 sw
tri -2596 1076 -446 6266 ne
rect -446 1075 445 6266
tri 445 1075 2596 6266 nw
tri 2596 1075 15125 6266 se
rect 15125 1075 36508 6266
rect -36508 185 -2596 1075
tri -2596 185 -446 1075 sw
tri -446 185 -77 1075 ne
rect -77 1074 445 1075
tri 2594 1074 2596 1075 se
rect 2596 1074 36508 1075
rect -77 185 76 1074
rect -36508 32 -446 185
tri -446 32 -77 185 sw
tri -77 33 -14 185 ne
rect -14 183 76 185
tri 76 184 445 1074 nw
tri 445 184 2594 1074 se
rect 2594 184 36508 1074
tri 443 183 445 184 se
rect 445 183 36508 184
rect -14 32 13 183
rect -36508 6 -77 32
tri -77 6 -14 32 sw
tri -14 6 -3 32 ne
rect -3 31 13 32
tri 13 31 76 183 nw
tri 76 31 443 183 se
rect 443 31 36508 183
rect -3 6 2 31
rect -36508 1 -14 6
tri -14 1 -3 6 sw
tri -3 2 -1 6 ne
rect -1 5 2 6
tri 2 5 13 31 nw
tri 13 5 76 31 se
rect 76 5 36508 31
rect -1 1 0 5
tri 0 1 2 5 nw
tri 2 1 13 5 se
rect 13 1 36508 5
rect -36508 0 -3 1
tri -3 0 -1 1 sw
tri -1 0 0 1 ne
tri 0 0 2 1 se
rect 2 0 36508 1
rect -36508 -1 -2 0
tri -2 -1 0 0 nw
tri 0 -1 1 0 ne
rect 1 -1 36508 0
rect -36508 -5 -13 -1
tri -13 -5 -2 -1 nw
tri -2 -5 0 -1 se
tri 0 -3 1 -1 sw
tri 2 -3 6 -1 ne
rect 6 -3 36508 -1
rect 0 -5 1 -3
rect -36508 -31 -76 -5
tri -76 -31 -13 -5 nw
tri -13 -31 -2 -5 se
rect -2 -14 1 -5
tri 1 -14 6 -3 sw
tri 6 -14 32 -3 ne
rect 32 -14 36508 -3
rect -2 -31 6 -14
rect -36508 -183 -443 -31
tri -443 -183 -76 -31 nw
tri -76 -183 -13 -31 se
rect -13 -77 6 -31
tri 6 -77 32 -14 sw
tri 33 -77 185 -14 ne
rect 185 -77 36508 -14
rect -13 -183 32 -77
rect -36508 -184 -445 -183
tri -445 -184 -443 -183 nw
rect -36508 -1074 -2594 -184
tri -2594 -1074 -445 -184 nw
tri -445 -1074 -76 -184 se
rect -76 -446 32 -183
tri 32 -446 185 -77 sw
tri 185 -446 1075 -77 ne
rect 1075 -446 36508 -77
rect -76 -1074 185 -446
rect -36508 -1075 -2596 -1074
tri -2596 -1075 -2594 -1074 nw
rect -36508 -6266 -15125 -1075
tri -15125 -6266 -2596 -1075 nw
tri -2596 -6266 -445 -1075 se
rect -445 -2596 185 -1074
tri 185 -2596 1075 -446 sw
tri 1076 -2596 6266 -446 ne
rect 6266 -2596 36508 -446
rect -445 -6266 1075 -2596
tri -36508 -15125 -15125 -6266 nw
tri -6266 -15125 -2596 -6266 se
rect -2596 -15125 1075 -6266
tri 1075 -15125 6266 -2596 sw
tri 6266 -15125 36508 -2596 ne
tri -15125 -36508 -6266 -15125 se
rect -6266 -36508 6266 -15125
tri 6266 -36508 15125 -15125 sw
<< properties >>
string GDS_END 10442368
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 10411100
string gencell sky130_fd_pr__rf_test_coil3
string library sky130
string parameter m=1
string path 881.450 -378.100 881.450 -75.000 
<< end >>
