magic
tech sky130B
magscale 1 2
timestamp 1676037725
<< dnwell >>
rect 80 80 1644 1644
<< nwell >>
rect 0 1364 1724 1724
rect 0 360 360 1364
rect 1364 360 1724 1364
rect 0 0 1724 360
<< pbase >>
rect 360 360 1364 1364
<< npn1p00 >>
rect 360 360 1364 1364
<< ndiff >>
rect 762 947 962 962
rect 762 777 777 947
rect 947 777 962 947
rect 762 762 962 777
<< ndiffc >>
rect 777 777 947 947
<< psubdiff >>
rect 520 1180 1204 1204
rect 520 1146 544 1180
rect 578 1146 641 1180
rect 675 1146 709 1180
rect 743 1146 777 1180
rect 811 1146 845 1180
rect 879 1146 913 1180
rect 947 1146 981 1180
rect 1015 1146 1049 1180
rect 1083 1146 1146 1180
rect 1180 1146 1204 1180
rect 520 1122 1204 1146
rect 520 1083 602 1122
rect 520 1049 544 1083
rect 578 1049 602 1083
rect 520 1015 602 1049
rect 520 981 544 1015
rect 578 981 602 1015
rect 520 947 602 981
rect 1122 1083 1204 1122
rect 1122 1049 1146 1083
rect 1180 1049 1204 1083
rect 1122 1015 1204 1049
rect 1122 981 1146 1015
rect 1180 981 1204 1015
rect 520 913 544 947
rect 578 913 602 947
rect 520 879 602 913
rect 520 845 544 879
rect 578 845 602 879
rect 520 811 602 845
rect 520 777 544 811
rect 578 777 602 811
rect 520 743 602 777
rect 1122 947 1204 981
rect 1122 913 1146 947
rect 1180 913 1204 947
rect 1122 879 1204 913
rect 1122 845 1146 879
rect 1180 845 1204 879
rect 1122 811 1204 845
rect 1122 777 1146 811
rect 1180 777 1204 811
rect 520 709 544 743
rect 578 709 602 743
rect 520 675 602 709
rect 520 641 544 675
rect 578 641 602 675
rect 520 602 602 641
rect 1122 743 1204 777
rect 1122 709 1146 743
rect 1180 709 1204 743
rect 1122 675 1204 709
rect 1122 641 1146 675
rect 1180 641 1204 675
rect 1122 602 1204 641
rect 520 578 1204 602
rect 520 544 544 578
rect 578 544 641 578
rect 675 544 709 578
rect 743 544 777 578
rect 811 544 845 578
rect 879 544 913 578
rect 947 544 981 578
rect 1015 544 1049 578
rect 1083 544 1146 578
rect 1180 544 1204 578
rect 520 520 1204 544
<< nsubdiff >>
rect 118 1582 1606 1606
rect 118 1548 142 1582
rect 176 1548 233 1582
rect 267 1548 301 1582
rect 335 1548 369 1582
rect 403 1548 437 1582
rect 471 1548 505 1582
rect 539 1548 573 1582
rect 607 1548 641 1582
rect 675 1548 709 1582
rect 743 1548 777 1582
rect 811 1548 845 1582
rect 879 1548 913 1582
rect 947 1548 981 1582
rect 1015 1548 1049 1582
rect 1083 1548 1117 1582
rect 1151 1548 1185 1582
rect 1219 1548 1253 1582
rect 1287 1548 1321 1582
rect 1355 1548 1389 1582
rect 1423 1548 1457 1582
rect 1491 1548 1548 1582
rect 1582 1548 1606 1582
rect 118 1524 1606 1548
rect 118 1491 200 1524
rect 118 1457 142 1491
rect 176 1457 200 1491
rect 118 1423 200 1457
rect 118 1389 142 1423
rect 176 1389 200 1423
rect 118 1355 200 1389
rect 118 1321 142 1355
rect 176 1321 200 1355
rect 118 1287 200 1321
rect 118 1253 142 1287
rect 176 1253 200 1287
rect 118 1219 200 1253
rect 118 1185 142 1219
rect 176 1185 200 1219
rect 1524 1491 1606 1524
rect 1524 1457 1548 1491
rect 1582 1457 1606 1491
rect 1524 1423 1606 1457
rect 1524 1389 1548 1423
rect 1582 1389 1606 1423
rect 1524 1355 1606 1389
rect 1524 1321 1548 1355
rect 1582 1321 1606 1355
rect 1524 1287 1606 1321
rect 1524 1253 1548 1287
rect 1582 1253 1606 1287
rect 1524 1219 1606 1253
rect 118 1151 200 1185
rect 118 1117 142 1151
rect 176 1117 200 1151
rect 118 1083 200 1117
rect 118 1049 142 1083
rect 176 1049 200 1083
rect 118 1015 200 1049
rect 118 981 142 1015
rect 176 981 200 1015
rect 118 947 200 981
rect 118 913 142 947
rect 176 913 200 947
rect 118 879 200 913
rect 118 845 142 879
rect 176 845 200 879
rect 118 811 200 845
rect 118 777 142 811
rect 176 777 200 811
rect 118 743 200 777
rect 118 709 142 743
rect 176 709 200 743
rect 118 675 200 709
rect 118 641 142 675
rect 176 641 200 675
rect 118 607 200 641
rect 118 573 142 607
rect 176 573 200 607
rect 118 539 200 573
rect 118 505 142 539
rect 176 505 200 539
rect 1524 1185 1548 1219
rect 1582 1185 1606 1219
rect 1524 1151 1606 1185
rect 1524 1117 1548 1151
rect 1582 1117 1606 1151
rect 1524 1083 1606 1117
rect 1524 1049 1548 1083
rect 1582 1049 1606 1083
rect 1524 1015 1606 1049
rect 1524 981 1548 1015
rect 1582 981 1606 1015
rect 1524 947 1606 981
rect 1524 913 1548 947
rect 1582 913 1606 947
rect 1524 879 1606 913
rect 1524 845 1548 879
rect 1582 845 1606 879
rect 1524 811 1606 845
rect 1524 777 1548 811
rect 1582 777 1606 811
rect 1524 743 1606 777
rect 1524 709 1548 743
rect 1582 709 1606 743
rect 1524 675 1606 709
rect 1524 641 1548 675
rect 1582 641 1606 675
rect 1524 607 1606 641
rect 1524 573 1548 607
rect 1582 573 1606 607
rect 1524 539 1606 573
rect 118 471 200 505
rect 118 437 142 471
rect 176 437 200 471
rect 118 403 200 437
rect 118 369 142 403
rect 176 369 200 403
rect 118 335 200 369
rect 118 301 142 335
rect 176 301 200 335
rect 118 267 200 301
rect 118 233 142 267
rect 176 233 200 267
rect 118 200 200 233
rect 1524 505 1548 539
rect 1582 505 1606 539
rect 1524 471 1606 505
rect 1524 437 1548 471
rect 1582 437 1606 471
rect 1524 403 1606 437
rect 1524 369 1548 403
rect 1582 369 1606 403
rect 1524 335 1606 369
rect 1524 301 1548 335
rect 1582 301 1606 335
rect 1524 267 1606 301
rect 1524 233 1548 267
rect 1582 233 1606 267
rect 1524 200 1606 233
rect 118 176 1606 200
rect 118 142 142 176
rect 176 142 233 176
rect 267 142 301 176
rect 335 142 369 176
rect 403 142 437 176
rect 471 142 505 176
rect 539 142 573 176
rect 607 142 641 176
rect 675 142 709 176
rect 743 142 777 176
rect 811 142 845 176
rect 879 142 913 176
rect 947 142 981 176
rect 1015 142 1049 176
rect 1083 142 1117 176
rect 1151 142 1185 176
rect 1219 142 1253 176
rect 1287 142 1321 176
rect 1355 142 1389 176
rect 1423 142 1457 176
rect 1491 142 1548 176
rect 1582 142 1606 176
rect 118 118 1606 142
<< psubdiffcont >>
rect 544 1146 578 1180
rect 641 1146 675 1180
rect 709 1146 743 1180
rect 777 1146 811 1180
rect 845 1146 879 1180
rect 913 1146 947 1180
rect 981 1146 1015 1180
rect 1049 1146 1083 1180
rect 1146 1146 1180 1180
rect 544 1049 578 1083
rect 544 981 578 1015
rect 1146 1049 1180 1083
rect 1146 981 1180 1015
rect 544 913 578 947
rect 544 845 578 879
rect 544 777 578 811
rect 1146 913 1180 947
rect 1146 845 1180 879
rect 1146 777 1180 811
rect 544 709 578 743
rect 544 641 578 675
rect 1146 709 1180 743
rect 1146 641 1180 675
rect 544 544 578 578
rect 641 544 675 578
rect 709 544 743 578
rect 777 544 811 578
rect 845 544 879 578
rect 913 544 947 578
rect 981 544 1015 578
rect 1049 544 1083 578
rect 1146 544 1180 578
<< nsubdiffcont >>
rect 142 1548 176 1582
rect 233 1548 267 1582
rect 301 1548 335 1582
rect 369 1548 403 1582
rect 437 1548 471 1582
rect 505 1548 539 1582
rect 573 1548 607 1582
rect 641 1548 675 1582
rect 709 1548 743 1582
rect 777 1548 811 1582
rect 845 1548 879 1582
rect 913 1548 947 1582
rect 981 1548 1015 1582
rect 1049 1548 1083 1582
rect 1117 1548 1151 1582
rect 1185 1548 1219 1582
rect 1253 1548 1287 1582
rect 1321 1548 1355 1582
rect 1389 1548 1423 1582
rect 1457 1548 1491 1582
rect 1548 1548 1582 1582
rect 142 1457 176 1491
rect 142 1389 176 1423
rect 142 1321 176 1355
rect 142 1253 176 1287
rect 142 1185 176 1219
rect 1548 1457 1582 1491
rect 1548 1389 1582 1423
rect 1548 1321 1582 1355
rect 1548 1253 1582 1287
rect 142 1117 176 1151
rect 142 1049 176 1083
rect 142 981 176 1015
rect 142 913 176 947
rect 142 845 176 879
rect 142 777 176 811
rect 142 709 176 743
rect 142 641 176 675
rect 142 573 176 607
rect 142 505 176 539
rect 1548 1185 1582 1219
rect 1548 1117 1582 1151
rect 1548 1049 1582 1083
rect 1548 981 1582 1015
rect 1548 913 1582 947
rect 1548 845 1582 879
rect 1548 777 1582 811
rect 1548 709 1582 743
rect 1548 641 1582 675
rect 1548 573 1582 607
rect 142 437 176 471
rect 142 369 176 403
rect 142 301 176 335
rect 142 233 176 267
rect 1548 505 1582 539
rect 1548 437 1582 471
rect 1548 369 1582 403
rect 1548 301 1582 335
rect 1548 233 1582 267
rect 142 142 176 176
rect 233 142 267 176
rect 301 142 335 176
rect 369 142 403 176
rect 437 142 471 176
rect 505 142 539 176
rect 573 142 607 176
rect 641 142 675 176
rect 709 142 743 176
rect 777 142 811 176
rect 845 142 879 176
rect 913 142 947 176
rect 981 142 1015 176
rect 1049 142 1083 176
rect 1117 142 1151 176
rect 1185 142 1219 176
rect 1253 142 1287 176
rect 1321 142 1355 176
rect 1389 142 1423 176
rect 1457 142 1491 176
rect 1548 142 1582 176
<< locali >>
rect 126 1582 1598 1598
rect 126 1548 142 1582
rect 176 1548 233 1582
rect 267 1548 301 1582
rect 339 1548 369 1582
rect 411 1548 437 1582
rect 483 1548 505 1582
rect 555 1548 573 1582
rect 627 1548 641 1582
rect 699 1548 709 1582
rect 771 1548 777 1582
rect 843 1548 845 1582
rect 879 1548 881 1582
rect 947 1548 953 1582
rect 1015 1548 1025 1582
rect 1083 1548 1097 1582
rect 1151 1548 1169 1582
rect 1219 1548 1241 1582
rect 1287 1548 1313 1582
rect 1355 1548 1385 1582
rect 1423 1548 1457 1582
rect 1491 1548 1548 1582
rect 1582 1548 1598 1582
rect 126 1532 1598 1548
rect 126 1491 192 1532
rect 126 1457 142 1491
rect 176 1457 192 1491
rect 126 1423 192 1457
rect 126 1385 142 1423
rect 176 1385 192 1423
rect 126 1355 192 1385
rect 126 1313 142 1355
rect 176 1313 192 1355
rect 126 1287 192 1313
rect 126 1241 142 1287
rect 176 1241 192 1287
rect 126 1219 192 1241
rect 126 1169 142 1219
rect 176 1169 192 1219
rect 1532 1491 1598 1532
rect 1532 1457 1548 1491
rect 1582 1457 1598 1491
rect 1532 1423 1598 1457
rect 1532 1385 1548 1423
rect 1582 1385 1598 1423
rect 1532 1355 1598 1385
rect 1532 1313 1548 1355
rect 1582 1313 1598 1355
rect 1532 1287 1598 1313
rect 1532 1241 1548 1287
rect 1582 1241 1598 1287
rect 1532 1219 1598 1241
rect 126 1151 192 1169
rect 126 1097 142 1151
rect 176 1097 192 1151
rect 126 1083 192 1097
rect 126 1025 142 1083
rect 176 1025 192 1083
rect 126 1015 192 1025
rect 126 953 142 1015
rect 176 953 192 1015
rect 126 947 192 953
rect 126 881 142 947
rect 176 881 192 947
rect 126 879 192 881
rect 126 845 142 879
rect 176 845 192 879
rect 126 843 192 845
rect 126 777 142 843
rect 176 777 192 843
rect 126 771 192 777
rect 126 709 142 771
rect 176 709 192 771
rect 126 699 192 709
rect 126 641 142 699
rect 176 641 192 699
rect 126 627 192 641
rect 126 573 142 627
rect 176 573 192 627
rect 126 555 192 573
rect 126 505 142 555
rect 176 505 192 555
rect 528 1180 1196 1196
rect 528 1146 544 1180
rect 578 1146 629 1180
rect 675 1146 701 1180
rect 743 1146 773 1180
rect 811 1146 845 1180
rect 879 1146 913 1180
rect 951 1146 981 1180
rect 1023 1146 1049 1180
rect 1095 1146 1146 1180
rect 1180 1146 1196 1180
rect 528 1130 1196 1146
rect 528 1095 594 1130
rect 528 1049 544 1095
rect 578 1049 594 1095
rect 528 1023 594 1049
rect 528 981 544 1023
rect 578 981 594 1023
rect 528 951 594 981
rect 1130 1095 1196 1130
rect 1130 1049 1146 1095
rect 1180 1049 1196 1095
rect 1130 1023 1196 1049
rect 1130 981 1146 1023
rect 1180 981 1196 1023
rect 528 913 544 951
rect 578 913 594 951
rect 528 879 594 913
rect 528 845 544 879
rect 578 845 594 879
rect 528 811 594 845
rect 528 773 544 811
rect 578 773 594 811
rect 528 743 594 773
rect 761 951 963 963
rect 761 773 773 951
rect 951 773 963 951
rect 761 761 963 773
rect 1130 951 1196 981
rect 1130 913 1146 951
rect 1180 913 1196 951
rect 1130 879 1196 913
rect 1130 845 1146 879
rect 1180 845 1196 879
rect 1130 811 1196 845
rect 1130 773 1146 811
rect 1180 773 1196 811
rect 528 701 544 743
rect 578 701 594 743
rect 528 675 594 701
rect 528 629 544 675
rect 578 629 594 675
rect 528 594 594 629
rect 1130 743 1196 773
rect 1130 701 1146 743
rect 1180 701 1196 743
rect 1130 675 1196 701
rect 1130 629 1146 675
rect 1180 629 1196 675
rect 1130 594 1196 629
rect 528 578 1196 594
rect 528 544 544 578
rect 578 544 629 578
rect 675 544 701 578
rect 743 544 773 578
rect 811 544 845 578
rect 879 544 913 578
rect 951 544 981 578
rect 1023 544 1049 578
rect 1095 544 1146 578
rect 1180 544 1196 578
rect 528 528 1196 544
rect 1532 1169 1548 1219
rect 1582 1169 1598 1219
rect 1532 1151 1598 1169
rect 1532 1097 1548 1151
rect 1582 1097 1598 1151
rect 1532 1083 1598 1097
rect 1532 1025 1548 1083
rect 1582 1025 1598 1083
rect 1532 1015 1598 1025
rect 1532 953 1548 1015
rect 1582 953 1598 1015
rect 1532 947 1598 953
rect 1532 881 1548 947
rect 1582 881 1598 947
rect 1532 879 1598 881
rect 1532 845 1548 879
rect 1582 845 1598 879
rect 1532 843 1598 845
rect 1532 777 1548 843
rect 1582 777 1598 843
rect 1532 771 1598 777
rect 1532 709 1548 771
rect 1582 709 1598 771
rect 1532 699 1598 709
rect 1532 641 1548 699
rect 1582 641 1598 699
rect 1532 627 1598 641
rect 1532 573 1548 627
rect 1582 573 1598 627
rect 1532 555 1598 573
rect 126 483 192 505
rect 126 437 142 483
rect 176 437 192 483
rect 126 411 192 437
rect 126 369 142 411
rect 176 369 192 411
rect 126 339 192 369
rect 126 301 142 339
rect 176 301 192 339
rect 126 267 192 301
rect 126 233 142 267
rect 176 233 192 267
rect 126 192 192 233
rect 1532 505 1548 555
rect 1582 505 1598 555
rect 1532 483 1598 505
rect 1532 437 1548 483
rect 1582 437 1598 483
rect 1532 411 1598 437
rect 1532 369 1548 411
rect 1582 369 1598 411
rect 1532 339 1598 369
rect 1532 301 1548 339
rect 1582 301 1598 339
rect 1532 267 1598 301
rect 1532 233 1548 267
rect 1582 233 1598 267
rect 1532 192 1598 233
rect 126 176 1598 192
rect 126 142 142 176
rect 176 142 233 176
rect 267 142 301 176
rect 339 142 369 176
rect 411 142 437 176
rect 483 142 505 176
rect 555 142 573 176
rect 627 142 641 176
rect 699 142 709 176
rect 771 142 777 176
rect 843 142 845 176
rect 879 142 881 176
rect 947 142 953 176
rect 1015 142 1025 176
rect 1083 142 1097 176
rect 1151 142 1169 176
rect 1219 142 1241 176
rect 1287 142 1313 176
rect 1355 142 1385 176
rect 1423 142 1457 176
rect 1491 142 1548 176
rect 1582 142 1598 176
rect 126 126 1598 142
<< viali >>
rect 142 1548 176 1582
rect 233 1548 267 1582
rect 305 1548 335 1582
rect 335 1548 339 1582
rect 377 1548 403 1582
rect 403 1548 411 1582
rect 449 1548 471 1582
rect 471 1548 483 1582
rect 521 1548 539 1582
rect 539 1548 555 1582
rect 593 1548 607 1582
rect 607 1548 627 1582
rect 665 1548 675 1582
rect 675 1548 699 1582
rect 737 1548 743 1582
rect 743 1548 771 1582
rect 809 1548 811 1582
rect 811 1548 843 1582
rect 881 1548 913 1582
rect 913 1548 915 1582
rect 953 1548 981 1582
rect 981 1548 987 1582
rect 1025 1548 1049 1582
rect 1049 1548 1059 1582
rect 1097 1548 1117 1582
rect 1117 1548 1131 1582
rect 1169 1548 1185 1582
rect 1185 1548 1203 1582
rect 1241 1548 1253 1582
rect 1253 1548 1275 1582
rect 1313 1548 1321 1582
rect 1321 1548 1347 1582
rect 1385 1548 1389 1582
rect 1389 1548 1419 1582
rect 1457 1548 1491 1582
rect 1548 1548 1582 1582
rect 142 1457 176 1491
rect 142 1389 176 1419
rect 142 1385 176 1389
rect 142 1321 176 1347
rect 142 1313 176 1321
rect 142 1253 176 1275
rect 142 1241 176 1253
rect 142 1185 176 1203
rect 142 1169 176 1185
rect 1548 1457 1582 1491
rect 1548 1389 1582 1419
rect 1548 1385 1582 1389
rect 1548 1321 1582 1347
rect 1548 1313 1582 1321
rect 1548 1253 1582 1275
rect 1548 1241 1582 1253
rect 142 1117 176 1131
rect 142 1097 176 1117
rect 142 1049 176 1059
rect 142 1025 176 1049
rect 142 981 176 987
rect 142 953 176 981
rect 142 913 176 915
rect 142 881 176 913
rect 142 811 176 843
rect 142 809 176 811
rect 142 743 176 771
rect 142 737 176 743
rect 142 675 176 699
rect 142 665 176 675
rect 142 607 176 627
rect 142 593 176 607
rect 142 539 176 555
rect 142 521 176 539
rect 544 1146 578 1180
rect 629 1146 641 1180
rect 641 1146 663 1180
rect 701 1146 709 1180
rect 709 1146 735 1180
rect 773 1146 777 1180
rect 777 1146 807 1180
rect 845 1146 879 1180
rect 917 1146 947 1180
rect 947 1146 951 1180
rect 989 1146 1015 1180
rect 1015 1146 1023 1180
rect 1061 1146 1083 1180
rect 1083 1146 1095 1180
rect 1146 1146 1180 1180
rect 544 1083 578 1095
rect 544 1061 578 1083
rect 544 1015 578 1023
rect 544 989 578 1015
rect 1146 1083 1180 1095
rect 1146 1061 1180 1083
rect 1146 1015 1180 1023
rect 1146 989 1180 1015
rect 544 947 578 951
rect 544 917 578 947
rect 544 845 578 879
rect 544 777 578 807
rect 544 773 578 777
rect 773 947 951 951
rect 773 777 777 947
rect 777 777 947 947
rect 947 777 951 947
rect 773 773 951 777
rect 1146 947 1180 951
rect 1146 917 1180 947
rect 1146 845 1180 879
rect 1146 777 1180 807
rect 1146 773 1180 777
rect 544 709 578 735
rect 544 701 578 709
rect 544 641 578 663
rect 544 629 578 641
rect 1146 709 1180 735
rect 1146 701 1180 709
rect 1146 641 1180 663
rect 1146 629 1180 641
rect 544 544 578 578
rect 629 544 641 578
rect 641 544 663 578
rect 701 544 709 578
rect 709 544 735 578
rect 773 544 777 578
rect 777 544 807 578
rect 845 544 879 578
rect 917 544 947 578
rect 947 544 951 578
rect 989 544 1015 578
rect 1015 544 1023 578
rect 1061 544 1083 578
rect 1083 544 1095 578
rect 1146 544 1180 578
rect 1548 1185 1582 1203
rect 1548 1169 1582 1185
rect 1548 1117 1582 1131
rect 1548 1097 1582 1117
rect 1548 1049 1582 1059
rect 1548 1025 1582 1049
rect 1548 981 1582 987
rect 1548 953 1582 981
rect 1548 913 1582 915
rect 1548 881 1582 913
rect 1548 811 1582 843
rect 1548 809 1582 811
rect 1548 743 1582 771
rect 1548 737 1582 743
rect 1548 675 1582 699
rect 1548 665 1582 675
rect 1548 607 1582 627
rect 1548 593 1582 607
rect 142 471 176 483
rect 142 449 176 471
rect 142 403 176 411
rect 142 377 176 403
rect 142 335 176 339
rect 142 305 176 335
rect 142 233 176 267
rect 1548 539 1582 555
rect 1548 521 1582 539
rect 1548 471 1582 483
rect 1548 449 1582 471
rect 1548 403 1582 411
rect 1548 377 1582 403
rect 1548 335 1582 339
rect 1548 305 1582 335
rect 1548 233 1582 267
rect 142 142 176 176
rect 233 142 267 176
rect 305 142 335 176
rect 335 142 339 176
rect 377 142 403 176
rect 403 142 411 176
rect 449 142 471 176
rect 471 142 483 176
rect 521 142 539 176
rect 539 142 555 176
rect 593 142 607 176
rect 607 142 627 176
rect 665 142 675 176
rect 675 142 699 176
rect 737 142 743 176
rect 743 142 771 176
rect 809 142 811 176
rect 811 142 843 176
rect 881 142 913 176
rect 913 142 915 176
rect 953 142 981 176
rect 981 142 987 176
rect 1025 142 1049 176
rect 1049 142 1059 176
rect 1097 142 1117 176
rect 1117 142 1131 176
rect 1169 142 1185 176
rect 1185 142 1203 176
rect 1241 142 1253 176
rect 1253 142 1275 176
rect 1313 142 1321 176
rect 1321 142 1347 176
rect 1385 142 1389 176
rect 1389 142 1419 176
rect 1457 142 1491 176
rect 1548 142 1582 176
<< metal1 >>
rect 130 1582 1594 1594
rect 130 1548 142 1582
rect 176 1548 233 1582
rect 267 1548 305 1582
rect 339 1548 377 1582
rect 411 1548 449 1582
rect 483 1548 521 1582
rect 555 1548 593 1582
rect 627 1548 665 1582
rect 699 1548 737 1582
rect 771 1548 809 1582
rect 843 1548 881 1582
rect 915 1548 953 1582
rect 987 1548 1025 1582
rect 1059 1548 1097 1582
rect 1131 1548 1169 1582
rect 1203 1548 1241 1582
rect 1275 1548 1313 1582
rect 1347 1548 1385 1582
rect 1419 1548 1457 1582
rect 1491 1548 1548 1582
rect 1582 1548 1594 1582
rect 130 1536 1594 1548
rect 130 1491 188 1536
rect 130 1457 142 1491
rect 176 1457 188 1491
rect 130 1419 188 1457
rect 130 1385 142 1419
rect 176 1385 188 1419
rect 130 1347 188 1385
rect 130 1313 142 1347
rect 176 1313 188 1347
rect 130 1275 188 1313
rect 130 1241 142 1275
rect 176 1241 188 1275
rect 130 1203 188 1241
rect 130 1169 142 1203
rect 176 1169 188 1203
rect 1536 1491 1594 1536
rect 1536 1457 1548 1491
rect 1582 1457 1594 1491
rect 1536 1419 1594 1457
rect 1536 1385 1548 1419
rect 1582 1385 1594 1419
rect 1536 1347 1594 1385
rect 1536 1313 1548 1347
rect 1582 1313 1594 1347
rect 1536 1275 1594 1313
rect 1536 1241 1548 1275
rect 1582 1241 1594 1275
rect 1536 1203 1594 1241
rect 130 1131 188 1169
rect 130 1097 142 1131
rect 176 1097 188 1131
rect 130 1059 188 1097
rect 130 1025 142 1059
rect 176 1025 188 1059
rect 130 987 188 1025
rect 130 953 142 987
rect 176 953 188 987
rect 130 915 188 953
rect 130 881 142 915
rect 176 881 188 915
rect 130 843 188 881
rect 130 809 142 843
rect 176 809 188 843
rect 130 771 188 809
rect 130 737 142 771
rect 176 737 188 771
rect 130 699 188 737
rect 130 665 142 699
rect 176 665 188 699
rect 130 627 188 665
rect 130 593 142 627
rect 176 593 188 627
rect 130 555 188 593
rect 130 521 142 555
rect 176 521 188 555
rect 532 1180 1192 1192
rect 532 1146 544 1180
rect 578 1146 629 1180
rect 663 1146 701 1180
rect 735 1146 773 1180
rect 807 1146 845 1180
rect 879 1146 917 1180
rect 951 1146 989 1180
rect 1023 1146 1061 1180
rect 1095 1146 1146 1180
rect 1180 1146 1192 1180
rect 532 1134 1192 1146
rect 532 1095 590 1134
rect 532 1061 544 1095
rect 578 1061 590 1095
rect 532 1023 590 1061
rect 532 989 544 1023
rect 578 989 590 1023
rect 532 951 590 989
rect 1134 1095 1192 1134
rect 1134 1061 1146 1095
rect 1180 1061 1192 1095
rect 1134 1023 1192 1061
rect 1134 989 1146 1023
rect 1180 989 1192 1023
rect 532 917 544 951
rect 578 917 590 951
rect 532 879 590 917
rect 532 845 544 879
rect 578 845 590 879
rect 532 807 590 845
rect 532 773 544 807
rect 578 773 590 807
rect 532 735 590 773
rect 761 951 963 963
rect 761 773 773 951
rect 951 773 963 951
rect 761 761 963 773
rect 1134 951 1192 989
rect 1134 917 1146 951
rect 1180 917 1192 951
rect 1134 879 1192 917
rect 1134 845 1146 879
rect 1180 845 1192 879
rect 1134 807 1192 845
rect 1134 773 1146 807
rect 1180 773 1192 807
rect 532 701 544 735
rect 578 701 590 735
rect 532 663 590 701
rect 532 629 544 663
rect 578 629 590 663
rect 532 590 590 629
rect 1134 735 1192 773
rect 1134 701 1146 735
rect 1180 701 1192 735
rect 1134 663 1192 701
rect 1134 629 1146 663
rect 1180 629 1192 663
rect 1134 590 1192 629
rect 532 578 1192 590
rect 532 544 544 578
rect 578 544 629 578
rect 663 544 701 578
rect 735 544 773 578
rect 807 544 845 578
rect 879 544 917 578
rect 951 544 989 578
rect 1023 544 1061 578
rect 1095 544 1146 578
rect 1180 544 1192 578
rect 532 532 1192 544
rect 1536 1169 1548 1203
rect 1582 1169 1594 1203
rect 1536 1131 1594 1169
rect 1536 1097 1548 1131
rect 1582 1097 1594 1131
rect 1536 1059 1594 1097
rect 1536 1025 1548 1059
rect 1582 1025 1594 1059
rect 1536 987 1594 1025
rect 1536 953 1548 987
rect 1582 953 1594 987
rect 1536 915 1594 953
rect 1536 881 1548 915
rect 1582 881 1594 915
rect 1536 843 1594 881
rect 1536 809 1548 843
rect 1582 809 1594 843
rect 1536 771 1594 809
rect 1536 737 1548 771
rect 1582 737 1594 771
rect 1536 699 1594 737
rect 1536 665 1548 699
rect 1582 665 1594 699
rect 1536 627 1594 665
rect 1536 593 1548 627
rect 1582 593 1594 627
rect 1536 555 1594 593
rect 130 483 188 521
rect 130 449 142 483
rect 176 449 188 483
rect 130 411 188 449
rect 130 377 142 411
rect 176 377 188 411
rect 130 339 188 377
rect 130 305 142 339
rect 176 305 188 339
rect 130 267 188 305
rect 130 233 142 267
rect 176 233 188 267
rect 130 188 188 233
rect 1536 521 1548 555
rect 1582 521 1594 555
rect 1536 483 1594 521
rect 1536 449 1548 483
rect 1582 449 1594 483
rect 1536 411 1594 449
rect 1536 377 1548 411
rect 1582 377 1594 411
rect 1536 339 1594 377
rect 1536 305 1548 339
rect 1582 305 1594 339
rect 1536 267 1594 305
rect 1536 233 1548 267
rect 1582 233 1594 267
rect 1536 188 1594 233
rect 130 176 1594 188
rect 130 142 142 176
rect 176 142 233 176
rect 267 142 305 176
rect 339 142 377 176
rect 411 142 449 176
rect 483 142 521 176
rect 555 142 593 176
rect 627 142 665 176
rect 699 142 737 176
rect 771 142 809 176
rect 843 142 881 176
rect 915 142 953 176
rect 987 142 1025 176
rect 1059 142 1097 176
rect 1131 142 1169 176
rect 1203 142 1241 176
rect 1275 142 1313 176
rect 1347 142 1385 176
rect 1419 142 1457 176
rect 1491 142 1548 176
rect 1582 142 1594 176
rect 130 130 1594 142
<< properties >>
string GDS_END 8739290
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 8717518
string gencell sky130_fd_pr__rf_npn_05v5_W1p00L1p00
string library sky130
string parameter m=1
string path 4.500 9.000 4.500 38.600 38.600 38.600 38.600 4.500 0.000 4.500 
<< end >>
