magic
tech sky130B
magscale 1 2
timestamp 1676037725
<< metal1 >>
tri 1870 16075 1904 16109 sw
tri 2723 16075 2731 16083 se
rect 1845 16047 2731 16075
tri 2697 16013 2731 16047 ne
rect 1870 15975 2649 16003
tri 1870 15923 1922 15975 nw
tri 2615 15941 2649 15975 ne
tri 2697 14974 2731 15008 se
tri 2122 14896 2156 14930 ne
rect 2406 14928 2788 14974
tri 1292 11234 1312 11254 sw
tri 1292 11154 1326 11188 nw
rect 3614 11164 3654 11200
tri 1240 11116 1250 11126 ne
rect 1250 11062 1282 11126
tri 1282 11116 1292 11126 nw
tri 1448 11106 1472 11130 sw
rect 3614 11106 3642 11164
tri 3772 11116 3783 11127 se
rect 3783 11116 4098 11127
rect 1448 11078 3642 11106
tri 3737 11081 3772 11116 se
rect 3772 11099 4098 11116
rect 3772 11081 3783 11099
tri 3783 11081 3801 11099 nw
tri 1250 11030 1282 11062 ne
tri 1282 11050 1308 11076 sw
tri 3706 11050 3737 11081 se
rect 3737 11050 3752 11081
tri 3752 11050 3783 11081 nw
rect 1282 11030 3724 11050
tri 1282 11022 1290 11030 ne
rect 1290 11022 3724 11030
tri 3724 11022 3752 11050 nw
tri 1085 10753 1235 10903 ne
tri 1292 10599 1322 10629 sw
tri 1949 10616 1993 10660 se
rect 1993 10632 2903 10660
tri 1993 10616 2009 10632 nw
tri 1905 10572 1949 10616 se
tri 1949 10572 1993 10616 nw
tri 1292 10519 1326 10553 nw
tri 1861 10528 1905 10572 se
tri 1905 10528 1949 10572 nw
tri 1200 10473 1228 10501 sw
tri 1817 10484 1861 10528 se
tri 1861 10484 1905 10528 nw
tri 1806 10473 1817 10484 se
rect 1817 10473 1822 10484
rect 1200 10445 1822 10473
tri 1822 10445 1861 10484 nw
tri 16397 2339 16403 2345 ne
tri 16531 2339 16537 2345 nw
tri 15136 1867 15142 1873 nw
tri 15252 1825 15301 1874 se
rect 15301 1825 15348 1873
rect 15262 1773 15348 1825
tri 15348 1773 15448 1873 nw
tri 14771 1209 14789 1227 se
tri 14982 1209 15000 1227 sw
tri 15247 1209 15379 1341 se
rect 15379 1213 16531 1341
rect 15379 1209 15391 1213
tri 15391 1209 15395 1213 nw
tri 14230 1079 14268 1117 sw
tri 15293 1111 15391 1209 nw
rect 14230 915 15502 1079
tri 16710 -367 16766 -311 se
rect 16123 -423 16766 -367
<< metal2 >>
tri 1295 16084 1345 16134 sw
tri 1754 16084 1818 16148 se
rect 1295 16047 1818 16084
rect 1379 15975 1818 16003
tri 1379 15919 1435 15975 nw
tri 1763 15920 1818 15975 ne
tri 2615 15090 2649 15124 se
tri 1717 11774 1719 11776 ne
rect 1719 11410 1835 11776
tri 1835 11741 1870 11776 nw
tri 1744 10819 1778 10853 se
tri 1834 10819 1868 10853 sw
rect 16095 7661 16390 7707
rect 16095 5106 16141 7661
tri 16141 5106 16161 5126 sw
tri 16095 5040 16161 5106 ne
tri 16161 5040 16227 5106 sw
tri 16161 4974 16227 5040 ne
tri 16227 4974 16293 5040 sw
tri 16227 4914 16287 4974 ne
rect 16287 4934 16293 4974
tri 16293 4934 16333 4974 sw
tri 16221 2975 16287 3041 se
rect 16287 3021 16333 4934
tri 16287 2975 16333 3021 nw
tri 16164 2918 16221 2975 se
rect 16221 2918 16230 2975
tri 16230 2918 16287 2975 nw
tri 15008 1850 15025 1867 ne
tri 14951 961 15025 1035 se
rect 15025 1013 15077 1867
tri 15077 1808 15136 1867 nw
tri 15134 1722 15185 1773 ne
tri 15025 961 15077 1013 nw
tri 15111 977 15185 1051 se
rect 15185 1029 15237 1773
tri 15237 1748 15262 1773 nw
tri 16158 1729 16164 1735 se
rect 16164 1729 16210 2918
tri 16210 2898 16230 2918 nw
tri 16445 2305 16479 2339 ne
rect 16479 1341 16531 2339
tri 15185 977 15237 1029 nw
tri 15095 961 15111 977 se
tri 14877 887 14951 961 se
rect 14951 903 14967 961
tri 14967 903 15025 961 nw
tri 15037 903 15095 961 se
rect 15095 903 15111 961
tri 15111 903 15185 977 nw
tri 14951 887 14967 903 nw
tri 14871 881 14877 887 se
rect 14877 881 14908 887
tri 14908 844 14951 887 nw
tri 15018 884 15037 903 se
rect 15037 884 15052 903
tri 15052 844 15111 903 nw
<< metal3 >>
tri 2121 14799 2151 14829 se
rect 2151 14801 2217 14990
rect 2151 14799 2215 14801
tri 2215 14799 2217 14801 nw
tri 2027 14705 2121 14799 se
tri 2121 14705 2215 14799 nw
tri 1933 14611 2027 14705 se
tri 2027 14611 2121 14705 nw
tri 1839 14517 1933 14611 se
tri 1933 14517 2027 14611 nw
tri 1773 14451 1839 14517 se
rect 1773 7114 1839 14451
tri 1839 14423 1933 14517 nw
tri 2907 10600 2922 10615 ne
tri 2851 7694 2922 7765 se
rect 2922 7694 2988 10615
tri 2988 10550 3053 10615 nw
tri 2988 7694 3007 7713 sw
tri 1773 7048 1839 7114 ne
tri 1839 7103 1878 7142 sw
rect 1839 7048 1878 7103
tri 1839 7009 1878 7048 ne
tri 1878 7009 1972 7103 sw
tri 1878 6915 1972 7009 ne
tri 1972 6915 2066 7009 sw
tri 1972 6821 2066 6915 ne
tri 2066 6821 2160 6915 sw
tri 2066 6727 2160 6821 ne
tri 2160 6727 2254 6821 sw
tri 2160 6633 2254 6727 ne
tri 2254 6633 2348 6727 sw
tri 2254 6605 2282 6633 ne
tri 2220 1227 2282 1289 se
rect 2282 1261 2348 6633
rect 2282 1227 2314 1261
tri 2314 1227 2348 1261 nw
rect 14510 2356 14996 2491
tri 14996 2356 15131 2491 sw
tri 1699 1133 1793 1227 se
rect 1793 1161 2248 1227
tri 2248 1161 2314 1227 nw
tri 1793 1133 1821 1161 nw
tri 1680 1114 1699 1133 se
rect 1699 1114 1746 1133
tri 1670 -363 1680 -353 se
rect 1680 -395 1746 1114
tri 1746 1086 1793 1133 nw
rect 14510 1111 15131 2356
tri 1746 -363 1826 -283 sw
use sky130_fd_io__gpiov2_amux_ctl_inv_1  sky130_fd_io__gpiov2_amux_ctl_inv_1_0
timestamp 1676037725
transform -1 0 14983 0 1 494
box 0 0 1 1
use sky130_fd_io__gpiov2_amux_ctl_inv_1  sky130_fd_io__gpiov2_amux_ctl_inv_1_1
timestamp 1676037725
transform -1 0 15292 0 1 494
box 0 0 1 1
use sky130_fd_io__gpiov2_amux_ctl_ls  sky130_fd_io__gpiov2_amux_ctl_ls_0
timestamp 1676037725
transform 1 0 14705 0 1 1344
box 53 163 2159 1426
use sky130_fd_io__gpiov2_amux_ctl_lshv2hv2  sky130_fd_io__gpiov2_amux_ctl_lshv2hv2_0
timestamp 1676037725
transform 1 0 748 0 1 13628
box 290 665 1808 3319
use sky130_fd_io__gpiov2_amux_ctl_lshv2hv  sky130_fd_io__gpiov2_amux_ctl_lshv2hv_0
timestamp 1676037725
transform -1 0 8787 0 1 10523
box 3564 882 6767 1429
use sky130_fd_io__tap_1  sky130_fd_io__tap_1_0
timestamp 1676037725
transform -1 0 14675 0 1 494
box -38 -49 134 715
use sky130_fd_pr__model__nfet_highvoltage__example_55959141808586  sky130_fd_pr__model__nfet_highvoltage__example_55959141808586_0
timestamp 1676037725
transform -1 0 1459 0 -1 11410
box -1 0 121 1
use sky130_fd_pr__model__pfet_highvoltage__example_55959141808421  sky130_fd_pr__model__pfet_highvoltage__example_55959141808421_0
timestamp 1676037725
transform 1 0 1286 0 -1 10835
box -1 0 297 1
<< properties >>
string GDS_END 43862376
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 43836720
<< end >>
