magic
tech sky130B
magscale 1 2
timestamp 1676037725
<< nwell >>
rect -38 261 866 582
<< pwell >>
rect 31 21 762 203
rect 31 17 63 21
rect 29 -17 63 17
<< scnmos >>
rect 119 47 149 177
rect 210 47 240 177
rect 294 47 324 177
rect 482 47 512 177
rect 566 47 596 177
rect 650 47 680 177
<< scpmoshvt >>
rect 119 297 149 497
rect 215 297 245 497
rect 287 297 317 497
rect 482 297 512 497
rect 554 297 584 497
rect 650 297 680 497
<< ndiff >>
rect 57 163 119 177
rect 57 129 65 163
rect 99 129 119 163
rect 57 95 119 129
rect 57 61 65 95
rect 99 61 119 95
rect 57 47 119 61
rect 149 95 210 177
rect 149 61 165 95
rect 199 61 210 95
rect 149 47 210 61
rect 240 163 294 177
rect 240 129 250 163
rect 284 129 294 163
rect 240 47 294 129
rect 324 95 376 177
rect 324 61 334 95
rect 368 61 376 95
rect 324 47 376 61
rect 430 95 482 177
rect 430 61 438 95
rect 472 61 482 95
rect 430 47 482 61
rect 512 163 566 177
rect 512 129 522 163
rect 556 129 566 163
rect 512 95 566 129
rect 512 61 522 95
rect 556 61 566 95
rect 512 47 566 61
rect 596 163 650 177
rect 596 129 606 163
rect 640 129 650 163
rect 596 95 650 129
rect 596 61 606 95
rect 640 61 650 95
rect 596 47 650 61
rect 680 163 736 177
rect 680 129 690 163
rect 724 129 736 163
rect 680 95 736 129
rect 680 61 690 95
rect 724 61 736 95
rect 680 47 736 61
<< pdiff >>
rect 51 477 119 497
rect 51 443 74 477
rect 108 443 119 477
rect 51 409 119 443
rect 51 375 74 409
rect 108 375 119 409
rect 51 341 119 375
rect 51 307 74 341
rect 108 307 119 341
rect 51 297 119 307
rect 149 477 215 497
rect 149 443 163 477
rect 197 443 215 477
rect 149 409 215 443
rect 149 375 163 409
rect 197 375 215 409
rect 149 297 215 375
rect 245 297 287 497
rect 317 477 482 497
rect 317 443 327 477
rect 361 443 438 477
rect 472 443 482 477
rect 317 409 482 443
rect 317 375 327 409
rect 361 375 438 409
rect 472 375 482 409
rect 317 297 482 375
rect 512 297 554 497
rect 584 477 650 497
rect 584 443 594 477
rect 628 443 650 477
rect 584 409 650 443
rect 584 375 594 409
rect 628 375 650 409
rect 584 297 650 375
rect 680 477 736 497
rect 680 443 694 477
rect 728 443 736 477
rect 680 409 736 443
rect 680 375 694 409
rect 728 375 736 409
rect 680 297 736 375
<< ndiffc >>
rect 65 129 99 163
rect 65 61 99 95
rect 165 61 199 95
rect 250 129 284 163
rect 334 61 368 95
rect 438 61 472 95
rect 522 129 556 163
rect 522 61 556 95
rect 606 129 640 163
rect 606 61 640 95
rect 690 129 724 163
rect 690 61 724 95
<< pdiffc >>
rect 74 443 108 477
rect 74 375 108 409
rect 74 307 108 341
rect 163 443 197 477
rect 163 375 197 409
rect 327 443 361 477
rect 438 443 472 477
rect 327 375 361 409
rect 438 375 472 409
rect 594 443 628 477
rect 594 375 628 409
rect 694 443 728 477
rect 694 375 728 409
<< poly >>
rect 119 497 149 523
rect 215 497 245 523
rect 287 497 317 523
rect 482 497 512 523
rect 554 497 584 523
rect 650 497 680 523
rect 119 265 149 297
rect 215 265 245 297
rect 23 249 149 265
rect 23 215 33 249
rect 67 215 149 249
rect 23 199 149 215
rect 191 249 245 265
rect 191 215 201 249
rect 235 215 245 249
rect 191 199 245 215
rect 287 265 317 297
rect 482 265 512 297
rect 287 249 357 265
rect 287 215 313 249
rect 347 215 357 249
rect 287 199 357 215
rect 438 249 512 265
rect 438 215 448 249
rect 482 215 512 249
rect 438 199 512 215
rect 554 265 584 297
rect 650 265 680 297
rect 554 249 608 265
rect 554 215 564 249
rect 598 215 608 249
rect 554 199 608 215
rect 650 249 721 265
rect 650 215 677 249
rect 711 215 721 249
rect 650 199 721 215
rect 119 177 149 199
rect 210 177 240 199
rect 294 177 324 199
rect 482 177 512 199
rect 566 177 596 199
rect 650 177 680 199
rect 119 21 149 47
rect 210 21 240 47
rect 294 21 324 47
rect 482 21 512 47
rect 566 21 596 47
rect 650 21 680 47
<< polycont >>
rect 33 215 67 249
rect 201 215 235 249
rect 313 215 347 249
rect 448 215 482 249
rect 564 215 598 249
rect 677 215 711 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 48 477 108 493
rect 48 443 74 477
rect 48 409 108 443
rect 48 375 74 409
rect 48 341 108 375
rect 147 477 197 527
rect 147 443 163 477
rect 147 409 197 443
rect 315 477 476 493
rect 315 443 327 477
rect 361 443 438 477
rect 472 443 476 477
rect 315 409 476 443
rect 578 477 644 527
rect 578 443 594 477
rect 628 443 644 477
rect 578 409 644 443
rect 147 375 163 409
rect 147 359 197 375
rect 231 375 327 409
rect 361 375 438 409
rect 472 375 544 409
rect 48 307 74 341
rect 231 325 265 375
rect 108 307 265 325
rect 48 291 265 307
rect 17 249 83 257
rect 17 215 33 249
rect 67 215 83 249
rect 17 199 83 215
rect 117 165 151 291
rect 299 265 363 341
rect 185 249 251 257
rect 185 215 201 249
rect 235 215 251 249
rect 287 249 363 265
rect 287 215 313 249
rect 347 215 363 249
rect 401 257 476 341
rect 510 325 544 375
rect 578 375 594 409
rect 628 375 644 409
rect 678 477 811 493
rect 678 443 694 477
rect 728 443 811 477
rect 678 409 811 443
rect 678 375 694 409
rect 728 375 811 409
rect 578 359 644 375
rect 510 291 694 325
rect 660 257 694 291
rect 401 249 498 257
rect 401 215 448 249
rect 482 215 498 249
rect 536 249 626 257
rect 536 215 564 249
rect 598 215 626 249
rect 660 249 727 257
rect 660 215 677 249
rect 711 215 727 249
rect 761 181 811 375
rect 49 163 151 165
rect 49 129 65 163
rect 99 129 151 163
rect 232 163 572 181
rect 232 129 250 163
rect 284 147 522 163
rect 284 129 309 147
rect 506 129 522 147
rect 556 129 572 163
rect 49 95 115 129
rect 438 95 472 111
rect 49 61 65 95
rect 99 61 115 95
rect 149 61 165 95
rect 199 61 334 95
rect 368 61 386 95
rect 49 51 115 61
rect 438 17 472 61
rect 506 95 572 129
rect 506 61 522 95
rect 556 61 572 95
rect 506 54 572 61
rect 606 163 640 181
rect 606 95 640 129
rect 606 17 640 61
rect 674 163 811 181
rect 674 129 690 163
rect 724 129 811 163
rect 674 95 811 129
rect 674 61 690 95
rect 724 61 811 95
rect 674 53 811 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
<< metal1 >>
rect 0 561 828 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 496 828 527
rect 0 17 828 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 -48 828 -17
<< labels >>
flabel locali s 401 221 435 255 0 FreeSans 400 0 0 0 A2
port 2 nsew signal input
flabel locali s 765 357 799 391 0 FreeSans 400 0 0 0 X
port 10 nsew signal output
flabel locali s 213 221 247 255 0 FreeSans 400 0 0 0 B1
port 3 nsew signal input
flabel locali s 29 221 63 255 0 FreeSans 400 0 0 0 C1
port 5 nsew signal input
flabel locali s 585 221 619 255 0 FreeSans 400 0 0 0 A1
port 1 nsew signal input
flabel locali s 401 289 435 323 0 FreeSans 400 0 0 0 A2
port 2 nsew signal input
flabel locali s 305 221 339 255 0 FreeSans 400 0 0 0 B2
port 4 nsew signal input
flabel locali s 305 289 339 323 0 FreeSans 400 0 0 0 B2
port 4 nsew signal input
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 6 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 9 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 o221a_1
rlabel metal1 s 0 -48 828 48 1 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 496 828 592 1 VPWR
port 9 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 828 544
string GDS_END 801168
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 793938
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 4.140 0.000 
<< end >>
