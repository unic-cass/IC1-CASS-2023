magic
tech sky130B
magscale 1 2
timestamp 1676037725
<< dnwell >>
rect 214 214 2578 2578
<< nwell >>
rect 134 2298 2658 2658
rect 134 494 494 2298
rect 2298 494 2658 2298
rect 134 134 2658 494
<< pwell >>
rect 0 2658 2792 2792
rect 0 134 134 2658
rect 628 628 2164 2164
rect 2658 134 2792 2658
rect 0 0 2792 134
<< ndiff >>
rect 896 1855 1896 1896
rect 896 937 937 1855
rect 1855 937 1896 1855
rect 896 896 1896 937
<< ndiffc >>
rect 937 937 1855 1855
<< psubdiff >>
rect 26 2742 2766 2766
rect 26 2708 50 2742
rect 84 2708 121 2742
rect 155 2708 189 2742
rect 223 2708 257 2742
rect 291 2708 325 2742
rect 359 2708 393 2742
rect 427 2708 461 2742
rect 495 2708 529 2742
rect 563 2708 597 2742
rect 631 2708 665 2742
rect 699 2708 733 2742
rect 767 2708 801 2742
rect 835 2708 869 2742
rect 903 2708 937 2742
rect 971 2708 1005 2742
rect 1039 2708 1073 2742
rect 1107 2708 1141 2742
rect 1175 2708 1209 2742
rect 1243 2708 1277 2742
rect 1311 2708 1345 2742
rect 1379 2708 1413 2742
rect 1447 2708 1481 2742
rect 1515 2708 1549 2742
rect 1583 2708 1617 2742
rect 1651 2708 1685 2742
rect 1719 2708 1753 2742
rect 1787 2708 1821 2742
rect 1855 2708 1889 2742
rect 1923 2708 1957 2742
rect 1991 2708 2025 2742
rect 2059 2708 2093 2742
rect 2127 2708 2161 2742
rect 2195 2708 2229 2742
rect 2263 2708 2297 2742
rect 2331 2708 2365 2742
rect 2399 2708 2433 2742
rect 2467 2708 2501 2742
rect 2535 2708 2569 2742
rect 2603 2708 2637 2742
rect 2671 2708 2708 2742
rect 2742 2708 2766 2742
rect 26 2684 2766 2708
rect 26 2671 108 2684
rect 26 2637 50 2671
rect 84 2637 108 2671
rect 26 2603 108 2637
rect 26 2569 50 2603
rect 84 2569 108 2603
rect 26 2535 108 2569
rect 2684 2671 2766 2684
rect 2684 2637 2708 2671
rect 2742 2637 2766 2671
rect 2684 2603 2766 2637
rect 2684 2569 2708 2603
rect 2742 2569 2766 2603
rect 26 2501 50 2535
rect 84 2501 108 2535
rect 26 2467 108 2501
rect 26 2433 50 2467
rect 84 2433 108 2467
rect 26 2399 108 2433
rect 26 2365 50 2399
rect 84 2365 108 2399
rect 26 2331 108 2365
rect 26 2297 50 2331
rect 84 2297 108 2331
rect 26 2263 108 2297
rect 26 2229 50 2263
rect 84 2229 108 2263
rect 26 2195 108 2229
rect 26 2161 50 2195
rect 84 2161 108 2195
rect 26 2127 108 2161
rect 26 2093 50 2127
rect 84 2093 108 2127
rect 26 2059 108 2093
rect 26 2025 50 2059
rect 84 2025 108 2059
rect 26 1991 108 2025
rect 26 1957 50 1991
rect 84 1957 108 1991
rect 26 1923 108 1957
rect 26 1889 50 1923
rect 84 1889 108 1923
rect 26 1855 108 1889
rect 26 1821 50 1855
rect 84 1821 108 1855
rect 26 1787 108 1821
rect 26 1753 50 1787
rect 84 1753 108 1787
rect 26 1719 108 1753
rect 26 1685 50 1719
rect 84 1685 108 1719
rect 26 1651 108 1685
rect 26 1617 50 1651
rect 84 1617 108 1651
rect 26 1583 108 1617
rect 26 1549 50 1583
rect 84 1549 108 1583
rect 26 1515 108 1549
rect 26 1481 50 1515
rect 84 1481 108 1515
rect 26 1447 108 1481
rect 26 1413 50 1447
rect 84 1413 108 1447
rect 26 1379 108 1413
rect 26 1345 50 1379
rect 84 1345 108 1379
rect 26 1311 108 1345
rect 26 1277 50 1311
rect 84 1277 108 1311
rect 26 1243 108 1277
rect 26 1209 50 1243
rect 84 1209 108 1243
rect 26 1175 108 1209
rect 26 1141 50 1175
rect 84 1141 108 1175
rect 26 1107 108 1141
rect 26 1073 50 1107
rect 84 1073 108 1107
rect 26 1039 108 1073
rect 26 1005 50 1039
rect 84 1005 108 1039
rect 26 971 108 1005
rect 26 937 50 971
rect 84 937 108 971
rect 26 903 108 937
rect 26 869 50 903
rect 84 869 108 903
rect 26 835 108 869
rect 26 801 50 835
rect 84 801 108 835
rect 26 767 108 801
rect 26 733 50 767
rect 84 733 108 767
rect 26 699 108 733
rect 26 665 50 699
rect 84 665 108 699
rect 26 631 108 665
rect 26 597 50 631
rect 84 597 108 631
rect 26 563 108 597
rect 26 529 50 563
rect 84 529 108 563
rect 26 495 108 529
rect 26 461 50 495
rect 84 461 108 495
rect 26 427 108 461
rect 26 393 50 427
rect 84 393 108 427
rect 26 359 108 393
rect 26 325 50 359
rect 84 325 108 359
rect 26 291 108 325
rect 26 257 50 291
rect 84 257 108 291
rect 26 223 108 257
rect 654 2114 2138 2138
rect 654 2080 678 2114
rect 712 2080 767 2114
rect 801 2080 835 2114
rect 869 2080 903 2114
rect 937 2080 971 2114
rect 1005 2080 1039 2114
rect 1073 2080 1107 2114
rect 1141 2080 1175 2114
rect 1209 2080 1243 2114
rect 1277 2080 1311 2114
rect 1345 2080 1379 2114
rect 1413 2080 1447 2114
rect 1481 2080 1515 2114
rect 1549 2080 1583 2114
rect 1617 2080 1651 2114
rect 1685 2080 1719 2114
rect 1753 2080 1787 2114
rect 1821 2080 1855 2114
rect 1889 2080 1923 2114
rect 1957 2080 1991 2114
rect 2025 2080 2080 2114
rect 2114 2080 2138 2114
rect 654 2056 2138 2080
rect 654 2025 736 2056
rect 654 1991 678 2025
rect 712 1991 736 2025
rect 654 1957 736 1991
rect 654 1923 678 1957
rect 712 1923 736 1957
rect 654 1889 736 1923
rect 2056 2025 2138 2056
rect 2056 1991 2080 2025
rect 2114 1991 2138 2025
rect 2056 1957 2138 1991
rect 2056 1923 2080 1957
rect 2114 1923 2138 1957
rect 654 1855 678 1889
rect 712 1855 736 1889
rect 654 1821 736 1855
rect 654 1787 678 1821
rect 712 1787 736 1821
rect 654 1753 736 1787
rect 654 1719 678 1753
rect 712 1719 736 1753
rect 654 1685 736 1719
rect 654 1651 678 1685
rect 712 1651 736 1685
rect 654 1617 736 1651
rect 654 1583 678 1617
rect 712 1583 736 1617
rect 654 1549 736 1583
rect 654 1515 678 1549
rect 712 1515 736 1549
rect 654 1481 736 1515
rect 654 1447 678 1481
rect 712 1447 736 1481
rect 654 1413 736 1447
rect 654 1379 678 1413
rect 712 1379 736 1413
rect 654 1345 736 1379
rect 654 1311 678 1345
rect 712 1311 736 1345
rect 654 1277 736 1311
rect 654 1243 678 1277
rect 712 1243 736 1277
rect 654 1209 736 1243
rect 654 1175 678 1209
rect 712 1175 736 1209
rect 654 1141 736 1175
rect 654 1107 678 1141
rect 712 1107 736 1141
rect 654 1073 736 1107
rect 654 1039 678 1073
rect 712 1039 736 1073
rect 654 1005 736 1039
rect 654 971 678 1005
rect 712 971 736 1005
rect 654 937 736 971
rect 654 903 678 937
rect 712 903 736 937
rect 654 869 736 903
rect 2056 1889 2138 1923
rect 2056 1855 2080 1889
rect 2114 1855 2138 1889
rect 2056 1821 2138 1855
rect 2056 1787 2080 1821
rect 2114 1787 2138 1821
rect 2056 1753 2138 1787
rect 2056 1719 2080 1753
rect 2114 1719 2138 1753
rect 2056 1685 2138 1719
rect 2056 1651 2080 1685
rect 2114 1651 2138 1685
rect 2056 1617 2138 1651
rect 2056 1583 2080 1617
rect 2114 1583 2138 1617
rect 2056 1549 2138 1583
rect 2056 1515 2080 1549
rect 2114 1515 2138 1549
rect 2056 1481 2138 1515
rect 2056 1447 2080 1481
rect 2114 1447 2138 1481
rect 2056 1413 2138 1447
rect 2056 1379 2080 1413
rect 2114 1379 2138 1413
rect 2056 1345 2138 1379
rect 2056 1311 2080 1345
rect 2114 1311 2138 1345
rect 2056 1277 2138 1311
rect 2056 1243 2080 1277
rect 2114 1243 2138 1277
rect 2056 1209 2138 1243
rect 2056 1175 2080 1209
rect 2114 1175 2138 1209
rect 2056 1141 2138 1175
rect 2056 1107 2080 1141
rect 2114 1107 2138 1141
rect 2056 1073 2138 1107
rect 2056 1039 2080 1073
rect 2114 1039 2138 1073
rect 2056 1005 2138 1039
rect 2056 971 2080 1005
rect 2114 971 2138 1005
rect 2056 937 2138 971
rect 2056 903 2080 937
rect 2114 903 2138 937
rect 654 835 678 869
rect 712 835 736 869
rect 654 801 736 835
rect 654 767 678 801
rect 712 767 736 801
rect 654 736 736 767
rect 2056 869 2138 903
rect 2056 835 2080 869
rect 2114 835 2138 869
rect 2056 801 2138 835
rect 2056 767 2080 801
rect 2114 767 2138 801
rect 2056 736 2138 767
rect 654 712 2138 736
rect 654 678 678 712
rect 712 678 767 712
rect 801 678 835 712
rect 869 678 903 712
rect 937 678 971 712
rect 1005 678 1039 712
rect 1073 678 1107 712
rect 1141 678 1175 712
rect 1209 678 1243 712
rect 1277 678 1311 712
rect 1345 678 1379 712
rect 1413 678 1447 712
rect 1481 678 1515 712
rect 1549 678 1583 712
rect 1617 678 1651 712
rect 1685 678 1719 712
rect 1753 678 1787 712
rect 1821 678 1855 712
rect 1889 678 1923 712
rect 1957 678 1991 712
rect 2025 678 2080 712
rect 2114 678 2138 712
rect 654 654 2138 678
rect 2684 2535 2766 2569
rect 2684 2501 2708 2535
rect 2742 2501 2766 2535
rect 2684 2467 2766 2501
rect 2684 2433 2708 2467
rect 2742 2433 2766 2467
rect 2684 2399 2766 2433
rect 2684 2365 2708 2399
rect 2742 2365 2766 2399
rect 2684 2331 2766 2365
rect 2684 2297 2708 2331
rect 2742 2297 2766 2331
rect 2684 2263 2766 2297
rect 2684 2229 2708 2263
rect 2742 2229 2766 2263
rect 2684 2195 2766 2229
rect 2684 2161 2708 2195
rect 2742 2161 2766 2195
rect 2684 2127 2766 2161
rect 2684 2093 2708 2127
rect 2742 2093 2766 2127
rect 2684 2059 2766 2093
rect 2684 2025 2708 2059
rect 2742 2025 2766 2059
rect 2684 1991 2766 2025
rect 2684 1957 2708 1991
rect 2742 1957 2766 1991
rect 2684 1923 2766 1957
rect 2684 1889 2708 1923
rect 2742 1889 2766 1923
rect 2684 1855 2766 1889
rect 2684 1821 2708 1855
rect 2742 1821 2766 1855
rect 2684 1787 2766 1821
rect 2684 1753 2708 1787
rect 2742 1753 2766 1787
rect 2684 1719 2766 1753
rect 2684 1685 2708 1719
rect 2742 1685 2766 1719
rect 2684 1651 2766 1685
rect 2684 1617 2708 1651
rect 2742 1617 2766 1651
rect 2684 1583 2766 1617
rect 2684 1549 2708 1583
rect 2742 1549 2766 1583
rect 2684 1515 2766 1549
rect 2684 1481 2708 1515
rect 2742 1481 2766 1515
rect 2684 1447 2766 1481
rect 2684 1413 2708 1447
rect 2742 1413 2766 1447
rect 2684 1379 2766 1413
rect 2684 1345 2708 1379
rect 2742 1345 2766 1379
rect 2684 1311 2766 1345
rect 2684 1277 2708 1311
rect 2742 1277 2766 1311
rect 2684 1243 2766 1277
rect 2684 1209 2708 1243
rect 2742 1209 2766 1243
rect 2684 1175 2766 1209
rect 2684 1141 2708 1175
rect 2742 1141 2766 1175
rect 2684 1107 2766 1141
rect 2684 1073 2708 1107
rect 2742 1073 2766 1107
rect 2684 1039 2766 1073
rect 2684 1005 2708 1039
rect 2742 1005 2766 1039
rect 2684 971 2766 1005
rect 2684 937 2708 971
rect 2742 937 2766 971
rect 2684 903 2766 937
rect 2684 869 2708 903
rect 2742 869 2766 903
rect 2684 835 2766 869
rect 2684 801 2708 835
rect 2742 801 2766 835
rect 2684 767 2766 801
rect 2684 733 2708 767
rect 2742 733 2766 767
rect 2684 699 2766 733
rect 2684 665 2708 699
rect 2742 665 2766 699
rect 2684 631 2766 665
rect 2684 597 2708 631
rect 2742 597 2766 631
rect 2684 563 2766 597
rect 2684 529 2708 563
rect 2742 529 2766 563
rect 2684 495 2766 529
rect 2684 461 2708 495
rect 2742 461 2766 495
rect 2684 427 2766 461
rect 2684 393 2708 427
rect 2742 393 2766 427
rect 2684 359 2766 393
rect 2684 325 2708 359
rect 2742 325 2766 359
rect 2684 291 2766 325
rect 2684 257 2708 291
rect 2742 257 2766 291
rect 26 189 50 223
rect 84 189 108 223
rect 26 155 108 189
rect 26 121 50 155
rect 84 121 108 155
rect 26 108 108 121
rect 2684 223 2766 257
rect 2684 189 2708 223
rect 2742 189 2766 223
rect 2684 155 2766 189
rect 2684 121 2708 155
rect 2742 121 2766 155
rect 2684 108 2766 121
rect 26 84 2766 108
rect 26 50 50 84
rect 84 50 121 84
rect 155 50 189 84
rect 223 50 257 84
rect 291 50 325 84
rect 359 50 393 84
rect 427 50 461 84
rect 495 50 529 84
rect 563 50 597 84
rect 631 50 665 84
rect 699 50 733 84
rect 767 50 801 84
rect 835 50 869 84
rect 903 50 937 84
rect 971 50 1005 84
rect 1039 50 1073 84
rect 1107 50 1141 84
rect 1175 50 1209 84
rect 1243 50 1277 84
rect 1311 50 1345 84
rect 1379 50 1413 84
rect 1447 50 1481 84
rect 1515 50 1549 84
rect 1583 50 1617 84
rect 1651 50 1685 84
rect 1719 50 1753 84
rect 1787 50 1821 84
rect 1855 50 1889 84
rect 1923 50 1957 84
rect 1991 50 2025 84
rect 2059 50 2093 84
rect 2127 50 2161 84
rect 2195 50 2229 84
rect 2263 50 2297 84
rect 2331 50 2365 84
rect 2399 50 2433 84
rect 2467 50 2501 84
rect 2535 50 2569 84
rect 2603 50 2637 84
rect 2671 50 2708 84
rect 2742 50 2766 84
rect 26 26 2766 50
<< nsubdiff >>
rect 252 2516 2540 2540
rect 252 2482 276 2516
rect 310 2482 359 2516
rect 393 2482 427 2516
rect 461 2482 495 2516
rect 529 2482 563 2516
rect 597 2482 631 2516
rect 665 2482 699 2516
rect 733 2482 767 2516
rect 801 2482 835 2516
rect 869 2482 903 2516
rect 937 2482 971 2516
rect 1005 2482 1039 2516
rect 1073 2482 1107 2516
rect 1141 2482 1175 2516
rect 1209 2482 1243 2516
rect 1277 2482 1311 2516
rect 1345 2482 1379 2516
rect 1413 2482 1447 2516
rect 1481 2482 1515 2516
rect 1549 2482 1583 2516
rect 1617 2482 1651 2516
rect 1685 2482 1719 2516
rect 1753 2482 1787 2516
rect 1821 2482 1855 2516
rect 1889 2482 1923 2516
rect 1957 2482 1991 2516
rect 2025 2482 2059 2516
rect 2093 2482 2127 2516
rect 2161 2482 2195 2516
rect 2229 2482 2263 2516
rect 2297 2482 2331 2516
rect 2365 2482 2399 2516
rect 2433 2482 2482 2516
rect 2516 2482 2540 2516
rect 252 2458 2540 2482
rect 252 2433 334 2458
rect 252 2399 276 2433
rect 310 2399 334 2433
rect 252 2365 334 2399
rect 252 2331 276 2365
rect 310 2331 334 2365
rect 252 2297 334 2331
rect 252 2263 276 2297
rect 310 2263 334 2297
rect 252 2229 334 2263
rect 252 2195 276 2229
rect 310 2195 334 2229
rect 252 2161 334 2195
rect 252 2127 276 2161
rect 310 2127 334 2161
rect 2458 2433 2540 2458
rect 2458 2399 2482 2433
rect 2516 2399 2540 2433
rect 2458 2365 2540 2399
rect 2458 2331 2482 2365
rect 2516 2331 2540 2365
rect 2458 2297 2540 2331
rect 2458 2263 2482 2297
rect 2516 2263 2540 2297
rect 2458 2229 2540 2263
rect 2458 2195 2482 2229
rect 2516 2195 2540 2229
rect 2458 2161 2540 2195
rect 252 2093 334 2127
rect 252 2059 276 2093
rect 310 2059 334 2093
rect 252 2025 334 2059
rect 252 1991 276 2025
rect 310 1991 334 2025
rect 252 1957 334 1991
rect 252 1923 276 1957
rect 310 1923 334 1957
rect 252 1889 334 1923
rect 252 1855 276 1889
rect 310 1855 334 1889
rect 252 1821 334 1855
rect 252 1787 276 1821
rect 310 1787 334 1821
rect 252 1753 334 1787
rect 252 1719 276 1753
rect 310 1719 334 1753
rect 252 1685 334 1719
rect 252 1651 276 1685
rect 310 1651 334 1685
rect 252 1617 334 1651
rect 252 1583 276 1617
rect 310 1583 334 1617
rect 252 1549 334 1583
rect 252 1515 276 1549
rect 310 1515 334 1549
rect 252 1481 334 1515
rect 252 1447 276 1481
rect 310 1447 334 1481
rect 252 1413 334 1447
rect 252 1379 276 1413
rect 310 1379 334 1413
rect 252 1345 334 1379
rect 252 1311 276 1345
rect 310 1311 334 1345
rect 252 1277 334 1311
rect 252 1243 276 1277
rect 310 1243 334 1277
rect 252 1209 334 1243
rect 252 1175 276 1209
rect 310 1175 334 1209
rect 252 1141 334 1175
rect 252 1107 276 1141
rect 310 1107 334 1141
rect 252 1073 334 1107
rect 252 1039 276 1073
rect 310 1039 334 1073
rect 252 1005 334 1039
rect 252 971 276 1005
rect 310 971 334 1005
rect 252 937 334 971
rect 252 903 276 937
rect 310 903 334 937
rect 252 869 334 903
rect 252 835 276 869
rect 310 835 334 869
rect 252 801 334 835
rect 252 767 276 801
rect 310 767 334 801
rect 252 733 334 767
rect 252 699 276 733
rect 310 699 334 733
rect 252 665 334 699
rect 252 631 276 665
rect 310 631 334 665
rect 2458 2127 2482 2161
rect 2516 2127 2540 2161
rect 2458 2093 2540 2127
rect 2458 2059 2482 2093
rect 2516 2059 2540 2093
rect 2458 2025 2540 2059
rect 2458 1991 2482 2025
rect 2516 1991 2540 2025
rect 2458 1957 2540 1991
rect 2458 1923 2482 1957
rect 2516 1923 2540 1957
rect 2458 1889 2540 1923
rect 2458 1855 2482 1889
rect 2516 1855 2540 1889
rect 2458 1821 2540 1855
rect 2458 1787 2482 1821
rect 2516 1787 2540 1821
rect 2458 1753 2540 1787
rect 2458 1719 2482 1753
rect 2516 1719 2540 1753
rect 2458 1685 2540 1719
rect 2458 1651 2482 1685
rect 2516 1651 2540 1685
rect 2458 1617 2540 1651
rect 2458 1583 2482 1617
rect 2516 1583 2540 1617
rect 2458 1549 2540 1583
rect 2458 1515 2482 1549
rect 2516 1515 2540 1549
rect 2458 1481 2540 1515
rect 2458 1447 2482 1481
rect 2516 1447 2540 1481
rect 2458 1413 2540 1447
rect 2458 1379 2482 1413
rect 2516 1379 2540 1413
rect 2458 1345 2540 1379
rect 2458 1311 2482 1345
rect 2516 1311 2540 1345
rect 2458 1277 2540 1311
rect 2458 1243 2482 1277
rect 2516 1243 2540 1277
rect 2458 1209 2540 1243
rect 2458 1175 2482 1209
rect 2516 1175 2540 1209
rect 2458 1141 2540 1175
rect 2458 1107 2482 1141
rect 2516 1107 2540 1141
rect 2458 1073 2540 1107
rect 2458 1039 2482 1073
rect 2516 1039 2540 1073
rect 2458 1005 2540 1039
rect 2458 971 2482 1005
rect 2516 971 2540 1005
rect 2458 937 2540 971
rect 2458 903 2482 937
rect 2516 903 2540 937
rect 2458 869 2540 903
rect 2458 835 2482 869
rect 2516 835 2540 869
rect 2458 801 2540 835
rect 2458 767 2482 801
rect 2516 767 2540 801
rect 2458 733 2540 767
rect 2458 699 2482 733
rect 2516 699 2540 733
rect 2458 665 2540 699
rect 252 597 334 631
rect 252 563 276 597
rect 310 563 334 597
rect 252 529 334 563
rect 252 495 276 529
rect 310 495 334 529
rect 252 461 334 495
rect 252 427 276 461
rect 310 427 334 461
rect 252 393 334 427
rect 252 359 276 393
rect 310 359 334 393
rect 252 334 334 359
rect 2458 631 2482 665
rect 2516 631 2540 665
rect 2458 597 2540 631
rect 2458 563 2482 597
rect 2516 563 2540 597
rect 2458 529 2540 563
rect 2458 495 2482 529
rect 2516 495 2540 529
rect 2458 461 2540 495
rect 2458 427 2482 461
rect 2516 427 2540 461
rect 2458 393 2540 427
rect 2458 359 2482 393
rect 2516 359 2540 393
rect 2458 334 2540 359
rect 252 310 2540 334
rect 252 276 276 310
rect 310 276 359 310
rect 393 276 427 310
rect 461 276 495 310
rect 529 276 563 310
rect 597 276 631 310
rect 665 276 699 310
rect 733 276 767 310
rect 801 276 835 310
rect 869 276 903 310
rect 937 276 971 310
rect 1005 276 1039 310
rect 1073 276 1107 310
rect 1141 276 1175 310
rect 1209 276 1243 310
rect 1277 276 1311 310
rect 1345 276 1379 310
rect 1413 276 1447 310
rect 1481 276 1515 310
rect 1549 276 1583 310
rect 1617 276 1651 310
rect 1685 276 1719 310
rect 1753 276 1787 310
rect 1821 276 1855 310
rect 1889 276 1923 310
rect 1957 276 1991 310
rect 2025 276 2059 310
rect 2093 276 2127 310
rect 2161 276 2195 310
rect 2229 276 2263 310
rect 2297 276 2331 310
rect 2365 276 2399 310
rect 2433 276 2482 310
rect 2516 276 2540 310
rect 252 252 2540 276
<< psubdiffcont >>
rect 50 2708 84 2742
rect 121 2708 155 2742
rect 189 2708 223 2742
rect 257 2708 291 2742
rect 325 2708 359 2742
rect 393 2708 427 2742
rect 461 2708 495 2742
rect 529 2708 563 2742
rect 597 2708 631 2742
rect 665 2708 699 2742
rect 733 2708 767 2742
rect 801 2708 835 2742
rect 869 2708 903 2742
rect 937 2708 971 2742
rect 1005 2708 1039 2742
rect 1073 2708 1107 2742
rect 1141 2708 1175 2742
rect 1209 2708 1243 2742
rect 1277 2708 1311 2742
rect 1345 2708 1379 2742
rect 1413 2708 1447 2742
rect 1481 2708 1515 2742
rect 1549 2708 1583 2742
rect 1617 2708 1651 2742
rect 1685 2708 1719 2742
rect 1753 2708 1787 2742
rect 1821 2708 1855 2742
rect 1889 2708 1923 2742
rect 1957 2708 1991 2742
rect 2025 2708 2059 2742
rect 2093 2708 2127 2742
rect 2161 2708 2195 2742
rect 2229 2708 2263 2742
rect 2297 2708 2331 2742
rect 2365 2708 2399 2742
rect 2433 2708 2467 2742
rect 2501 2708 2535 2742
rect 2569 2708 2603 2742
rect 2637 2708 2671 2742
rect 2708 2708 2742 2742
rect 50 2637 84 2671
rect 50 2569 84 2603
rect 2708 2637 2742 2671
rect 2708 2569 2742 2603
rect 50 2501 84 2535
rect 50 2433 84 2467
rect 50 2365 84 2399
rect 50 2297 84 2331
rect 50 2229 84 2263
rect 50 2161 84 2195
rect 50 2093 84 2127
rect 50 2025 84 2059
rect 50 1957 84 1991
rect 50 1889 84 1923
rect 50 1821 84 1855
rect 50 1753 84 1787
rect 50 1685 84 1719
rect 50 1617 84 1651
rect 50 1549 84 1583
rect 50 1481 84 1515
rect 50 1413 84 1447
rect 50 1345 84 1379
rect 50 1277 84 1311
rect 50 1209 84 1243
rect 50 1141 84 1175
rect 50 1073 84 1107
rect 50 1005 84 1039
rect 50 937 84 971
rect 50 869 84 903
rect 50 801 84 835
rect 50 733 84 767
rect 50 665 84 699
rect 50 597 84 631
rect 50 529 84 563
rect 50 461 84 495
rect 50 393 84 427
rect 50 325 84 359
rect 50 257 84 291
rect 678 2080 712 2114
rect 767 2080 801 2114
rect 835 2080 869 2114
rect 903 2080 937 2114
rect 971 2080 1005 2114
rect 1039 2080 1073 2114
rect 1107 2080 1141 2114
rect 1175 2080 1209 2114
rect 1243 2080 1277 2114
rect 1311 2080 1345 2114
rect 1379 2080 1413 2114
rect 1447 2080 1481 2114
rect 1515 2080 1549 2114
rect 1583 2080 1617 2114
rect 1651 2080 1685 2114
rect 1719 2080 1753 2114
rect 1787 2080 1821 2114
rect 1855 2080 1889 2114
rect 1923 2080 1957 2114
rect 1991 2080 2025 2114
rect 2080 2080 2114 2114
rect 678 1991 712 2025
rect 678 1923 712 1957
rect 2080 1991 2114 2025
rect 2080 1923 2114 1957
rect 678 1855 712 1889
rect 678 1787 712 1821
rect 678 1719 712 1753
rect 678 1651 712 1685
rect 678 1583 712 1617
rect 678 1515 712 1549
rect 678 1447 712 1481
rect 678 1379 712 1413
rect 678 1311 712 1345
rect 678 1243 712 1277
rect 678 1175 712 1209
rect 678 1107 712 1141
rect 678 1039 712 1073
rect 678 971 712 1005
rect 678 903 712 937
rect 2080 1855 2114 1889
rect 2080 1787 2114 1821
rect 2080 1719 2114 1753
rect 2080 1651 2114 1685
rect 2080 1583 2114 1617
rect 2080 1515 2114 1549
rect 2080 1447 2114 1481
rect 2080 1379 2114 1413
rect 2080 1311 2114 1345
rect 2080 1243 2114 1277
rect 2080 1175 2114 1209
rect 2080 1107 2114 1141
rect 2080 1039 2114 1073
rect 2080 971 2114 1005
rect 2080 903 2114 937
rect 678 835 712 869
rect 678 767 712 801
rect 2080 835 2114 869
rect 2080 767 2114 801
rect 678 678 712 712
rect 767 678 801 712
rect 835 678 869 712
rect 903 678 937 712
rect 971 678 1005 712
rect 1039 678 1073 712
rect 1107 678 1141 712
rect 1175 678 1209 712
rect 1243 678 1277 712
rect 1311 678 1345 712
rect 1379 678 1413 712
rect 1447 678 1481 712
rect 1515 678 1549 712
rect 1583 678 1617 712
rect 1651 678 1685 712
rect 1719 678 1753 712
rect 1787 678 1821 712
rect 1855 678 1889 712
rect 1923 678 1957 712
rect 1991 678 2025 712
rect 2080 678 2114 712
rect 2708 2501 2742 2535
rect 2708 2433 2742 2467
rect 2708 2365 2742 2399
rect 2708 2297 2742 2331
rect 2708 2229 2742 2263
rect 2708 2161 2742 2195
rect 2708 2093 2742 2127
rect 2708 2025 2742 2059
rect 2708 1957 2742 1991
rect 2708 1889 2742 1923
rect 2708 1821 2742 1855
rect 2708 1753 2742 1787
rect 2708 1685 2742 1719
rect 2708 1617 2742 1651
rect 2708 1549 2742 1583
rect 2708 1481 2742 1515
rect 2708 1413 2742 1447
rect 2708 1345 2742 1379
rect 2708 1277 2742 1311
rect 2708 1209 2742 1243
rect 2708 1141 2742 1175
rect 2708 1073 2742 1107
rect 2708 1005 2742 1039
rect 2708 937 2742 971
rect 2708 869 2742 903
rect 2708 801 2742 835
rect 2708 733 2742 767
rect 2708 665 2742 699
rect 2708 597 2742 631
rect 2708 529 2742 563
rect 2708 461 2742 495
rect 2708 393 2742 427
rect 2708 325 2742 359
rect 2708 257 2742 291
rect 50 189 84 223
rect 50 121 84 155
rect 2708 189 2742 223
rect 2708 121 2742 155
rect 50 50 84 84
rect 121 50 155 84
rect 189 50 223 84
rect 257 50 291 84
rect 325 50 359 84
rect 393 50 427 84
rect 461 50 495 84
rect 529 50 563 84
rect 597 50 631 84
rect 665 50 699 84
rect 733 50 767 84
rect 801 50 835 84
rect 869 50 903 84
rect 937 50 971 84
rect 1005 50 1039 84
rect 1073 50 1107 84
rect 1141 50 1175 84
rect 1209 50 1243 84
rect 1277 50 1311 84
rect 1345 50 1379 84
rect 1413 50 1447 84
rect 1481 50 1515 84
rect 1549 50 1583 84
rect 1617 50 1651 84
rect 1685 50 1719 84
rect 1753 50 1787 84
rect 1821 50 1855 84
rect 1889 50 1923 84
rect 1957 50 1991 84
rect 2025 50 2059 84
rect 2093 50 2127 84
rect 2161 50 2195 84
rect 2229 50 2263 84
rect 2297 50 2331 84
rect 2365 50 2399 84
rect 2433 50 2467 84
rect 2501 50 2535 84
rect 2569 50 2603 84
rect 2637 50 2671 84
rect 2708 50 2742 84
<< nsubdiffcont >>
rect 276 2482 310 2516
rect 359 2482 393 2516
rect 427 2482 461 2516
rect 495 2482 529 2516
rect 563 2482 597 2516
rect 631 2482 665 2516
rect 699 2482 733 2516
rect 767 2482 801 2516
rect 835 2482 869 2516
rect 903 2482 937 2516
rect 971 2482 1005 2516
rect 1039 2482 1073 2516
rect 1107 2482 1141 2516
rect 1175 2482 1209 2516
rect 1243 2482 1277 2516
rect 1311 2482 1345 2516
rect 1379 2482 1413 2516
rect 1447 2482 1481 2516
rect 1515 2482 1549 2516
rect 1583 2482 1617 2516
rect 1651 2482 1685 2516
rect 1719 2482 1753 2516
rect 1787 2482 1821 2516
rect 1855 2482 1889 2516
rect 1923 2482 1957 2516
rect 1991 2482 2025 2516
rect 2059 2482 2093 2516
rect 2127 2482 2161 2516
rect 2195 2482 2229 2516
rect 2263 2482 2297 2516
rect 2331 2482 2365 2516
rect 2399 2482 2433 2516
rect 2482 2482 2516 2516
rect 276 2399 310 2433
rect 276 2331 310 2365
rect 276 2263 310 2297
rect 276 2195 310 2229
rect 276 2127 310 2161
rect 2482 2399 2516 2433
rect 2482 2331 2516 2365
rect 2482 2263 2516 2297
rect 2482 2195 2516 2229
rect 276 2059 310 2093
rect 276 1991 310 2025
rect 276 1923 310 1957
rect 276 1855 310 1889
rect 276 1787 310 1821
rect 276 1719 310 1753
rect 276 1651 310 1685
rect 276 1583 310 1617
rect 276 1515 310 1549
rect 276 1447 310 1481
rect 276 1379 310 1413
rect 276 1311 310 1345
rect 276 1243 310 1277
rect 276 1175 310 1209
rect 276 1107 310 1141
rect 276 1039 310 1073
rect 276 971 310 1005
rect 276 903 310 937
rect 276 835 310 869
rect 276 767 310 801
rect 276 699 310 733
rect 276 631 310 665
rect 2482 2127 2516 2161
rect 2482 2059 2516 2093
rect 2482 1991 2516 2025
rect 2482 1923 2516 1957
rect 2482 1855 2516 1889
rect 2482 1787 2516 1821
rect 2482 1719 2516 1753
rect 2482 1651 2516 1685
rect 2482 1583 2516 1617
rect 2482 1515 2516 1549
rect 2482 1447 2516 1481
rect 2482 1379 2516 1413
rect 2482 1311 2516 1345
rect 2482 1243 2516 1277
rect 2482 1175 2516 1209
rect 2482 1107 2516 1141
rect 2482 1039 2516 1073
rect 2482 971 2516 1005
rect 2482 903 2516 937
rect 2482 835 2516 869
rect 2482 767 2516 801
rect 2482 699 2516 733
rect 276 563 310 597
rect 276 495 310 529
rect 276 427 310 461
rect 276 359 310 393
rect 2482 631 2516 665
rect 2482 563 2516 597
rect 2482 495 2516 529
rect 2482 427 2516 461
rect 2482 359 2516 393
rect 276 276 310 310
rect 359 276 393 310
rect 427 276 461 310
rect 495 276 529 310
rect 563 276 597 310
rect 631 276 665 310
rect 699 276 733 310
rect 767 276 801 310
rect 835 276 869 310
rect 903 276 937 310
rect 971 276 1005 310
rect 1039 276 1073 310
rect 1107 276 1141 310
rect 1175 276 1209 310
rect 1243 276 1277 310
rect 1311 276 1345 310
rect 1379 276 1413 310
rect 1447 276 1481 310
rect 1515 276 1549 310
rect 1583 276 1617 310
rect 1651 276 1685 310
rect 1719 276 1753 310
rect 1787 276 1821 310
rect 1855 276 1889 310
rect 1923 276 1957 310
rect 1991 276 2025 310
rect 2059 276 2093 310
rect 2127 276 2161 310
rect 2195 276 2229 310
rect 2263 276 2297 310
rect 2331 276 2365 310
rect 2399 276 2433 310
rect 2482 276 2516 310
<< locali >>
rect 34 2742 2758 2758
rect 34 2708 50 2742
rect 84 2708 121 2742
rect 223 2708 227 2742
rect 291 2708 299 2742
rect 359 2708 371 2742
rect 427 2708 443 2742
rect 495 2708 515 2742
rect 563 2708 587 2742
rect 631 2708 659 2742
rect 699 2708 731 2742
rect 767 2708 801 2742
rect 837 2708 869 2742
rect 909 2708 937 2742
rect 981 2708 1005 2742
rect 1053 2708 1073 2742
rect 1125 2708 1141 2742
rect 1197 2708 1209 2742
rect 1269 2708 1277 2742
rect 1341 2708 1345 2742
rect 1447 2708 1451 2742
rect 1515 2708 1523 2742
rect 1583 2708 1595 2742
rect 1651 2708 1667 2742
rect 1719 2708 1739 2742
rect 1787 2708 1811 2742
rect 1855 2708 1883 2742
rect 1923 2708 1955 2742
rect 1991 2708 2025 2742
rect 2061 2708 2093 2742
rect 2133 2708 2161 2742
rect 2205 2708 2229 2742
rect 2277 2708 2297 2742
rect 2349 2708 2365 2742
rect 2421 2708 2433 2742
rect 2493 2708 2501 2742
rect 2565 2708 2569 2742
rect 2671 2708 2708 2742
rect 2742 2708 2758 2742
rect 34 2692 2758 2708
rect 34 2671 100 2692
rect 34 2569 50 2671
rect 84 2569 100 2671
rect 34 2565 100 2569
rect 34 2501 50 2565
rect 84 2501 100 2565
rect 2692 2671 2758 2692
rect 2692 2569 2708 2671
rect 2742 2569 2758 2671
rect 2692 2565 2758 2569
rect 34 2493 100 2501
rect 34 2433 50 2493
rect 84 2433 100 2493
rect 34 2421 100 2433
rect 34 2365 50 2421
rect 84 2365 100 2421
rect 34 2349 100 2365
rect 34 2297 50 2349
rect 84 2297 100 2349
rect 34 2277 100 2297
rect 34 2229 50 2277
rect 84 2229 100 2277
rect 34 2205 100 2229
rect 34 2161 50 2205
rect 84 2161 100 2205
rect 34 2133 100 2161
rect 34 2093 50 2133
rect 84 2093 100 2133
rect 34 2061 100 2093
rect 34 2025 50 2061
rect 84 2025 100 2061
rect 34 1991 100 2025
rect 34 1955 50 1991
rect 84 1955 100 1991
rect 34 1923 100 1955
rect 34 1883 50 1923
rect 84 1883 100 1923
rect 34 1855 100 1883
rect 34 1811 50 1855
rect 84 1811 100 1855
rect 34 1787 100 1811
rect 34 1739 50 1787
rect 84 1739 100 1787
rect 34 1719 100 1739
rect 34 1667 50 1719
rect 84 1667 100 1719
rect 34 1651 100 1667
rect 34 1595 50 1651
rect 84 1595 100 1651
rect 34 1583 100 1595
rect 34 1523 50 1583
rect 84 1523 100 1583
rect 34 1515 100 1523
rect 34 1451 50 1515
rect 84 1451 100 1515
rect 34 1447 100 1451
rect 34 1345 50 1447
rect 84 1345 100 1447
rect 34 1341 100 1345
rect 34 1277 50 1341
rect 84 1277 100 1341
rect 34 1269 100 1277
rect 34 1209 50 1269
rect 84 1209 100 1269
rect 34 1197 100 1209
rect 34 1141 50 1197
rect 84 1141 100 1197
rect 34 1125 100 1141
rect 34 1073 50 1125
rect 84 1073 100 1125
rect 34 1053 100 1073
rect 34 1005 50 1053
rect 84 1005 100 1053
rect 34 981 100 1005
rect 34 937 50 981
rect 84 937 100 981
rect 34 909 100 937
rect 34 869 50 909
rect 84 869 100 909
rect 34 837 100 869
rect 34 801 50 837
rect 84 801 100 837
rect 34 767 100 801
rect 34 731 50 767
rect 84 731 100 767
rect 34 699 100 731
rect 34 659 50 699
rect 84 659 100 699
rect 34 631 100 659
rect 34 587 50 631
rect 84 587 100 631
rect 34 563 100 587
rect 34 515 50 563
rect 84 515 100 563
rect 34 495 100 515
rect 34 443 50 495
rect 84 443 100 495
rect 34 427 100 443
rect 34 371 50 427
rect 84 371 100 427
rect 34 359 100 371
rect 34 299 50 359
rect 84 299 100 359
rect 34 291 100 299
rect 34 227 50 291
rect 84 227 100 291
rect 260 2516 2532 2532
rect 260 2482 276 2516
rect 310 2482 359 2516
rect 405 2482 427 2516
rect 477 2482 495 2516
rect 549 2482 563 2516
rect 621 2482 631 2516
rect 693 2482 699 2516
rect 765 2482 767 2516
rect 801 2482 803 2516
rect 869 2482 875 2516
rect 937 2482 947 2516
rect 1005 2482 1019 2516
rect 1073 2482 1091 2516
rect 1141 2482 1163 2516
rect 1209 2482 1235 2516
rect 1277 2482 1307 2516
rect 1345 2482 1379 2516
rect 1413 2482 1447 2516
rect 1485 2482 1515 2516
rect 1557 2482 1583 2516
rect 1629 2482 1651 2516
rect 1701 2482 1719 2516
rect 1773 2482 1787 2516
rect 1845 2482 1855 2516
rect 1917 2482 1923 2516
rect 1989 2482 1991 2516
rect 2025 2482 2027 2516
rect 2093 2482 2099 2516
rect 2161 2482 2171 2516
rect 2229 2482 2243 2516
rect 2297 2482 2315 2516
rect 2365 2482 2387 2516
rect 2433 2482 2482 2516
rect 2516 2482 2532 2516
rect 260 2466 2532 2482
rect 260 2433 326 2466
rect 260 2387 276 2433
rect 310 2387 326 2433
rect 260 2365 326 2387
rect 260 2315 276 2365
rect 310 2315 326 2365
rect 260 2297 326 2315
rect 260 2243 276 2297
rect 310 2243 326 2297
rect 260 2229 326 2243
rect 260 2171 276 2229
rect 310 2171 326 2229
rect 260 2161 326 2171
rect 260 2099 276 2161
rect 310 2099 326 2161
rect 2466 2433 2532 2466
rect 2466 2387 2482 2433
rect 2516 2387 2532 2433
rect 2466 2365 2532 2387
rect 2466 2315 2482 2365
rect 2516 2315 2532 2365
rect 2466 2297 2532 2315
rect 2466 2243 2482 2297
rect 2516 2243 2532 2297
rect 2466 2229 2532 2243
rect 2466 2171 2482 2229
rect 2516 2171 2532 2229
rect 2466 2161 2532 2171
rect 260 2093 326 2099
rect 260 2027 276 2093
rect 310 2027 326 2093
rect 260 2025 326 2027
rect 260 1991 276 2025
rect 310 1991 326 2025
rect 260 1989 326 1991
rect 260 1923 276 1989
rect 310 1923 326 1989
rect 260 1917 326 1923
rect 260 1855 276 1917
rect 310 1855 326 1917
rect 260 1845 326 1855
rect 260 1787 276 1845
rect 310 1787 326 1845
rect 260 1773 326 1787
rect 260 1719 276 1773
rect 310 1719 326 1773
rect 260 1701 326 1719
rect 260 1651 276 1701
rect 310 1651 326 1701
rect 260 1629 326 1651
rect 260 1583 276 1629
rect 310 1583 326 1629
rect 260 1557 326 1583
rect 260 1515 276 1557
rect 310 1515 326 1557
rect 260 1485 326 1515
rect 260 1447 276 1485
rect 310 1447 326 1485
rect 260 1413 326 1447
rect 260 1379 276 1413
rect 310 1379 326 1413
rect 260 1345 326 1379
rect 260 1307 276 1345
rect 310 1307 326 1345
rect 260 1277 326 1307
rect 260 1235 276 1277
rect 310 1235 326 1277
rect 260 1209 326 1235
rect 260 1163 276 1209
rect 310 1163 326 1209
rect 260 1141 326 1163
rect 260 1091 276 1141
rect 310 1091 326 1141
rect 260 1073 326 1091
rect 260 1019 276 1073
rect 310 1019 326 1073
rect 260 1005 326 1019
rect 260 947 276 1005
rect 310 947 326 1005
rect 260 937 326 947
rect 260 875 276 937
rect 310 875 326 937
rect 260 869 326 875
rect 260 803 276 869
rect 310 803 326 869
rect 260 801 326 803
rect 260 767 276 801
rect 310 767 326 801
rect 260 765 326 767
rect 260 699 276 765
rect 310 699 326 765
rect 260 693 326 699
rect 260 631 276 693
rect 310 631 326 693
rect 662 2114 2130 2130
rect 662 2080 678 2114
rect 712 2080 767 2114
rect 801 2080 835 2114
rect 873 2080 903 2114
rect 945 2080 971 2114
rect 1017 2080 1039 2114
rect 1089 2080 1107 2114
rect 1161 2080 1175 2114
rect 1233 2080 1243 2114
rect 1305 2080 1311 2114
rect 1377 2080 1379 2114
rect 1413 2080 1415 2114
rect 1481 2080 1487 2114
rect 1549 2080 1559 2114
rect 1617 2080 1631 2114
rect 1685 2080 1703 2114
rect 1753 2080 1775 2114
rect 1821 2080 1847 2114
rect 1889 2080 1919 2114
rect 1957 2080 1991 2114
rect 2025 2080 2080 2114
rect 2114 2080 2130 2114
rect 662 2064 2130 2080
rect 662 2025 728 2064
rect 662 1991 678 2025
rect 712 1991 728 2025
rect 662 1957 728 1991
rect 662 1919 678 1957
rect 712 1919 728 1957
rect 662 1889 728 1919
rect 662 1847 678 1889
rect 712 1847 728 1889
rect 2064 2025 2130 2064
rect 2064 1991 2080 2025
rect 2114 1991 2130 2025
rect 2064 1957 2130 1991
rect 2064 1919 2080 1957
rect 2114 1919 2130 1957
rect 2064 1889 2130 1919
rect 662 1821 728 1847
rect 662 1775 678 1821
rect 712 1775 728 1821
rect 662 1753 728 1775
rect 662 1703 678 1753
rect 712 1703 728 1753
rect 662 1685 728 1703
rect 662 1631 678 1685
rect 712 1631 728 1685
rect 662 1617 728 1631
rect 662 1559 678 1617
rect 712 1559 728 1617
rect 662 1549 728 1559
rect 662 1487 678 1549
rect 712 1487 728 1549
rect 662 1481 728 1487
rect 662 1415 678 1481
rect 712 1415 728 1481
rect 662 1413 728 1415
rect 662 1379 678 1413
rect 712 1379 728 1413
rect 662 1377 728 1379
rect 662 1311 678 1377
rect 712 1311 728 1377
rect 662 1305 728 1311
rect 662 1243 678 1305
rect 712 1243 728 1305
rect 662 1233 728 1243
rect 662 1175 678 1233
rect 712 1175 728 1233
rect 662 1161 728 1175
rect 662 1107 678 1161
rect 712 1107 728 1161
rect 662 1089 728 1107
rect 662 1039 678 1089
rect 712 1039 728 1089
rect 662 1017 728 1039
rect 662 971 678 1017
rect 712 971 728 1017
rect 662 945 728 971
rect 662 903 678 945
rect 712 903 728 945
rect 921 1855 1871 1871
rect 921 937 937 1855
rect 1855 937 1871 1855
rect 921 921 1871 937
rect 2064 1847 2080 1889
rect 2114 1847 2130 1889
rect 2064 1821 2130 1847
rect 2064 1775 2080 1821
rect 2114 1775 2130 1821
rect 2064 1753 2130 1775
rect 2064 1703 2080 1753
rect 2114 1703 2130 1753
rect 2064 1685 2130 1703
rect 2064 1631 2080 1685
rect 2114 1631 2130 1685
rect 2064 1617 2130 1631
rect 2064 1559 2080 1617
rect 2114 1559 2130 1617
rect 2064 1549 2130 1559
rect 2064 1487 2080 1549
rect 2114 1487 2130 1549
rect 2064 1481 2130 1487
rect 2064 1415 2080 1481
rect 2114 1415 2130 1481
rect 2064 1413 2130 1415
rect 2064 1379 2080 1413
rect 2114 1379 2130 1413
rect 2064 1377 2130 1379
rect 2064 1311 2080 1377
rect 2114 1311 2130 1377
rect 2064 1305 2130 1311
rect 2064 1243 2080 1305
rect 2114 1243 2130 1305
rect 2064 1233 2130 1243
rect 2064 1175 2080 1233
rect 2114 1175 2130 1233
rect 2064 1161 2130 1175
rect 2064 1107 2080 1161
rect 2114 1107 2130 1161
rect 2064 1089 2130 1107
rect 2064 1039 2080 1089
rect 2114 1039 2130 1089
rect 2064 1017 2130 1039
rect 2064 971 2080 1017
rect 2114 971 2130 1017
rect 2064 945 2130 971
rect 662 873 728 903
rect 662 835 678 873
rect 712 835 728 873
rect 662 801 728 835
rect 662 767 678 801
rect 712 767 728 801
rect 662 728 728 767
rect 2064 903 2080 945
rect 2114 903 2130 945
rect 2064 873 2130 903
rect 2064 835 2080 873
rect 2114 835 2130 873
rect 2064 801 2130 835
rect 2064 767 2080 801
rect 2114 767 2130 801
rect 2064 728 2130 767
rect 662 712 2130 728
rect 662 678 678 712
rect 712 678 767 712
rect 801 678 835 712
rect 873 678 903 712
rect 945 678 971 712
rect 1017 678 1039 712
rect 1089 678 1107 712
rect 1161 678 1175 712
rect 1233 678 1243 712
rect 1305 678 1311 712
rect 1377 678 1379 712
rect 1413 678 1415 712
rect 1481 678 1487 712
rect 1549 678 1559 712
rect 1617 678 1631 712
rect 1685 678 1703 712
rect 1753 678 1775 712
rect 1821 678 1847 712
rect 1889 678 1919 712
rect 1957 678 1991 712
rect 2025 678 2080 712
rect 2114 678 2130 712
rect 662 662 2130 678
rect 2466 2099 2482 2161
rect 2516 2099 2532 2161
rect 2466 2093 2532 2099
rect 2466 2027 2482 2093
rect 2516 2027 2532 2093
rect 2466 2025 2532 2027
rect 2466 1991 2482 2025
rect 2516 1991 2532 2025
rect 2466 1989 2532 1991
rect 2466 1923 2482 1989
rect 2516 1923 2532 1989
rect 2466 1917 2532 1923
rect 2466 1855 2482 1917
rect 2516 1855 2532 1917
rect 2466 1845 2532 1855
rect 2466 1787 2482 1845
rect 2516 1787 2532 1845
rect 2466 1773 2532 1787
rect 2466 1719 2482 1773
rect 2516 1719 2532 1773
rect 2466 1701 2532 1719
rect 2466 1651 2482 1701
rect 2516 1651 2532 1701
rect 2466 1629 2532 1651
rect 2466 1583 2482 1629
rect 2516 1583 2532 1629
rect 2466 1557 2532 1583
rect 2466 1515 2482 1557
rect 2516 1515 2532 1557
rect 2466 1485 2532 1515
rect 2466 1447 2482 1485
rect 2516 1447 2532 1485
rect 2466 1413 2532 1447
rect 2466 1379 2482 1413
rect 2516 1379 2532 1413
rect 2466 1345 2532 1379
rect 2466 1307 2482 1345
rect 2516 1307 2532 1345
rect 2466 1277 2532 1307
rect 2466 1235 2482 1277
rect 2516 1235 2532 1277
rect 2466 1209 2532 1235
rect 2466 1163 2482 1209
rect 2516 1163 2532 1209
rect 2466 1141 2532 1163
rect 2466 1091 2482 1141
rect 2516 1091 2532 1141
rect 2466 1073 2532 1091
rect 2466 1019 2482 1073
rect 2516 1019 2532 1073
rect 2466 1005 2532 1019
rect 2466 947 2482 1005
rect 2516 947 2532 1005
rect 2466 937 2532 947
rect 2466 875 2482 937
rect 2516 875 2532 937
rect 2466 869 2532 875
rect 2466 803 2482 869
rect 2516 803 2532 869
rect 2466 801 2532 803
rect 2466 767 2482 801
rect 2516 767 2532 801
rect 2466 765 2532 767
rect 2466 699 2482 765
rect 2516 699 2532 765
rect 2466 693 2532 699
rect 260 621 326 631
rect 260 563 276 621
rect 310 563 326 621
rect 260 549 326 563
rect 260 495 276 549
rect 310 495 326 549
rect 260 477 326 495
rect 260 427 276 477
rect 310 427 326 477
rect 260 405 326 427
rect 260 359 276 405
rect 310 359 326 405
rect 260 326 326 359
rect 2466 631 2482 693
rect 2516 631 2532 693
rect 2466 621 2532 631
rect 2466 563 2482 621
rect 2516 563 2532 621
rect 2466 549 2532 563
rect 2466 495 2482 549
rect 2516 495 2532 549
rect 2466 477 2532 495
rect 2466 427 2482 477
rect 2516 427 2532 477
rect 2466 405 2532 427
rect 2466 359 2482 405
rect 2516 359 2532 405
rect 2466 326 2532 359
rect 260 310 2532 326
rect 260 276 276 310
rect 310 276 359 310
rect 405 276 427 310
rect 477 276 495 310
rect 549 276 563 310
rect 621 276 631 310
rect 693 276 699 310
rect 765 276 767 310
rect 801 276 803 310
rect 869 276 875 310
rect 937 276 947 310
rect 1005 276 1019 310
rect 1073 276 1091 310
rect 1141 276 1163 310
rect 1209 276 1235 310
rect 1277 276 1307 310
rect 1345 276 1379 310
rect 1413 276 1447 310
rect 1485 276 1515 310
rect 1557 276 1583 310
rect 1629 276 1651 310
rect 1701 276 1719 310
rect 1773 276 1787 310
rect 1845 276 1855 310
rect 1917 276 1923 310
rect 1989 276 1991 310
rect 2025 276 2027 310
rect 2093 276 2099 310
rect 2161 276 2171 310
rect 2229 276 2243 310
rect 2297 276 2315 310
rect 2365 276 2387 310
rect 2433 276 2482 310
rect 2516 276 2532 310
rect 260 260 2532 276
rect 2692 2501 2708 2565
rect 2742 2501 2758 2565
rect 2692 2493 2758 2501
rect 2692 2433 2708 2493
rect 2742 2433 2758 2493
rect 2692 2421 2758 2433
rect 2692 2365 2708 2421
rect 2742 2365 2758 2421
rect 2692 2349 2758 2365
rect 2692 2297 2708 2349
rect 2742 2297 2758 2349
rect 2692 2277 2758 2297
rect 2692 2229 2708 2277
rect 2742 2229 2758 2277
rect 2692 2205 2758 2229
rect 2692 2161 2708 2205
rect 2742 2161 2758 2205
rect 2692 2133 2758 2161
rect 2692 2093 2708 2133
rect 2742 2093 2758 2133
rect 2692 2061 2758 2093
rect 2692 2025 2708 2061
rect 2742 2025 2758 2061
rect 2692 1991 2758 2025
rect 2692 1955 2708 1991
rect 2742 1955 2758 1991
rect 2692 1923 2758 1955
rect 2692 1883 2708 1923
rect 2742 1883 2758 1923
rect 2692 1855 2758 1883
rect 2692 1811 2708 1855
rect 2742 1811 2758 1855
rect 2692 1787 2758 1811
rect 2692 1739 2708 1787
rect 2742 1739 2758 1787
rect 2692 1719 2758 1739
rect 2692 1667 2708 1719
rect 2742 1667 2758 1719
rect 2692 1651 2758 1667
rect 2692 1595 2708 1651
rect 2742 1595 2758 1651
rect 2692 1583 2758 1595
rect 2692 1523 2708 1583
rect 2742 1523 2758 1583
rect 2692 1515 2758 1523
rect 2692 1451 2708 1515
rect 2742 1451 2758 1515
rect 2692 1447 2758 1451
rect 2692 1345 2708 1447
rect 2742 1345 2758 1447
rect 2692 1341 2758 1345
rect 2692 1277 2708 1341
rect 2742 1277 2758 1341
rect 2692 1269 2758 1277
rect 2692 1209 2708 1269
rect 2742 1209 2758 1269
rect 2692 1197 2758 1209
rect 2692 1141 2708 1197
rect 2742 1141 2758 1197
rect 2692 1125 2758 1141
rect 2692 1073 2708 1125
rect 2742 1073 2758 1125
rect 2692 1053 2758 1073
rect 2692 1005 2708 1053
rect 2742 1005 2758 1053
rect 2692 981 2758 1005
rect 2692 937 2708 981
rect 2742 937 2758 981
rect 2692 909 2758 937
rect 2692 869 2708 909
rect 2742 869 2758 909
rect 2692 837 2758 869
rect 2692 801 2708 837
rect 2742 801 2758 837
rect 2692 767 2758 801
rect 2692 731 2708 767
rect 2742 731 2758 767
rect 2692 699 2758 731
rect 2692 659 2708 699
rect 2742 659 2758 699
rect 2692 631 2758 659
rect 2692 587 2708 631
rect 2742 587 2758 631
rect 2692 563 2758 587
rect 2692 515 2708 563
rect 2742 515 2758 563
rect 2692 495 2758 515
rect 2692 443 2708 495
rect 2742 443 2758 495
rect 2692 427 2758 443
rect 2692 371 2708 427
rect 2742 371 2758 427
rect 2692 359 2758 371
rect 2692 299 2708 359
rect 2742 299 2758 359
rect 2692 291 2758 299
rect 34 223 100 227
rect 34 121 50 223
rect 84 121 100 223
rect 34 100 100 121
rect 2692 227 2708 291
rect 2742 227 2758 291
rect 2692 223 2758 227
rect 2692 121 2708 223
rect 2742 121 2758 223
rect 2692 100 2758 121
rect 34 84 2758 100
rect 34 50 50 84
rect 84 50 121 84
rect 223 50 227 84
rect 291 50 299 84
rect 359 50 371 84
rect 427 50 443 84
rect 495 50 515 84
rect 563 50 587 84
rect 631 50 659 84
rect 699 50 731 84
rect 767 50 801 84
rect 837 50 869 84
rect 909 50 937 84
rect 981 50 1005 84
rect 1053 50 1073 84
rect 1125 50 1141 84
rect 1197 50 1209 84
rect 1269 50 1277 84
rect 1341 50 1345 84
rect 1447 50 1451 84
rect 1515 50 1523 84
rect 1583 50 1595 84
rect 1651 50 1667 84
rect 1719 50 1739 84
rect 1787 50 1811 84
rect 1855 50 1883 84
rect 1923 50 1955 84
rect 1991 50 2025 84
rect 2061 50 2093 84
rect 2133 50 2161 84
rect 2205 50 2229 84
rect 2277 50 2297 84
rect 2349 50 2365 84
rect 2421 50 2433 84
rect 2493 50 2501 84
rect 2565 50 2569 84
rect 2671 50 2708 84
rect 2742 50 2758 84
rect 34 34 2758 50
<< viali >>
rect 50 2708 84 2742
rect 155 2708 189 2742
rect 227 2708 257 2742
rect 257 2708 261 2742
rect 299 2708 325 2742
rect 325 2708 333 2742
rect 371 2708 393 2742
rect 393 2708 405 2742
rect 443 2708 461 2742
rect 461 2708 477 2742
rect 515 2708 529 2742
rect 529 2708 549 2742
rect 587 2708 597 2742
rect 597 2708 621 2742
rect 659 2708 665 2742
rect 665 2708 693 2742
rect 731 2708 733 2742
rect 733 2708 765 2742
rect 803 2708 835 2742
rect 835 2708 837 2742
rect 875 2708 903 2742
rect 903 2708 909 2742
rect 947 2708 971 2742
rect 971 2708 981 2742
rect 1019 2708 1039 2742
rect 1039 2708 1053 2742
rect 1091 2708 1107 2742
rect 1107 2708 1125 2742
rect 1163 2708 1175 2742
rect 1175 2708 1197 2742
rect 1235 2708 1243 2742
rect 1243 2708 1269 2742
rect 1307 2708 1311 2742
rect 1311 2708 1341 2742
rect 1379 2708 1413 2742
rect 1451 2708 1481 2742
rect 1481 2708 1485 2742
rect 1523 2708 1549 2742
rect 1549 2708 1557 2742
rect 1595 2708 1617 2742
rect 1617 2708 1629 2742
rect 1667 2708 1685 2742
rect 1685 2708 1701 2742
rect 1739 2708 1753 2742
rect 1753 2708 1773 2742
rect 1811 2708 1821 2742
rect 1821 2708 1845 2742
rect 1883 2708 1889 2742
rect 1889 2708 1917 2742
rect 1955 2708 1957 2742
rect 1957 2708 1989 2742
rect 2027 2708 2059 2742
rect 2059 2708 2061 2742
rect 2099 2708 2127 2742
rect 2127 2708 2133 2742
rect 2171 2708 2195 2742
rect 2195 2708 2205 2742
rect 2243 2708 2263 2742
rect 2263 2708 2277 2742
rect 2315 2708 2331 2742
rect 2331 2708 2349 2742
rect 2387 2708 2399 2742
rect 2399 2708 2421 2742
rect 2459 2708 2467 2742
rect 2467 2708 2493 2742
rect 2531 2708 2535 2742
rect 2535 2708 2565 2742
rect 2603 2708 2637 2742
rect 2708 2708 2742 2742
rect 50 2603 84 2637
rect 50 2535 84 2565
rect 50 2531 84 2535
rect 2708 2603 2742 2637
rect 50 2467 84 2493
rect 50 2459 84 2467
rect 50 2399 84 2421
rect 50 2387 84 2399
rect 50 2331 84 2349
rect 50 2315 84 2331
rect 50 2263 84 2277
rect 50 2243 84 2263
rect 50 2195 84 2205
rect 50 2171 84 2195
rect 50 2127 84 2133
rect 50 2099 84 2127
rect 50 2059 84 2061
rect 50 2027 84 2059
rect 50 1957 84 1989
rect 50 1955 84 1957
rect 50 1889 84 1917
rect 50 1883 84 1889
rect 50 1821 84 1845
rect 50 1811 84 1821
rect 50 1753 84 1773
rect 50 1739 84 1753
rect 50 1685 84 1701
rect 50 1667 84 1685
rect 50 1617 84 1629
rect 50 1595 84 1617
rect 50 1549 84 1557
rect 50 1523 84 1549
rect 50 1481 84 1485
rect 50 1451 84 1481
rect 50 1379 84 1413
rect 50 1311 84 1341
rect 50 1307 84 1311
rect 50 1243 84 1269
rect 50 1235 84 1243
rect 50 1175 84 1197
rect 50 1163 84 1175
rect 50 1107 84 1125
rect 50 1091 84 1107
rect 50 1039 84 1053
rect 50 1019 84 1039
rect 50 971 84 981
rect 50 947 84 971
rect 50 903 84 909
rect 50 875 84 903
rect 50 835 84 837
rect 50 803 84 835
rect 50 733 84 765
rect 50 731 84 733
rect 50 665 84 693
rect 50 659 84 665
rect 50 597 84 621
rect 50 587 84 597
rect 50 529 84 549
rect 50 515 84 529
rect 50 461 84 477
rect 50 443 84 461
rect 50 393 84 405
rect 50 371 84 393
rect 50 325 84 333
rect 50 299 84 325
rect 50 257 84 261
rect 50 227 84 257
rect 276 2482 310 2516
rect 371 2482 393 2516
rect 393 2482 405 2516
rect 443 2482 461 2516
rect 461 2482 477 2516
rect 515 2482 529 2516
rect 529 2482 549 2516
rect 587 2482 597 2516
rect 597 2482 621 2516
rect 659 2482 665 2516
rect 665 2482 693 2516
rect 731 2482 733 2516
rect 733 2482 765 2516
rect 803 2482 835 2516
rect 835 2482 837 2516
rect 875 2482 903 2516
rect 903 2482 909 2516
rect 947 2482 971 2516
rect 971 2482 981 2516
rect 1019 2482 1039 2516
rect 1039 2482 1053 2516
rect 1091 2482 1107 2516
rect 1107 2482 1125 2516
rect 1163 2482 1175 2516
rect 1175 2482 1197 2516
rect 1235 2482 1243 2516
rect 1243 2482 1269 2516
rect 1307 2482 1311 2516
rect 1311 2482 1341 2516
rect 1379 2482 1413 2516
rect 1451 2482 1481 2516
rect 1481 2482 1485 2516
rect 1523 2482 1549 2516
rect 1549 2482 1557 2516
rect 1595 2482 1617 2516
rect 1617 2482 1629 2516
rect 1667 2482 1685 2516
rect 1685 2482 1701 2516
rect 1739 2482 1753 2516
rect 1753 2482 1773 2516
rect 1811 2482 1821 2516
rect 1821 2482 1845 2516
rect 1883 2482 1889 2516
rect 1889 2482 1917 2516
rect 1955 2482 1957 2516
rect 1957 2482 1989 2516
rect 2027 2482 2059 2516
rect 2059 2482 2061 2516
rect 2099 2482 2127 2516
rect 2127 2482 2133 2516
rect 2171 2482 2195 2516
rect 2195 2482 2205 2516
rect 2243 2482 2263 2516
rect 2263 2482 2277 2516
rect 2315 2482 2331 2516
rect 2331 2482 2349 2516
rect 2387 2482 2399 2516
rect 2399 2482 2421 2516
rect 2482 2482 2516 2516
rect 276 2399 310 2421
rect 276 2387 310 2399
rect 276 2331 310 2349
rect 276 2315 310 2331
rect 276 2263 310 2277
rect 276 2243 310 2263
rect 276 2195 310 2205
rect 276 2171 310 2195
rect 276 2127 310 2133
rect 276 2099 310 2127
rect 2482 2399 2516 2421
rect 2482 2387 2516 2399
rect 2482 2331 2516 2349
rect 2482 2315 2516 2331
rect 2482 2263 2516 2277
rect 2482 2243 2516 2263
rect 2482 2195 2516 2205
rect 2482 2171 2516 2195
rect 276 2059 310 2061
rect 276 2027 310 2059
rect 276 1957 310 1989
rect 276 1955 310 1957
rect 276 1889 310 1917
rect 276 1883 310 1889
rect 276 1821 310 1845
rect 276 1811 310 1821
rect 276 1753 310 1773
rect 276 1739 310 1753
rect 276 1685 310 1701
rect 276 1667 310 1685
rect 276 1617 310 1629
rect 276 1595 310 1617
rect 276 1549 310 1557
rect 276 1523 310 1549
rect 276 1481 310 1485
rect 276 1451 310 1481
rect 276 1379 310 1413
rect 276 1311 310 1341
rect 276 1307 310 1311
rect 276 1243 310 1269
rect 276 1235 310 1243
rect 276 1175 310 1197
rect 276 1163 310 1175
rect 276 1107 310 1125
rect 276 1091 310 1107
rect 276 1039 310 1053
rect 276 1019 310 1039
rect 276 971 310 981
rect 276 947 310 971
rect 276 903 310 909
rect 276 875 310 903
rect 276 835 310 837
rect 276 803 310 835
rect 276 733 310 765
rect 276 731 310 733
rect 276 665 310 693
rect 276 659 310 665
rect 678 2080 712 2114
rect 767 2080 801 2114
rect 839 2080 869 2114
rect 869 2080 873 2114
rect 911 2080 937 2114
rect 937 2080 945 2114
rect 983 2080 1005 2114
rect 1005 2080 1017 2114
rect 1055 2080 1073 2114
rect 1073 2080 1089 2114
rect 1127 2080 1141 2114
rect 1141 2080 1161 2114
rect 1199 2080 1209 2114
rect 1209 2080 1233 2114
rect 1271 2080 1277 2114
rect 1277 2080 1305 2114
rect 1343 2080 1345 2114
rect 1345 2080 1377 2114
rect 1415 2080 1447 2114
rect 1447 2080 1449 2114
rect 1487 2080 1515 2114
rect 1515 2080 1521 2114
rect 1559 2080 1583 2114
rect 1583 2080 1593 2114
rect 1631 2080 1651 2114
rect 1651 2080 1665 2114
rect 1703 2080 1719 2114
rect 1719 2080 1737 2114
rect 1775 2080 1787 2114
rect 1787 2080 1809 2114
rect 1847 2080 1855 2114
rect 1855 2080 1881 2114
rect 1919 2080 1923 2114
rect 1923 2080 1953 2114
rect 1991 2080 2025 2114
rect 2080 2080 2114 2114
rect 678 1991 712 2025
rect 678 1923 712 1953
rect 678 1919 712 1923
rect 678 1855 712 1881
rect 678 1847 712 1855
rect 2080 1991 2114 2025
rect 2080 1923 2114 1953
rect 2080 1919 2114 1923
rect 678 1787 712 1809
rect 678 1775 712 1787
rect 678 1719 712 1737
rect 678 1703 712 1719
rect 678 1651 712 1665
rect 678 1631 712 1651
rect 678 1583 712 1593
rect 678 1559 712 1583
rect 678 1515 712 1521
rect 678 1487 712 1515
rect 678 1447 712 1449
rect 678 1415 712 1447
rect 678 1345 712 1377
rect 678 1343 712 1345
rect 678 1277 712 1305
rect 678 1271 712 1277
rect 678 1209 712 1233
rect 678 1199 712 1209
rect 678 1141 712 1161
rect 678 1127 712 1141
rect 678 1073 712 1089
rect 678 1055 712 1073
rect 678 1005 712 1017
rect 678 983 712 1005
rect 678 937 712 945
rect 678 911 712 937
rect 947 947 1845 1845
rect 2080 1855 2114 1881
rect 2080 1847 2114 1855
rect 2080 1787 2114 1809
rect 2080 1775 2114 1787
rect 2080 1719 2114 1737
rect 2080 1703 2114 1719
rect 2080 1651 2114 1665
rect 2080 1631 2114 1651
rect 2080 1583 2114 1593
rect 2080 1559 2114 1583
rect 2080 1515 2114 1521
rect 2080 1487 2114 1515
rect 2080 1447 2114 1449
rect 2080 1415 2114 1447
rect 2080 1345 2114 1377
rect 2080 1343 2114 1345
rect 2080 1277 2114 1305
rect 2080 1271 2114 1277
rect 2080 1209 2114 1233
rect 2080 1199 2114 1209
rect 2080 1141 2114 1161
rect 2080 1127 2114 1141
rect 2080 1073 2114 1089
rect 2080 1055 2114 1073
rect 2080 1005 2114 1017
rect 2080 983 2114 1005
rect 678 869 712 873
rect 678 839 712 869
rect 678 767 712 801
rect 2080 937 2114 945
rect 2080 911 2114 937
rect 2080 869 2114 873
rect 2080 839 2114 869
rect 2080 767 2114 801
rect 678 678 712 712
rect 767 678 801 712
rect 839 678 869 712
rect 869 678 873 712
rect 911 678 937 712
rect 937 678 945 712
rect 983 678 1005 712
rect 1005 678 1017 712
rect 1055 678 1073 712
rect 1073 678 1089 712
rect 1127 678 1141 712
rect 1141 678 1161 712
rect 1199 678 1209 712
rect 1209 678 1233 712
rect 1271 678 1277 712
rect 1277 678 1305 712
rect 1343 678 1345 712
rect 1345 678 1377 712
rect 1415 678 1447 712
rect 1447 678 1449 712
rect 1487 678 1515 712
rect 1515 678 1521 712
rect 1559 678 1583 712
rect 1583 678 1593 712
rect 1631 678 1651 712
rect 1651 678 1665 712
rect 1703 678 1719 712
rect 1719 678 1737 712
rect 1775 678 1787 712
rect 1787 678 1809 712
rect 1847 678 1855 712
rect 1855 678 1881 712
rect 1919 678 1923 712
rect 1923 678 1953 712
rect 1991 678 2025 712
rect 2080 678 2114 712
rect 2482 2127 2516 2133
rect 2482 2099 2516 2127
rect 2482 2059 2516 2061
rect 2482 2027 2516 2059
rect 2482 1957 2516 1989
rect 2482 1955 2516 1957
rect 2482 1889 2516 1917
rect 2482 1883 2516 1889
rect 2482 1821 2516 1845
rect 2482 1811 2516 1821
rect 2482 1753 2516 1773
rect 2482 1739 2516 1753
rect 2482 1685 2516 1701
rect 2482 1667 2516 1685
rect 2482 1617 2516 1629
rect 2482 1595 2516 1617
rect 2482 1549 2516 1557
rect 2482 1523 2516 1549
rect 2482 1481 2516 1485
rect 2482 1451 2516 1481
rect 2482 1379 2516 1413
rect 2482 1311 2516 1341
rect 2482 1307 2516 1311
rect 2482 1243 2516 1269
rect 2482 1235 2516 1243
rect 2482 1175 2516 1197
rect 2482 1163 2516 1175
rect 2482 1107 2516 1125
rect 2482 1091 2516 1107
rect 2482 1039 2516 1053
rect 2482 1019 2516 1039
rect 2482 971 2516 981
rect 2482 947 2516 971
rect 2482 903 2516 909
rect 2482 875 2516 903
rect 2482 835 2516 837
rect 2482 803 2516 835
rect 2482 733 2516 765
rect 2482 731 2516 733
rect 276 597 310 621
rect 276 587 310 597
rect 276 529 310 549
rect 276 515 310 529
rect 276 461 310 477
rect 276 443 310 461
rect 276 393 310 405
rect 276 371 310 393
rect 2482 665 2516 693
rect 2482 659 2516 665
rect 2482 597 2516 621
rect 2482 587 2516 597
rect 2482 529 2516 549
rect 2482 515 2516 529
rect 2482 461 2516 477
rect 2482 443 2516 461
rect 2482 393 2516 405
rect 2482 371 2516 393
rect 276 276 310 310
rect 371 276 393 310
rect 393 276 405 310
rect 443 276 461 310
rect 461 276 477 310
rect 515 276 529 310
rect 529 276 549 310
rect 587 276 597 310
rect 597 276 621 310
rect 659 276 665 310
rect 665 276 693 310
rect 731 276 733 310
rect 733 276 765 310
rect 803 276 835 310
rect 835 276 837 310
rect 875 276 903 310
rect 903 276 909 310
rect 947 276 971 310
rect 971 276 981 310
rect 1019 276 1039 310
rect 1039 276 1053 310
rect 1091 276 1107 310
rect 1107 276 1125 310
rect 1163 276 1175 310
rect 1175 276 1197 310
rect 1235 276 1243 310
rect 1243 276 1269 310
rect 1307 276 1311 310
rect 1311 276 1341 310
rect 1379 276 1413 310
rect 1451 276 1481 310
rect 1481 276 1485 310
rect 1523 276 1549 310
rect 1549 276 1557 310
rect 1595 276 1617 310
rect 1617 276 1629 310
rect 1667 276 1685 310
rect 1685 276 1701 310
rect 1739 276 1753 310
rect 1753 276 1773 310
rect 1811 276 1821 310
rect 1821 276 1845 310
rect 1883 276 1889 310
rect 1889 276 1917 310
rect 1955 276 1957 310
rect 1957 276 1989 310
rect 2027 276 2059 310
rect 2059 276 2061 310
rect 2099 276 2127 310
rect 2127 276 2133 310
rect 2171 276 2195 310
rect 2195 276 2205 310
rect 2243 276 2263 310
rect 2263 276 2277 310
rect 2315 276 2331 310
rect 2331 276 2349 310
rect 2387 276 2399 310
rect 2399 276 2421 310
rect 2482 276 2516 310
rect 2708 2535 2742 2565
rect 2708 2531 2742 2535
rect 2708 2467 2742 2493
rect 2708 2459 2742 2467
rect 2708 2399 2742 2421
rect 2708 2387 2742 2399
rect 2708 2331 2742 2349
rect 2708 2315 2742 2331
rect 2708 2263 2742 2277
rect 2708 2243 2742 2263
rect 2708 2195 2742 2205
rect 2708 2171 2742 2195
rect 2708 2127 2742 2133
rect 2708 2099 2742 2127
rect 2708 2059 2742 2061
rect 2708 2027 2742 2059
rect 2708 1957 2742 1989
rect 2708 1955 2742 1957
rect 2708 1889 2742 1917
rect 2708 1883 2742 1889
rect 2708 1821 2742 1845
rect 2708 1811 2742 1821
rect 2708 1753 2742 1773
rect 2708 1739 2742 1753
rect 2708 1685 2742 1701
rect 2708 1667 2742 1685
rect 2708 1617 2742 1629
rect 2708 1595 2742 1617
rect 2708 1549 2742 1557
rect 2708 1523 2742 1549
rect 2708 1481 2742 1485
rect 2708 1451 2742 1481
rect 2708 1379 2742 1413
rect 2708 1311 2742 1341
rect 2708 1307 2742 1311
rect 2708 1243 2742 1269
rect 2708 1235 2742 1243
rect 2708 1175 2742 1197
rect 2708 1163 2742 1175
rect 2708 1107 2742 1125
rect 2708 1091 2742 1107
rect 2708 1039 2742 1053
rect 2708 1019 2742 1039
rect 2708 971 2742 981
rect 2708 947 2742 971
rect 2708 903 2742 909
rect 2708 875 2742 903
rect 2708 835 2742 837
rect 2708 803 2742 835
rect 2708 733 2742 765
rect 2708 731 2742 733
rect 2708 665 2742 693
rect 2708 659 2742 665
rect 2708 597 2742 621
rect 2708 587 2742 597
rect 2708 529 2742 549
rect 2708 515 2742 529
rect 2708 461 2742 477
rect 2708 443 2742 461
rect 2708 393 2742 405
rect 2708 371 2742 393
rect 2708 325 2742 333
rect 2708 299 2742 325
rect 50 155 84 189
rect 2708 257 2742 261
rect 2708 227 2742 257
rect 2708 155 2742 189
rect 50 50 84 84
rect 155 50 189 84
rect 227 50 257 84
rect 257 50 261 84
rect 299 50 325 84
rect 325 50 333 84
rect 371 50 393 84
rect 393 50 405 84
rect 443 50 461 84
rect 461 50 477 84
rect 515 50 529 84
rect 529 50 549 84
rect 587 50 597 84
rect 597 50 621 84
rect 659 50 665 84
rect 665 50 693 84
rect 731 50 733 84
rect 733 50 765 84
rect 803 50 835 84
rect 835 50 837 84
rect 875 50 903 84
rect 903 50 909 84
rect 947 50 971 84
rect 971 50 981 84
rect 1019 50 1039 84
rect 1039 50 1053 84
rect 1091 50 1107 84
rect 1107 50 1125 84
rect 1163 50 1175 84
rect 1175 50 1197 84
rect 1235 50 1243 84
rect 1243 50 1269 84
rect 1307 50 1311 84
rect 1311 50 1341 84
rect 1379 50 1413 84
rect 1451 50 1481 84
rect 1481 50 1485 84
rect 1523 50 1549 84
rect 1549 50 1557 84
rect 1595 50 1617 84
rect 1617 50 1629 84
rect 1667 50 1685 84
rect 1685 50 1701 84
rect 1739 50 1753 84
rect 1753 50 1773 84
rect 1811 50 1821 84
rect 1821 50 1845 84
rect 1883 50 1889 84
rect 1889 50 1917 84
rect 1955 50 1957 84
rect 1957 50 1989 84
rect 2027 50 2059 84
rect 2059 50 2061 84
rect 2099 50 2127 84
rect 2127 50 2133 84
rect 2171 50 2195 84
rect 2195 50 2205 84
rect 2243 50 2263 84
rect 2263 50 2277 84
rect 2315 50 2331 84
rect 2331 50 2349 84
rect 2387 50 2399 84
rect 2399 50 2421 84
rect 2459 50 2467 84
rect 2467 50 2493 84
rect 2531 50 2535 84
rect 2535 50 2565 84
rect 2603 50 2637 84
rect 2708 50 2742 84
<< metal1 >>
rect 38 2742 2754 2754
rect 38 2708 50 2742
rect 84 2708 155 2742
rect 189 2708 227 2742
rect 261 2708 299 2742
rect 333 2708 371 2742
rect 405 2708 443 2742
rect 477 2708 515 2742
rect 549 2708 587 2742
rect 621 2708 659 2742
rect 693 2708 731 2742
rect 765 2708 803 2742
rect 837 2708 875 2742
rect 909 2708 947 2742
rect 981 2708 1019 2742
rect 1053 2708 1091 2742
rect 1125 2708 1163 2742
rect 1197 2708 1235 2742
rect 1269 2708 1307 2742
rect 1341 2708 1379 2742
rect 1413 2708 1451 2742
rect 1485 2708 1523 2742
rect 1557 2708 1595 2742
rect 1629 2708 1667 2742
rect 1701 2708 1739 2742
rect 1773 2708 1811 2742
rect 1845 2708 1883 2742
rect 1917 2708 1955 2742
rect 1989 2708 2027 2742
rect 2061 2708 2099 2742
rect 2133 2708 2171 2742
rect 2205 2708 2243 2742
rect 2277 2708 2315 2742
rect 2349 2708 2387 2742
rect 2421 2708 2459 2742
rect 2493 2708 2531 2742
rect 2565 2708 2603 2742
rect 2637 2708 2708 2742
rect 2742 2708 2754 2742
rect 38 2696 2754 2708
rect 38 2637 96 2696
rect 38 2603 50 2637
rect 84 2603 96 2637
rect 38 2565 96 2603
rect 38 2531 50 2565
rect 84 2531 96 2565
rect 38 2493 96 2531
rect 2696 2637 2754 2696
rect 2696 2603 2708 2637
rect 2742 2603 2754 2637
rect 2696 2565 2754 2603
rect 2696 2531 2708 2565
rect 2742 2531 2754 2565
rect 38 2459 50 2493
rect 84 2459 96 2493
rect 38 2421 96 2459
rect 38 2387 50 2421
rect 84 2387 96 2421
rect 38 2349 96 2387
rect 38 2315 50 2349
rect 84 2315 96 2349
rect 38 2277 96 2315
rect 38 2243 50 2277
rect 84 2243 96 2277
rect 38 2205 96 2243
rect 38 2171 50 2205
rect 84 2171 96 2205
rect 38 2133 96 2171
rect 38 2099 50 2133
rect 84 2099 96 2133
rect 38 2061 96 2099
rect 38 2027 50 2061
rect 84 2027 96 2061
rect 38 1989 96 2027
rect 38 1955 50 1989
rect 84 1955 96 1989
rect 38 1917 96 1955
rect 38 1883 50 1917
rect 84 1883 96 1917
rect 38 1845 96 1883
rect 38 1811 50 1845
rect 84 1811 96 1845
rect 38 1773 96 1811
rect 38 1739 50 1773
rect 84 1739 96 1773
rect 38 1701 96 1739
rect 38 1667 50 1701
rect 84 1667 96 1701
rect 38 1629 96 1667
rect 38 1595 50 1629
rect 84 1595 96 1629
rect 38 1557 96 1595
rect 38 1523 50 1557
rect 84 1523 96 1557
rect 38 1485 96 1523
rect 38 1451 50 1485
rect 84 1451 96 1485
rect 38 1413 96 1451
rect 38 1379 50 1413
rect 84 1379 96 1413
rect 38 1341 96 1379
rect 38 1307 50 1341
rect 84 1307 96 1341
rect 38 1269 96 1307
rect 38 1235 50 1269
rect 84 1235 96 1269
rect 38 1197 96 1235
rect 38 1163 50 1197
rect 84 1163 96 1197
rect 38 1125 96 1163
rect 38 1091 50 1125
rect 84 1091 96 1125
rect 38 1053 96 1091
rect 38 1019 50 1053
rect 84 1019 96 1053
rect 38 981 96 1019
rect 38 947 50 981
rect 84 947 96 981
rect 38 909 96 947
rect 38 875 50 909
rect 84 875 96 909
rect 38 837 96 875
rect 38 803 50 837
rect 84 803 96 837
rect 38 765 96 803
rect 38 731 50 765
rect 84 731 96 765
rect 38 693 96 731
rect 38 659 50 693
rect 84 659 96 693
rect 38 621 96 659
rect 38 587 50 621
rect 84 587 96 621
rect 38 549 96 587
rect 38 515 50 549
rect 84 515 96 549
rect 38 477 96 515
rect 38 443 50 477
rect 84 443 96 477
rect 38 405 96 443
rect 38 371 50 405
rect 84 371 96 405
rect 38 333 96 371
rect 38 299 50 333
rect 84 299 96 333
rect 38 261 96 299
rect 264 2516 2528 2528
rect 264 2482 276 2516
rect 310 2482 371 2516
rect 405 2482 443 2516
rect 477 2482 515 2516
rect 549 2482 587 2516
rect 621 2482 659 2516
rect 693 2482 731 2516
rect 765 2482 803 2516
rect 837 2482 875 2516
rect 909 2482 947 2516
rect 981 2482 1019 2516
rect 1053 2482 1091 2516
rect 1125 2482 1163 2516
rect 1197 2482 1235 2516
rect 1269 2482 1307 2516
rect 1341 2482 1379 2516
rect 1413 2482 1451 2516
rect 1485 2482 1523 2516
rect 1557 2482 1595 2516
rect 1629 2482 1667 2516
rect 1701 2482 1739 2516
rect 1773 2482 1811 2516
rect 1845 2482 1883 2516
rect 1917 2482 1955 2516
rect 1989 2482 2027 2516
rect 2061 2482 2099 2516
rect 2133 2482 2171 2516
rect 2205 2482 2243 2516
rect 2277 2482 2315 2516
rect 2349 2482 2387 2516
rect 2421 2482 2482 2516
rect 2516 2482 2528 2516
rect 264 2470 2528 2482
rect 264 2421 322 2470
rect 264 2387 276 2421
rect 310 2387 322 2421
rect 264 2349 322 2387
rect 264 2315 276 2349
rect 310 2315 322 2349
rect 264 2277 322 2315
rect 264 2243 276 2277
rect 310 2243 322 2277
rect 264 2205 322 2243
rect 264 2171 276 2205
rect 310 2171 322 2205
rect 264 2133 322 2171
rect 264 2099 276 2133
rect 310 2099 322 2133
rect 2470 2421 2528 2470
rect 2470 2387 2482 2421
rect 2516 2387 2528 2421
rect 2470 2349 2528 2387
rect 2470 2315 2482 2349
rect 2516 2315 2528 2349
rect 2470 2277 2528 2315
rect 2470 2243 2482 2277
rect 2516 2243 2528 2277
rect 2470 2205 2528 2243
rect 2470 2171 2482 2205
rect 2516 2171 2528 2205
rect 2470 2133 2528 2171
rect 264 2061 322 2099
rect 264 2027 276 2061
rect 310 2027 322 2061
rect 264 1989 322 2027
rect 264 1955 276 1989
rect 310 1955 322 1989
rect 264 1917 322 1955
rect 264 1883 276 1917
rect 310 1883 322 1917
rect 264 1845 322 1883
rect 264 1811 276 1845
rect 310 1811 322 1845
rect 264 1773 322 1811
rect 264 1739 276 1773
rect 310 1739 322 1773
rect 264 1701 322 1739
rect 264 1667 276 1701
rect 310 1667 322 1701
rect 264 1629 322 1667
rect 264 1595 276 1629
rect 310 1595 322 1629
rect 264 1557 322 1595
rect 264 1523 276 1557
rect 310 1523 322 1557
rect 264 1485 322 1523
rect 264 1451 276 1485
rect 310 1451 322 1485
rect 264 1413 322 1451
rect 264 1379 276 1413
rect 310 1379 322 1413
rect 264 1341 322 1379
rect 264 1307 276 1341
rect 310 1307 322 1341
rect 264 1269 322 1307
rect 264 1235 276 1269
rect 310 1235 322 1269
rect 264 1197 322 1235
rect 264 1163 276 1197
rect 310 1163 322 1197
rect 264 1125 322 1163
rect 264 1091 276 1125
rect 310 1091 322 1125
rect 264 1053 322 1091
rect 264 1019 276 1053
rect 310 1019 322 1053
rect 264 981 322 1019
rect 264 947 276 981
rect 310 947 322 981
rect 264 909 322 947
rect 264 875 276 909
rect 310 875 322 909
rect 264 837 322 875
rect 264 803 276 837
rect 310 803 322 837
rect 264 765 322 803
rect 264 731 276 765
rect 310 731 322 765
rect 264 693 322 731
rect 264 659 276 693
rect 310 659 322 693
rect 666 2114 2126 2126
rect 666 2080 678 2114
rect 712 2080 767 2114
rect 801 2080 839 2114
rect 873 2080 911 2114
rect 945 2080 983 2114
rect 1017 2080 1055 2114
rect 1089 2080 1127 2114
rect 1161 2080 1199 2114
rect 1233 2080 1271 2114
rect 1305 2080 1343 2114
rect 1377 2080 1415 2114
rect 1449 2080 1487 2114
rect 1521 2080 1559 2114
rect 1593 2080 1631 2114
rect 1665 2080 1703 2114
rect 1737 2080 1775 2114
rect 1809 2080 1847 2114
rect 1881 2080 1919 2114
rect 1953 2080 1991 2114
rect 2025 2080 2080 2114
rect 2114 2080 2126 2114
rect 666 2068 2126 2080
rect 666 2025 724 2068
rect 666 1991 678 2025
rect 712 1991 724 2025
rect 666 1953 724 1991
rect 666 1919 678 1953
rect 712 1919 724 1953
rect 666 1881 724 1919
rect 666 1847 678 1881
rect 712 1847 724 1881
rect 2068 2025 2126 2068
rect 2068 1991 2080 2025
rect 2114 1991 2126 2025
rect 2068 1953 2126 1991
rect 2068 1919 2080 1953
rect 2114 1919 2126 1953
rect 2068 1881 2126 1919
rect 666 1809 724 1847
rect 666 1775 678 1809
rect 712 1775 724 1809
rect 666 1737 724 1775
rect 666 1703 678 1737
rect 712 1703 724 1737
rect 666 1665 724 1703
rect 666 1631 678 1665
rect 712 1631 724 1665
rect 666 1593 724 1631
rect 666 1559 678 1593
rect 712 1559 724 1593
rect 666 1521 724 1559
rect 666 1487 678 1521
rect 712 1487 724 1521
rect 666 1449 724 1487
rect 666 1415 678 1449
rect 712 1415 724 1449
rect 666 1377 724 1415
rect 666 1343 678 1377
rect 712 1343 724 1377
rect 666 1305 724 1343
rect 666 1271 678 1305
rect 712 1271 724 1305
rect 666 1233 724 1271
rect 666 1199 678 1233
rect 712 1199 724 1233
rect 666 1161 724 1199
rect 666 1127 678 1161
rect 712 1127 724 1161
rect 666 1089 724 1127
rect 666 1055 678 1089
rect 712 1055 724 1089
rect 666 1017 724 1055
rect 666 983 678 1017
rect 712 983 724 1017
rect 666 945 724 983
rect 666 911 678 945
rect 712 911 724 945
rect 935 1845 1857 1857
rect 935 947 947 1845
rect 1845 947 1857 1845
rect 935 935 1857 947
rect 2068 1847 2080 1881
rect 2114 1847 2126 1881
rect 2068 1809 2126 1847
rect 2068 1775 2080 1809
rect 2114 1775 2126 1809
rect 2068 1737 2126 1775
rect 2068 1703 2080 1737
rect 2114 1703 2126 1737
rect 2068 1665 2126 1703
rect 2068 1631 2080 1665
rect 2114 1631 2126 1665
rect 2068 1593 2126 1631
rect 2068 1559 2080 1593
rect 2114 1559 2126 1593
rect 2068 1521 2126 1559
rect 2068 1487 2080 1521
rect 2114 1487 2126 1521
rect 2068 1449 2126 1487
rect 2068 1415 2080 1449
rect 2114 1415 2126 1449
rect 2068 1377 2126 1415
rect 2068 1343 2080 1377
rect 2114 1343 2126 1377
rect 2068 1305 2126 1343
rect 2068 1271 2080 1305
rect 2114 1271 2126 1305
rect 2068 1233 2126 1271
rect 2068 1199 2080 1233
rect 2114 1199 2126 1233
rect 2068 1161 2126 1199
rect 2068 1127 2080 1161
rect 2114 1127 2126 1161
rect 2068 1089 2126 1127
rect 2068 1055 2080 1089
rect 2114 1055 2126 1089
rect 2068 1017 2126 1055
rect 2068 983 2080 1017
rect 2114 983 2126 1017
rect 2068 945 2126 983
rect 666 873 724 911
rect 666 839 678 873
rect 712 839 724 873
rect 666 801 724 839
rect 666 767 678 801
rect 712 767 724 801
rect 666 724 724 767
rect 2068 911 2080 945
rect 2114 911 2126 945
rect 2068 873 2126 911
rect 2068 839 2080 873
rect 2114 839 2126 873
rect 2068 801 2126 839
rect 2068 767 2080 801
rect 2114 767 2126 801
rect 2068 724 2126 767
rect 666 712 2126 724
rect 666 678 678 712
rect 712 678 767 712
rect 801 678 839 712
rect 873 678 911 712
rect 945 678 983 712
rect 1017 678 1055 712
rect 1089 678 1127 712
rect 1161 678 1199 712
rect 1233 678 1271 712
rect 1305 678 1343 712
rect 1377 678 1415 712
rect 1449 678 1487 712
rect 1521 678 1559 712
rect 1593 678 1631 712
rect 1665 678 1703 712
rect 1737 678 1775 712
rect 1809 678 1847 712
rect 1881 678 1919 712
rect 1953 678 1991 712
rect 2025 678 2080 712
rect 2114 678 2126 712
rect 666 666 2126 678
rect 2470 2099 2482 2133
rect 2516 2099 2528 2133
rect 2470 2061 2528 2099
rect 2470 2027 2482 2061
rect 2516 2027 2528 2061
rect 2470 1989 2528 2027
rect 2470 1955 2482 1989
rect 2516 1955 2528 1989
rect 2470 1917 2528 1955
rect 2470 1883 2482 1917
rect 2516 1883 2528 1917
rect 2470 1845 2528 1883
rect 2470 1811 2482 1845
rect 2516 1811 2528 1845
rect 2470 1773 2528 1811
rect 2470 1739 2482 1773
rect 2516 1739 2528 1773
rect 2470 1701 2528 1739
rect 2470 1667 2482 1701
rect 2516 1667 2528 1701
rect 2470 1629 2528 1667
rect 2470 1595 2482 1629
rect 2516 1595 2528 1629
rect 2470 1557 2528 1595
rect 2470 1523 2482 1557
rect 2516 1523 2528 1557
rect 2470 1485 2528 1523
rect 2470 1451 2482 1485
rect 2516 1451 2528 1485
rect 2470 1413 2528 1451
rect 2470 1379 2482 1413
rect 2516 1379 2528 1413
rect 2470 1341 2528 1379
rect 2470 1307 2482 1341
rect 2516 1307 2528 1341
rect 2470 1269 2528 1307
rect 2470 1235 2482 1269
rect 2516 1235 2528 1269
rect 2470 1197 2528 1235
rect 2470 1163 2482 1197
rect 2516 1163 2528 1197
rect 2470 1125 2528 1163
rect 2470 1091 2482 1125
rect 2516 1091 2528 1125
rect 2470 1053 2528 1091
rect 2470 1019 2482 1053
rect 2516 1019 2528 1053
rect 2470 981 2528 1019
rect 2470 947 2482 981
rect 2516 947 2528 981
rect 2470 909 2528 947
rect 2470 875 2482 909
rect 2516 875 2528 909
rect 2470 837 2528 875
rect 2470 803 2482 837
rect 2516 803 2528 837
rect 2470 765 2528 803
rect 2470 731 2482 765
rect 2516 731 2528 765
rect 2470 693 2528 731
rect 264 621 322 659
rect 264 587 276 621
rect 310 587 322 621
rect 264 549 322 587
rect 264 515 276 549
rect 310 515 322 549
rect 264 477 322 515
rect 264 443 276 477
rect 310 443 322 477
rect 264 405 322 443
rect 264 371 276 405
rect 310 371 322 405
rect 264 322 322 371
rect 2470 659 2482 693
rect 2516 659 2528 693
rect 2470 621 2528 659
rect 2470 587 2482 621
rect 2516 587 2528 621
rect 2470 549 2528 587
rect 2470 515 2482 549
rect 2516 515 2528 549
rect 2470 477 2528 515
rect 2470 443 2482 477
rect 2516 443 2528 477
rect 2470 405 2528 443
rect 2470 371 2482 405
rect 2516 371 2528 405
rect 2470 322 2528 371
rect 264 310 2528 322
rect 264 276 276 310
rect 310 276 371 310
rect 405 276 443 310
rect 477 276 515 310
rect 549 276 587 310
rect 621 276 659 310
rect 693 276 731 310
rect 765 276 803 310
rect 837 276 875 310
rect 909 276 947 310
rect 981 276 1019 310
rect 1053 276 1091 310
rect 1125 276 1163 310
rect 1197 276 1235 310
rect 1269 276 1307 310
rect 1341 276 1379 310
rect 1413 276 1451 310
rect 1485 276 1523 310
rect 1557 276 1595 310
rect 1629 276 1667 310
rect 1701 276 1739 310
rect 1773 276 1811 310
rect 1845 276 1883 310
rect 1917 276 1955 310
rect 1989 276 2027 310
rect 2061 276 2099 310
rect 2133 276 2171 310
rect 2205 276 2243 310
rect 2277 276 2315 310
rect 2349 276 2387 310
rect 2421 276 2482 310
rect 2516 276 2528 310
rect 264 264 2528 276
rect 2696 2493 2754 2531
rect 2696 2459 2708 2493
rect 2742 2459 2754 2493
rect 2696 2421 2754 2459
rect 2696 2387 2708 2421
rect 2742 2387 2754 2421
rect 2696 2349 2754 2387
rect 2696 2315 2708 2349
rect 2742 2315 2754 2349
rect 2696 2277 2754 2315
rect 2696 2243 2708 2277
rect 2742 2243 2754 2277
rect 2696 2205 2754 2243
rect 2696 2171 2708 2205
rect 2742 2171 2754 2205
rect 2696 2133 2754 2171
rect 2696 2099 2708 2133
rect 2742 2099 2754 2133
rect 2696 2061 2754 2099
rect 2696 2027 2708 2061
rect 2742 2027 2754 2061
rect 2696 1989 2754 2027
rect 2696 1955 2708 1989
rect 2742 1955 2754 1989
rect 2696 1917 2754 1955
rect 2696 1883 2708 1917
rect 2742 1883 2754 1917
rect 2696 1845 2754 1883
rect 2696 1811 2708 1845
rect 2742 1811 2754 1845
rect 2696 1773 2754 1811
rect 2696 1739 2708 1773
rect 2742 1739 2754 1773
rect 2696 1701 2754 1739
rect 2696 1667 2708 1701
rect 2742 1667 2754 1701
rect 2696 1629 2754 1667
rect 2696 1595 2708 1629
rect 2742 1595 2754 1629
rect 2696 1557 2754 1595
rect 2696 1523 2708 1557
rect 2742 1523 2754 1557
rect 2696 1485 2754 1523
rect 2696 1451 2708 1485
rect 2742 1451 2754 1485
rect 2696 1413 2754 1451
rect 2696 1379 2708 1413
rect 2742 1379 2754 1413
rect 2696 1341 2754 1379
rect 2696 1307 2708 1341
rect 2742 1307 2754 1341
rect 2696 1269 2754 1307
rect 2696 1235 2708 1269
rect 2742 1235 2754 1269
rect 2696 1197 2754 1235
rect 2696 1163 2708 1197
rect 2742 1163 2754 1197
rect 2696 1125 2754 1163
rect 2696 1091 2708 1125
rect 2742 1091 2754 1125
rect 2696 1053 2754 1091
rect 2696 1019 2708 1053
rect 2742 1019 2754 1053
rect 2696 981 2754 1019
rect 2696 947 2708 981
rect 2742 947 2754 981
rect 2696 909 2754 947
rect 2696 875 2708 909
rect 2742 875 2754 909
rect 2696 837 2754 875
rect 2696 803 2708 837
rect 2742 803 2754 837
rect 2696 765 2754 803
rect 2696 731 2708 765
rect 2742 731 2754 765
rect 2696 693 2754 731
rect 2696 659 2708 693
rect 2742 659 2754 693
rect 2696 621 2754 659
rect 2696 587 2708 621
rect 2742 587 2754 621
rect 2696 549 2754 587
rect 2696 515 2708 549
rect 2742 515 2754 549
rect 2696 477 2754 515
rect 2696 443 2708 477
rect 2742 443 2754 477
rect 2696 405 2754 443
rect 2696 371 2708 405
rect 2742 371 2754 405
rect 2696 333 2754 371
rect 2696 299 2708 333
rect 2742 299 2754 333
rect 38 227 50 261
rect 84 227 96 261
rect 38 189 96 227
rect 38 155 50 189
rect 84 155 96 189
rect 38 96 96 155
rect 2696 261 2754 299
rect 2696 227 2708 261
rect 2742 227 2754 261
rect 2696 189 2754 227
rect 2696 155 2708 189
rect 2742 155 2754 189
rect 2696 96 2754 155
rect 38 84 2754 96
rect 38 50 50 84
rect 84 50 155 84
rect 189 50 227 84
rect 261 50 299 84
rect 333 50 371 84
rect 405 50 443 84
rect 477 50 515 84
rect 549 50 587 84
rect 621 50 659 84
rect 693 50 731 84
rect 765 50 803 84
rect 837 50 875 84
rect 909 50 947 84
rect 981 50 1019 84
rect 1053 50 1091 84
rect 1125 50 1163 84
rect 1197 50 1235 84
rect 1269 50 1307 84
rect 1341 50 1379 84
rect 1413 50 1451 84
rect 1485 50 1523 84
rect 1557 50 1595 84
rect 1629 50 1667 84
rect 1701 50 1739 84
rect 1773 50 1811 84
rect 1845 50 1883 84
rect 1917 50 1955 84
rect 1989 50 2027 84
rect 2061 50 2099 84
rect 2133 50 2171 84
rect 2205 50 2243 84
rect 2277 50 2315 84
rect 2349 50 2387 84
rect 2421 50 2459 84
rect 2493 50 2531 84
rect 2565 50 2603 84
rect 2637 50 2708 84
rect 2742 50 2754 84
rect 38 38 2754 50
<< properties >>
string GDS_END 9117514
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 9039998
string path 7.850 12.350 7.850 61.950 61.950 61.950 61.950 7.850 3.350 7.850 
<< end >>
