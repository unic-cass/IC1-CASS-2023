// This is the unpowered netlist.
module egd_top_wrapper (la_data_in_65,
    wb_clk_i,
    la_data_in_58_43,
    la_data_in_60_59,
    la_data_out_23_16,
    la_data_out_26_24,
    la_data_out_30_27);
 input la_data_in_65;
 input wb_clk_i;
 input [15:0] la_data_in_58_43;
 input [1:0] la_data_in_60_59;
 output [7:0] la_data_out_23_16;
 output [2:0] la_data_out_26_24;
 output [3:0] la_data_out_30_27;

 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire _3360_;
 wire _3361_;
 wire _3362_;
 wire _3363_;
 wire _3364_;
 wire _3365_;
 wire _3366_;
 wire _3367_;
 wire _3368_;
 wire _3369_;
 wire clknet_0__2913_;
 wire clknet_0__2914_;
 wire clknet_0__2915_;
 wire clknet_0__2916_;
 wire clknet_0__2917_;
 wire clknet_0__2918_;
 wire clknet_0__2919_;
 wire clknet_0__2920_;
 wire clknet_0__2921_;
 wire clknet_0__2922_;
 wire clknet_0__2923_;
 wire clknet_0__2924_;
 wire clknet_0__2925_;
 wire clknet_0__2926_;
 wire clknet_0__2927_;
 wire clknet_1_0__leaf__2913_;
 wire clknet_1_0__leaf__2914_;
 wire clknet_1_0__leaf__2915_;
 wire clknet_1_0__leaf__2916_;
 wire clknet_1_0__leaf__2917_;
 wire clknet_1_0__leaf__2918_;
 wire clknet_1_0__leaf__2919_;
 wire clknet_1_0__leaf__2920_;
 wire clknet_1_0__leaf__2921_;
 wire clknet_1_0__leaf__2922_;
 wire clknet_1_0__leaf__2923_;
 wire clknet_1_0__leaf__2924_;
 wire clknet_1_0__leaf__2925_;
 wire clknet_1_0__leaf__2926_;
 wire clknet_1_0__leaf__2927_;
 wire clknet_1_1__leaf__2913_;
 wire clknet_1_1__leaf__2914_;
 wire clknet_1_1__leaf__2915_;
 wire clknet_1_1__leaf__2916_;
 wire clknet_1_1__leaf__2917_;
 wire clknet_1_1__leaf__2918_;
 wire clknet_1_1__leaf__2919_;
 wire clknet_1_1__leaf__2920_;
 wire clknet_1_1__leaf__2921_;
 wire clknet_1_1__leaf__2922_;
 wire clknet_1_1__leaf__2923_;
 wire clknet_1_1__leaf__2924_;
 wire clknet_1_1__leaf__2925_;
 wire clknet_1_1__leaf__2926_;
 wire clknet_1_1__leaf__2927_;
 wire \egd_top.BitStream_buffer.BS_buffer[0] ;
 wire \egd_top.BitStream_buffer.BS_buffer[100] ;
 wire \egd_top.BitStream_buffer.BS_buffer[101] ;
 wire \egd_top.BitStream_buffer.BS_buffer[102] ;
 wire \egd_top.BitStream_buffer.BS_buffer[103] ;
 wire \egd_top.BitStream_buffer.BS_buffer[104] ;
 wire \egd_top.BitStream_buffer.BS_buffer[105] ;
 wire \egd_top.BitStream_buffer.BS_buffer[106] ;
 wire \egd_top.BitStream_buffer.BS_buffer[107] ;
 wire \egd_top.BitStream_buffer.BS_buffer[108] ;
 wire \egd_top.BitStream_buffer.BS_buffer[109] ;
 wire \egd_top.BitStream_buffer.BS_buffer[10] ;
 wire \egd_top.BitStream_buffer.BS_buffer[110] ;
 wire \egd_top.BitStream_buffer.BS_buffer[111] ;
 wire \egd_top.BitStream_buffer.BS_buffer[112] ;
 wire \egd_top.BitStream_buffer.BS_buffer[113] ;
 wire \egd_top.BitStream_buffer.BS_buffer[114] ;
 wire \egd_top.BitStream_buffer.BS_buffer[115] ;
 wire \egd_top.BitStream_buffer.BS_buffer[116] ;
 wire \egd_top.BitStream_buffer.BS_buffer[117] ;
 wire \egd_top.BitStream_buffer.BS_buffer[118] ;
 wire \egd_top.BitStream_buffer.BS_buffer[119] ;
 wire \egd_top.BitStream_buffer.BS_buffer[11] ;
 wire \egd_top.BitStream_buffer.BS_buffer[120] ;
 wire \egd_top.BitStream_buffer.BS_buffer[121] ;
 wire \egd_top.BitStream_buffer.BS_buffer[122] ;
 wire \egd_top.BitStream_buffer.BS_buffer[123] ;
 wire \egd_top.BitStream_buffer.BS_buffer[124] ;
 wire \egd_top.BitStream_buffer.BS_buffer[125] ;
 wire \egd_top.BitStream_buffer.BS_buffer[126] ;
 wire \egd_top.BitStream_buffer.BS_buffer[127] ;
 wire \egd_top.BitStream_buffer.BS_buffer[12] ;
 wire \egd_top.BitStream_buffer.BS_buffer[13] ;
 wire \egd_top.BitStream_buffer.BS_buffer[14] ;
 wire \egd_top.BitStream_buffer.BS_buffer[15] ;
 wire \egd_top.BitStream_buffer.BS_buffer[16] ;
 wire \egd_top.BitStream_buffer.BS_buffer[17] ;
 wire \egd_top.BitStream_buffer.BS_buffer[18] ;
 wire \egd_top.BitStream_buffer.BS_buffer[19] ;
 wire \egd_top.BitStream_buffer.BS_buffer[1] ;
 wire \egd_top.BitStream_buffer.BS_buffer[20] ;
 wire \egd_top.BitStream_buffer.BS_buffer[21] ;
 wire \egd_top.BitStream_buffer.BS_buffer[22] ;
 wire \egd_top.BitStream_buffer.BS_buffer[23] ;
 wire \egd_top.BitStream_buffer.BS_buffer[24] ;
 wire \egd_top.BitStream_buffer.BS_buffer[25] ;
 wire \egd_top.BitStream_buffer.BS_buffer[26] ;
 wire \egd_top.BitStream_buffer.BS_buffer[27] ;
 wire \egd_top.BitStream_buffer.BS_buffer[28] ;
 wire \egd_top.BitStream_buffer.BS_buffer[29] ;
 wire \egd_top.BitStream_buffer.BS_buffer[2] ;
 wire \egd_top.BitStream_buffer.BS_buffer[30] ;
 wire \egd_top.BitStream_buffer.BS_buffer[31] ;
 wire \egd_top.BitStream_buffer.BS_buffer[32] ;
 wire \egd_top.BitStream_buffer.BS_buffer[33] ;
 wire \egd_top.BitStream_buffer.BS_buffer[34] ;
 wire \egd_top.BitStream_buffer.BS_buffer[35] ;
 wire \egd_top.BitStream_buffer.BS_buffer[36] ;
 wire \egd_top.BitStream_buffer.BS_buffer[37] ;
 wire \egd_top.BitStream_buffer.BS_buffer[38] ;
 wire \egd_top.BitStream_buffer.BS_buffer[39] ;
 wire \egd_top.BitStream_buffer.BS_buffer[3] ;
 wire \egd_top.BitStream_buffer.BS_buffer[40] ;
 wire \egd_top.BitStream_buffer.BS_buffer[41] ;
 wire \egd_top.BitStream_buffer.BS_buffer[42] ;
 wire \egd_top.BitStream_buffer.BS_buffer[43] ;
 wire \egd_top.BitStream_buffer.BS_buffer[44] ;
 wire \egd_top.BitStream_buffer.BS_buffer[45] ;
 wire \egd_top.BitStream_buffer.BS_buffer[46] ;
 wire \egd_top.BitStream_buffer.BS_buffer[47] ;
 wire \egd_top.BitStream_buffer.BS_buffer[48] ;
 wire \egd_top.BitStream_buffer.BS_buffer[49] ;
 wire \egd_top.BitStream_buffer.BS_buffer[4] ;
 wire \egd_top.BitStream_buffer.BS_buffer[50] ;
 wire \egd_top.BitStream_buffer.BS_buffer[51] ;
 wire \egd_top.BitStream_buffer.BS_buffer[52] ;
 wire \egd_top.BitStream_buffer.BS_buffer[53] ;
 wire \egd_top.BitStream_buffer.BS_buffer[54] ;
 wire \egd_top.BitStream_buffer.BS_buffer[55] ;
 wire \egd_top.BitStream_buffer.BS_buffer[56] ;
 wire \egd_top.BitStream_buffer.BS_buffer[57] ;
 wire \egd_top.BitStream_buffer.BS_buffer[58] ;
 wire \egd_top.BitStream_buffer.BS_buffer[59] ;
 wire \egd_top.BitStream_buffer.BS_buffer[5] ;
 wire \egd_top.BitStream_buffer.BS_buffer[60] ;
 wire \egd_top.BitStream_buffer.BS_buffer[61] ;
 wire \egd_top.BitStream_buffer.BS_buffer[62] ;
 wire \egd_top.BitStream_buffer.BS_buffer[63] ;
 wire \egd_top.BitStream_buffer.BS_buffer[64] ;
 wire \egd_top.BitStream_buffer.BS_buffer[65] ;
 wire \egd_top.BitStream_buffer.BS_buffer[66] ;
 wire \egd_top.BitStream_buffer.BS_buffer[67] ;
 wire \egd_top.BitStream_buffer.BS_buffer[68] ;
 wire \egd_top.BitStream_buffer.BS_buffer[69] ;
 wire \egd_top.BitStream_buffer.BS_buffer[6] ;
 wire \egd_top.BitStream_buffer.BS_buffer[70] ;
 wire \egd_top.BitStream_buffer.BS_buffer[71] ;
 wire \egd_top.BitStream_buffer.BS_buffer[72] ;
 wire \egd_top.BitStream_buffer.BS_buffer[73] ;
 wire \egd_top.BitStream_buffer.BS_buffer[74] ;
 wire \egd_top.BitStream_buffer.BS_buffer[75] ;
 wire \egd_top.BitStream_buffer.BS_buffer[76] ;
 wire \egd_top.BitStream_buffer.BS_buffer[77] ;
 wire \egd_top.BitStream_buffer.BS_buffer[78] ;
 wire \egd_top.BitStream_buffer.BS_buffer[79] ;
 wire \egd_top.BitStream_buffer.BS_buffer[7] ;
 wire \egd_top.BitStream_buffer.BS_buffer[80] ;
 wire \egd_top.BitStream_buffer.BS_buffer[81] ;
 wire \egd_top.BitStream_buffer.BS_buffer[82] ;
 wire \egd_top.BitStream_buffer.BS_buffer[83] ;
 wire \egd_top.BitStream_buffer.BS_buffer[84] ;
 wire \egd_top.BitStream_buffer.BS_buffer[85] ;
 wire \egd_top.BitStream_buffer.BS_buffer[86] ;
 wire \egd_top.BitStream_buffer.BS_buffer[87] ;
 wire \egd_top.BitStream_buffer.BS_buffer[88] ;
 wire \egd_top.BitStream_buffer.BS_buffer[89] ;
 wire \egd_top.BitStream_buffer.BS_buffer[8] ;
 wire \egd_top.BitStream_buffer.BS_buffer[90] ;
 wire \egd_top.BitStream_buffer.BS_buffer[91] ;
 wire \egd_top.BitStream_buffer.BS_buffer[92] ;
 wire \egd_top.BitStream_buffer.BS_buffer[93] ;
 wire \egd_top.BitStream_buffer.BS_buffer[94] ;
 wire \egd_top.BitStream_buffer.BS_buffer[95] ;
 wire \egd_top.BitStream_buffer.BS_buffer[96] ;
 wire \egd_top.BitStream_buffer.BS_buffer[97] ;
 wire \egd_top.BitStream_buffer.BS_buffer[98] ;
 wire \egd_top.BitStream_buffer.BS_buffer[99] ;
 wire \egd_top.BitStream_buffer.BS_buffer[9] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[10] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[11] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[12] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[13] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[14] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[15] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[1] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[2] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[3] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[4] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[5] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[6] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[7] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[8] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[9] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_valid_n ;
 wire \egd_top.BitStream_buffer.buffer_index[4] ;
 wire \egd_top.BitStream_buffer.buffer_index[5] ;
 wire \egd_top.BitStream_buffer.buffer_index[6] ;
 wire \egd_top.BitStream_buffer.exp_golomb_len[1] ;
 wire \egd_top.BitStream_buffer.exp_golomb_len[2] ;
 wire \egd_top.BitStream_buffer.exp_golomb_len[3] ;
 wire \egd_top.BitStream_buffer.pc[1] ;
 wire \egd_top.BitStream_buffer.pc[2] ;
 wire \egd_top.BitStream_buffer.pc[3] ;
 wire \egd_top.BitStream_buffer.pc[4] ;
 wire \egd_top.BitStream_buffer.pc[5] ;
 wire \egd_top.BitStream_buffer.pc[6] ;
 wire \egd_top.BitStream_buffer.pc_previous[0] ;
 wire \egd_top.BitStream_buffer.pc_previous[1] ;
 wire \egd_top.BitStream_buffer.pc_previous[2] ;
 wire \egd_top.BitStream_buffer.pc_previous[3] ;
 wire \egd_top.BitStream_buffer.pc_previous[4] ;
 wire \egd_top.BitStream_buffer.pc_previous[5] ;
 wire \egd_top.BitStream_buffer.pc_previous[6] ;
 wire \egd_top.exp_golomb_decoding.te_range[2] ;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_1217_));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(_1447_));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_1635_));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_1692_));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_1814_));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(_2369_));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(net5));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_191 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_198 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_357 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_538 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_214 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_228 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_553 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_254 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_554 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_280 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_46 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_491 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_471 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_479 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_504 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_140 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_466 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_79 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_67 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_228 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_410 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_471 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_507 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_554 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_79 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_79 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_495 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_552 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_331 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_59 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_508 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_423 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_60 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_527 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_532 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_224 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_366 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_536 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_76 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_451 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_519 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_413 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_394 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_310 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_200 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_168 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_534 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_394 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_536 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_476 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_536 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_140 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_254 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_366 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_480 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_479 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_504 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_367 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_482 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_133 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_370 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_535 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_476 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_507 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_469 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_535 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_410 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_422 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_396 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_424 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_107 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_392 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_396 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_480 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_186 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_469 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_424 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_451 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_275 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_327 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_394 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_92 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__inv_2 _3370_ (.A(net33),
    .Y(_2928_));
 sky130_fd_sc_hd__nand2_1 _3371_ (.A(net32),
    .B(net31),
    .Y(_2929_));
 sky130_fd_sc_hd__inv_2 _3372_ (.A(net34),
    .Y(_2930_));
 sky130_fd_sc_hd__o21ai_1 _3373_ (.A1(_2928_),
    .A2(_2929_),
    .B1(_2930_),
    .Y(_2931_));
 sky130_fd_sc_hd__buf_6 _3374_ (.A(net19),
    .X(_2932_));
 sky130_fd_sc_hd__buf_2 _3375_ (.A(_2932_),
    .X(_2933_));
 sky130_fd_sc_hd__and2_1 _3376_ (.A(_2931_),
    .B(_2933_),
    .X(_2934_));
 sky130_fd_sc_hd__clkbuf_1 _3377_ (.A(_2934_),
    .X(_0321_));
 sky130_fd_sc_hd__a21o_1 _3378_ (.A1(_2928_),
    .A2(_2929_),
    .B1(_2931_),
    .X(_2935_));
 sky130_fd_sc_hd__nand2_1 _3379_ (.A(net34),
    .B(net33),
    .Y(_2936_));
 sky130_fd_sc_hd__inv_2 _3380_ (.A(_2932_),
    .Y(_2937_));
 sky130_fd_sc_hd__clkbuf_4 _3381_ (.A(_2937_),
    .X(_2938_));
 sky130_fd_sc_hd__a21oi_1 _3382_ (.A1(_2935_),
    .A2(_2936_),
    .B1(_2938_),
    .Y(_0320_));
 sky130_fd_sc_hd__inv_2 _3383_ (.A(net31),
    .Y(_2939_));
 sky130_fd_sc_hd__nor2_1 _3384_ (.A(net33),
    .B(net32),
    .Y(_2940_));
 sky130_fd_sc_hd__nor2_1 _3385_ (.A(_2930_),
    .B(_2940_),
    .Y(_2941_));
 sky130_fd_sc_hd__nor2_1 _3386_ (.A(_2939_),
    .B(_2941_),
    .Y(_2942_));
 sky130_fd_sc_hd__a21o_1 _3387_ (.A1(_2942_),
    .A2(net32),
    .B1(_2937_),
    .X(_2943_));
 sky130_fd_sc_hd__o21ba_1 _3388_ (.A1(net32),
    .A2(_2942_),
    .B1_N(_2943_),
    .X(_2944_));
 sky130_fd_sc_hd__clkbuf_1 _3389_ (.A(_2944_),
    .X(_0319_));
 sky130_fd_sc_hd__inv_2 _3390_ (.A(_2941_),
    .Y(_2945_));
 sky130_fd_sc_hd__nor2_1 _3391_ (.A(net31),
    .B(_2945_),
    .Y(_2946_));
 sky130_fd_sc_hd__or3_1 _3392_ (.A(_2937_),
    .B(_2942_),
    .C(_2946_),
    .X(_2947_));
 sky130_fd_sc_hd__inv_2 _3393_ (.A(_2947_),
    .Y(_0318_));
 sky130_fd_sc_hd__inv_2 _3394_ (.A(net30),
    .Y(_2948_));
 sky130_fd_sc_hd__nor2_1 _3395_ (.A(net29),
    .B(net28),
    .Y(_2949_));
 sky130_fd_sc_hd__nor2_1 _3396_ (.A(_2948_),
    .B(_2949_),
    .Y(_2950_));
 sky130_fd_sc_hd__a21o_1 _3397_ (.A1(net29),
    .A2(net28),
    .B1(net30),
    .X(_2951_));
 sky130_fd_sc_hd__and2b_1 _3398_ (.A_N(_2950_),
    .B(_2951_),
    .X(_2952_));
 sky130_fd_sc_hd__inv_2 _3399_ (.A(net29),
    .Y(_2953_));
 sky130_fd_sc_hd__nand2_4 _3400_ (.A(\egd_top.BitStream_buffer.pc[2] ),
    .B(\egd_top.BitStream_buffer.pc[3] ),
    .Y(_2954_));
 sky130_fd_sc_hd__inv_2 _3401_ (.A(net18),
    .Y(_2955_));
 sky130_fd_sc_hd__inv_2 _3402_ (.A(net17),
    .Y(_2956_));
 sky130_fd_sc_hd__nand2_1 _3403_ (.A(_2955_),
    .B(_2956_),
    .Y(_2957_));
 sky130_fd_sc_hd__or2_1 _3404_ (.A(\egd_top.BitStream_buffer.pc_previous[0] ),
    .B(_2957_),
    .X(_2958_));
 sky130_fd_sc_hd__buf_6 _3405_ (.A(_2957_),
    .X(_2959_));
 sky130_fd_sc_hd__nand2_4 _3406_ (.A(_2959_),
    .B(\egd_top.BitStream_buffer.pc_previous[0] ),
    .Y(_2960_));
 sky130_fd_sc_hd__nand2_2 _3407_ (.A(_2958_),
    .B(_2960_),
    .Y(_2961_));
 sky130_fd_sc_hd__inv_2 _3408_ (.A(_2961_),
    .Y(_2962_));
 sky130_fd_sc_hd__nand2_2 _3409_ (.A(_2962_),
    .B(\egd_top.BitStream_buffer.pc[1] ),
    .Y(_2963_));
 sky130_fd_sc_hd__nor2_2 _3410_ (.A(_2954_),
    .B(_2963_),
    .Y(_2964_));
 sky130_fd_sc_hd__inv_2 _3411_ (.A(\egd_top.BitStream_buffer.pc[6] ),
    .Y(_2965_));
 sky130_fd_sc_hd__and3_1 _3412_ (.A(_2965_),
    .B(\egd_top.BitStream_buffer.pc[4] ),
    .C(\egd_top.BitStream_buffer.pc[5] ),
    .X(_2966_));
 sky130_fd_sc_hd__and2_1 _3413_ (.A(_2964_),
    .B(_2966_),
    .X(_2967_));
 sky130_fd_sc_hd__nor2_1 _3414_ (.A(\egd_top.BitStream_buffer.pc[6] ),
    .B(_2967_),
    .Y(_2968_));
 sky130_fd_sc_hd__inv_2 _3415_ (.A(_2949_),
    .Y(_2969_));
 sky130_fd_sc_hd__nor2_1 _3416_ (.A(net30),
    .B(_2969_),
    .Y(_2970_));
 sky130_fd_sc_hd__inv_2 _3417_ (.A(net198),
    .Y(_2971_));
 sky130_fd_sc_hd__inv_2 _3418_ (.A(net196),
    .Y(_2972_));
 sky130_fd_sc_hd__and3_2 _3419_ (.A(_2971_),
    .B(_2972_),
    .C(net200),
    .X(_2973_));
 sky130_fd_sc_hd__nand3_1 _3420_ (.A(_2968_),
    .B(_2970_),
    .C(_2973_),
    .Y(_2974_));
 sky130_fd_sc_hd__nor2_1 _3421_ (.A(_2950_),
    .B(_2970_),
    .Y(_2975_));
 sky130_fd_sc_hd__inv_2 _3422_ (.A(_2975_),
    .Y(_2976_));
 sky130_fd_sc_hd__nand2_1 _3423_ (.A(_2974_),
    .B(_2976_),
    .Y(_2977_));
 sky130_fd_sc_hd__inv_2 _3424_ (.A(net200),
    .Y(_2978_));
 sky130_fd_sc_hd__and3_2 _3425_ (.A(_2978_),
    .B(_2971_),
    .C(_2972_),
    .X(_2979_));
 sky130_fd_sc_hd__and4_1 _3426_ (.A(\egd_top.BitStream_buffer.pc_previous[0] ),
    .B(\egd_top.BitStream_buffer.pc_previous[1] ),
    .C(\egd_top.BitStream_buffer.pc_previous[2] ),
    .D(\egd_top.BitStream_buffer.pc_previous[3] ),
    .X(_2980_));
 sky130_fd_sc_hd__a31o_1 _3427_ (.A1(_2980_),
    .A2(\egd_top.BitStream_buffer.pc_previous[4] ),
    .A3(\egd_top.BitStream_buffer.pc_previous[5] ),
    .B1(\egd_top.BitStream_buffer.pc_previous[6] ),
    .X(_2981_));
 sky130_fd_sc_hd__nand2_1 _3428_ (.A(_2968_),
    .B(_2981_),
    .Y(_2982_));
 sky130_fd_sc_hd__or2_1 _3429_ (.A(\egd_top.BitStream_buffer.pc_previous[6] ),
    .B(_2965_),
    .X(_2983_));
 sky130_fd_sc_hd__a21boi_1 _3430_ (.A1(_2982_),
    .A2(_2983_),
    .B1_N(_2970_),
    .Y(_2984_));
 sky130_fd_sc_hd__a31o_1 _3431_ (.A1(\egd_top.BitStream_buffer.pc[6] ),
    .A2(_2970_),
    .A3(_2979_),
    .B1(_2984_),
    .X(_2985_));
 sky130_fd_sc_hd__a311o_1 _3432_ (.A1(net30),
    .A2(_2953_),
    .A3(net28),
    .B1(_2977_),
    .C1(_2985_),
    .X(_2986_));
 sky130_fd_sc_hd__and4_1 _3433_ (.A(_2928_),
    .B(_2939_),
    .C(net34),
    .D(net32),
    .X(_2987_));
 sky130_fd_sc_hd__nand2_2 _3434_ (.A(_2986_),
    .B(_2987_),
    .Y(_2988_));
 sky130_fd_sc_hd__clkbuf_4 _3435_ (.A(_2932_),
    .X(_2989_));
 sky130_fd_sc_hd__nand2_1 _3436_ (.A(_2988_),
    .B(_2948_),
    .Y(_2990_));
 sky130_fd_sc_hd__o211a_1 _3437_ (.A1(_2952_),
    .A2(_2988_),
    .B1(_2989_),
    .C1(_2990_),
    .X(_0317_));
 sky130_fd_sc_hd__nor2_1 _3438_ (.A(_2949_),
    .B(_2951_),
    .Y(_2991_));
 sky130_fd_sc_hd__nand2_1 _3439_ (.A(_2988_),
    .B(_2953_),
    .Y(_2992_));
 sky130_fd_sc_hd__o211a_1 _3440_ (.A1(_2991_),
    .A2(_2988_),
    .B1(_2989_),
    .C1(_2992_),
    .X(_0316_));
 sky130_fd_sc_hd__o21ai_1 _3441_ (.A1(net28),
    .A2(_2976_),
    .B1(_2974_),
    .Y(_2993_));
 sky130_fd_sc_hd__o21bai_1 _3442_ (.A1(_2985_),
    .A2(_2993_),
    .B1_N(_2988_),
    .Y(_2994_));
 sky130_fd_sc_hd__nand2_1 _3443_ (.A(_2988_),
    .B(net28),
    .Y(_2995_));
 sky130_fd_sc_hd__a21oi_1 _3444_ (.A1(_2994_),
    .A2(_2995_),
    .B1(_2938_),
    .Y(_0315_));
 sky130_fd_sc_hd__buf_2 _3445_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_valid_n ),
    .X(_2996_));
 sky130_fd_sc_hd__inv_2 _3446_ (.A(_2996_),
    .Y(_2997_));
 sky130_fd_sc_hd__o21ai_1 _3447_ (.A1(_2997_),
    .A2(_2987_),
    .B1(_2989_),
    .Y(_0314_));
 sky130_fd_sc_hd__clkbuf_4 _3448_ (.A(\egd_top.BitStream_buffer.BS_buffer[112] ),
    .X(_2998_));
 sky130_fd_sc_hd__nand2_1 _3449_ (.A(_2948_),
    .B(_2953_),
    .Y(_2999_));
 sky130_fd_sc_hd__nand2_1 _3450_ (.A(net30),
    .B(net29),
    .Y(_3000_));
 sky130_fd_sc_hd__nand2_1 _3451_ (.A(_2940_),
    .B(_2930_),
    .Y(_3001_));
 sky130_fd_sc_hd__a22o_4 _3452_ (.A1(_2999_),
    .A2(_3000_),
    .B1(_2945_),
    .B2(_3001_),
    .X(_3002_));
 sky130_fd_sc_hd__nand2_1 _3453_ (.A(_3002_),
    .B(net201),
    .Y(_3003_));
 sky130_fd_sc_hd__or2_1 _3454_ (.A(_2971_),
    .B(_3003_),
    .X(_3004_));
 sky130_fd_sc_hd__or2_1 _3455_ (.A(_2978_),
    .B(_3004_),
    .X(_3005_));
 sky130_fd_sc_hd__buf_2 _3456_ (.A(_3005_),
    .X(_3006_));
 sky130_fd_sc_hd__buf_4 _3457_ (.A(_3006_),
    .X(_3007_));
 sky130_fd_sc_hd__mux2_1 _3458_ (.A0(net7),
    .A1(_2998_),
    .S(_3007_),
    .X(_3008_));
 sky130_fd_sc_hd__and2_1 _3459_ (.A(_3008_),
    .B(_2933_),
    .X(_3009_));
 sky130_fd_sc_hd__clkbuf_1 _3460_ (.A(_3009_),
    .X(_0313_));
 sky130_fd_sc_hd__clkbuf_4 _3461_ (.A(\egd_top.BitStream_buffer.BS_buffer[113] ),
    .X(_3010_));
 sky130_fd_sc_hd__mux2_1 _3462_ (.A0(net6),
    .A1(_3010_),
    .S(_3007_),
    .X(_3011_));
 sky130_fd_sc_hd__and2_1 _3463_ (.A(_3011_),
    .B(_2933_),
    .X(_3012_));
 sky130_fd_sc_hd__clkbuf_1 _3464_ (.A(_3012_),
    .X(_0312_));
 sky130_fd_sc_hd__clkbuf_4 _3465_ (.A(\egd_top.BitStream_buffer.BS_buffer[114] ),
    .X(_3013_));
 sky130_fd_sc_hd__mux2_1 _3466_ (.A0(net5),
    .A1(_3013_),
    .S(_3007_),
    .X(_3014_));
 sky130_fd_sc_hd__and2_1 _3467_ (.A(_3014_),
    .B(_2933_),
    .X(_3015_));
 sky130_fd_sc_hd__clkbuf_1 _3468_ (.A(_3015_),
    .X(_0311_));
 sky130_fd_sc_hd__clkbuf_4 _3469_ (.A(\egd_top.BitStream_buffer.BS_buffer[115] ),
    .X(_3016_));
 sky130_fd_sc_hd__mux2_1 _3470_ (.A0(net4),
    .A1(_3016_),
    .S(_3007_),
    .X(_3017_));
 sky130_fd_sc_hd__and2_1 _3471_ (.A(_3017_),
    .B(_2933_),
    .X(_3018_));
 sky130_fd_sc_hd__clkbuf_1 _3472_ (.A(_3018_),
    .X(_0310_));
 sky130_fd_sc_hd__clkbuf_4 _3473_ (.A(\egd_top.BitStream_buffer.BS_buffer[116] ),
    .X(_3019_));
 sky130_fd_sc_hd__mux2_1 _3474_ (.A0(net3),
    .A1(_3019_),
    .S(_3007_),
    .X(_3020_));
 sky130_fd_sc_hd__and2_1 _3475_ (.A(_3020_),
    .B(_2933_),
    .X(_3021_));
 sky130_fd_sc_hd__clkbuf_1 _3476_ (.A(_3021_),
    .X(_0309_));
 sky130_fd_sc_hd__clkbuf_4 _3477_ (.A(\egd_top.BitStream_buffer.BS_buffer[117] ),
    .X(_3022_));
 sky130_fd_sc_hd__mux2_1 _3478_ (.A0(net2),
    .A1(_3022_),
    .S(_3007_),
    .X(_3023_));
 sky130_fd_sc_hd__and2_1 _3479_ (.A(_3023_),
    .B(_2933_),
    .X(_3024_));
 sky130_fd_sc_hd__clkbuf_1 _3480_ (.A(_3024_),
    .X(_0308_));
 sky130_fd_sc_hd__clkbuf_4 _3481_ (.A(\egd_top.BitStream_buffer.BS_buffer[118] ),
    .X(_3025_));
 sky130_fd_sc_hd__mux2_1 _3482_ (.A0(net16),
    .A1(_3025_),
    .S(_3007_),
    .X(_3026_));
 sky130_fd_sc_hd__and2_1 _3483_ (.A(_3026_),
    .B(_2933_),
    .X(_3027_));
 sky130_fd_sc_hd__clkbuf_1 _3484_ (.A(_3027_),
    .X(_0307_));
 sky130_fd_sc_hd__clkbuf_4 _3485_ (.A(\egd_top.BitStream_buffer.BS_buffer[119] ),
    .X(_3028_));
 sky130_fd_sc_hd__mux2_1 _3486_ (.A0(net15),
    .A1(_3028_),
    .S(_3007_),
    .X(_3029_));
 sky130_fd_sc_hd__and2_1 _3487_ (.A(_3029_),
    .B(_2933_),
    .X(_3030_));
 sky130_fd_sc_hd__clkbuf_1 _3488_ (.A(_3030_),
    .X(_0306_));
 sky130_fd_sc_hd__clkbuf_4 _3489_ (.A(\egd_top.BitStream_buffer.BS_buffer[120] ),
    .X(_3031_));
 sky130_fd_sc_hd__mux2_1 _3490_ (.A0(net14),
    .A1(_3031_),
    .S(_3007_),
    .X(_3032_));
 sky130_fd_sc_hd__and2_1 _3491_ (.A(_3032_),
    .B(_2933_),
    .X(_3033_));
 sky130_fd_sc_hd__clkbuf_1 _3492_ (.A(_3033_),
    .X(_0305_));
 sky130_fd_sc_hd__clkbuf_4 _3493_ (.A(\egd_top.BitStream_buffer.BS_buffer[121] ),
    .X(_3034_));
 sky130_fd_sc_hd__mux2_1 _3494_ (.A0(net13),
    .A1(_3034_),
    .S(_3007_),
    .X(_3035_));
 sky130_fd_sc_hd__and2_1 _3495_ (.A(_3035_),
    .B(_2933_),
    .X(_3036_));
 sky130_fd_sc_hd__clkbuf_1 _3496_ (.A(_3036_),
    .X(_0304_));
 sky130_fd_sc_hd__clkbuf_4 _3497_ (.A(\egd_top.BitStream_buffer.BS_buffer[122] ),
    .X(_3037_));
 sky130_fd_sc_hd__mux2_1 _3498_ (.A0(net12),
    .A1(_3037_),
    .S(_3007_),
    .X(_3038_));
 sky130_fd_sc_hd__and2_1 _3499_ (.A(_3038_),
    .B(_2933_),
    .X(_3039_));
 sky130_fd_sc_hd__clkbuf_1 _3500_ (.A(_3039_),
    .X(_0303_));
 sky130_fd_sc_hd__clkbuf_4 _3501_ (.A(\egd_top.BitStream_buffer.BS_buffer[123] ),
    .X(_3040_));
 sky130_fd_sc_hd__mux2_1 _3502_ (.A0(net11),
    .A1(_3040_),
    .S(_3006_),
    .X(_3041_));
 sky130_fd_sc_hd__buf_2 _3503_ (.A(_2932_),
    .X(_3042_));
 sky130_fd_sc_hd__and2_1 _3504_ (.A(_3041_),
    .B(_3042_),
    .X(_3043_));
 sky130_fd_sc_hd__clkbuf_1 _3505_ (.A(_3043_),
    .X(_0302_));
 sky130_fd_sc_hd__clkbuf_4 _3506_ (.A(\egd_top.BitStream_buffer.BS_buffer[124] ),
    .X(_3044_));
 sky130_fd_sc_hd__mux2_1 _3507_ (.A0(net10),
    .A1(_3044_),
    .S(_3006_),
    .X(_3045_));
 sky130_fd_sc_hd__and2_1 _3508_ (.A(_3045_),
    .B(_3042_),
    .X(_3046_));
 sky130_fd_sc_hd__clkbuf_1 _3509_ (.A(_3046_),
    .X(_0301_));
 sky130_fd_sc_hd__clkbuf_4 _3510_ (.A(\egd_top.BitStream_buffer.BS_buffer[125] ),
    .X(_3047_));
 sky130_fd_sc_hd__mux2_1 _3511_ (.A0(net9),
    .A1(_3047_),
    .S(_3006_),
    .X(_3048_));
 sky130_fd_sc_hd__and2_1 _3512_ (.A(_3048_),
    .B(_3042_),
    .X(_3049_));
 sky130_fd_sc_hd__clkbuf_1 _3513_ (.A(_3049_),
    .X(_0300_));
 sky130_fd_sc_hd__clkbuf_4 _3514_ (.A(\egd_top.BitStream_buffer.BS_buffer[126] ),
    .X(_3050_));
 sky130_fd_sc_hd__mux2_1 _3515_ (.A0(net8),
    .A1(_3050_),
    .S(_3006_),
    .X(_3051_));
 sky130_fd_sc_hd__and2_1 _3516_ (.A(_3051_),
    .B(_3042_),
    .X(_3052_));
 sky130_fd_sc_hd__clkbuf_1 _3517_ (.A(_3052_),
    .X(_0299_));
 sky130_fd_sc_hd__clkbuf_4 _3518_ (.A(\egd_top.BitStream_buffer.BS_buffer[127] ),
    .X(_3053_));
 sky130_fd_sc_hd__mux2_1 _3519_ (.A0(net1),
    .A1(_3053_),
    .S(_3006_),
    .X(_3054_));
 sky130_fd_sc_hd__and2_1 _3520_ (.A(_3054_),
    .B(_3042_),
    .X(_3055_));
 sky130_fd_sc_hd__clkbuf_1 _3521_ (.A(_3055_),
    .X(_0298_));
 sky130_fd_sc_hd__clkbuf_4 _3522_ (.A(_2996_),
    .X(_3056_));
 sky130_fd_sc_hd__clkbuf_4 _3523_ (.A(\egd_top.BitStream_buffer.BS_buffer[74] ),
    .X(_3057_));
 sky130_fd_sc_hd__nand2_2 _3524_ (.A(_2961_),
    .B(\egd_top.BitStream_buffer.pc[1] ),
    .Y(_3058_));
 sky130_fd_sc_hd__inv_2 _3525_ (.A(_3058_),
    .Y(_3059_));
 sky130_fd_sc_hd__inv_2 _3526_ (.A(\egd_top.BitStream_buffer.pc[2] ),
    .Y(_3060_));
 sky130_fd_sc_hd__and3_4 _3527_ (.A(_3059_),
    .B(_3060_),
    .C(\egd_top.BitStream_buffer.pc[3] ),
    .X(_3061_));
 sky130_fd_sc_hd__inv_2 _3528_ (.A(\egd_top.BitStream_buffer.pc[4] ),
    .Y(_3062_));
 sky130_fd_sc_hd__inv_2 _3529_ (.A(\egd_top.BitStream_buffer.pc[5] ),
    .Y(_3063_));
 sky130_fd_sc_hd__and3_1 _3530_ (.A(_3062_),
    .B(_3063_),
    .C(\egd_top.BitStream_buffer.pc[6] ),
    .X(_3064_));
 sky130_fd_sc_hd__buf_2 _3531_ (.A(_3064_),
    .X(_3065_));
 sky130_fd_sc_hd__and2_1 _3532_ (.A(_3061_),
    .B(_3065_),
    .X(_3066_));
 sky130_fd_sc_hd__buf_1 _3533_ (.A(_3066_),
    .X(_3067_));
 sky130_fd_sc_hd__clkbuf_4 _3534_ (.A(_3067_),
    .X(_3068_));
 sky130_fd_sc_hd__clkbuf_4 _3535_ (.A(\egd_top.BitStream_buffer.BS_buffer[75] ),
    .X(_3069_));
 sky130_fd_sc_hd__inv_2 _3536_ (.A(_2963_),
    .Y(_3070_));
 sky130_fd_sc_hd__and3_1 _3537_ (.A(_3070_),
    .B(_3060_),
    .C(\egd_top.BitStream_buffer.pc[3] ),
    .X(_3071_));
 sky130_fd_sc_hd__buf_2 _3538_ (.A(_3071_),
    .X(_3072_));
 sky130_fd_sc_hd__and2_1 _3539_ (.A(_3072_),
    .B(_3065_),
    .X(_3073_));
 sky130_fd_sc_hd__buf_1 _3540_ (.A(_3073_),
    .X(_3074_));
 sky130_fd_sc_hd__buf_4 _3541_ (.A(_3074_),
    .X(_3075_));
 sky130_fd_sc_hd__clkbuf_4 _3542_ (.A(\egd_top.BitStream_buffer.BS_buffer[72] ),
    .X(_3076_));
 sky130_fd_sc_hd__inv_2 _3543_ (.A(_3076_),
    .Y(_3077_));
 sky130_fd_sc_hd__inv_2 _3544_ (.A(\egd_top.BitStream_buffer.pc[1] ),
    .Y(_3078_));
 sky130_fd_sc_hd__nand2_2 _3545_ (.A(_2961_),
    .B(_3078_),
    .Y(_3079_));
 sky130_fd_sc_hd__inv_2 _3546_ (.A(_3079_),
    .Y(_3080_));
 sky130_fd_sc_hd__and3_1 _3547_ (.A(_3080_),
    .B(_3060_),
    .C(\egd_top.BitStream_buffer.pc[3] ),
    .X(_3081_));
 sky130_fd_sc_hd__clkbuf_4 _3548_ (.A(_3081_),
    .X(_3082_));
 sky130_fd_sc_hd__nand2_1 _3549_ (.A(_3082_),
    .B(_3065_),
    .Y(_3083_));
 sky130_fd_sc_hd__clkbuf_4 _3550_ (.A(_3083_),
    .X(_3084_));
 sky130_fd_sc_hd__clkbuf_4 _3551_ (.A(\egd_top.BitStream_buffer.BS_buffer[73] ),
    .X(_3085_));
 sky130_fd_sc_hd__inv_2 _3552_ (.A(_3085_),
    .Y(_3086_));
 sky130_fd_sc_hd__nand2_2 _3553_ (.A(_2962_),
    .B(_3078_),
    .Y(_3087_));
 sky130_fd_sc_hd__inv_2 _3554_ (.A(_3087_),
    .Y(_3088_));
 sky130_fd_sc_hd__and3_1 _3555_ (.A(_3088_),
    .B(_3060_),
    .C(\egd_top.BitStream_buffer.pc[3] ),
    .X(_3089_));
 sky130_fd_sc_hd__clkbuf_4 _3556_ (.A(_3089_),
    .X(_3090_));
 sky130_fd_sc_hd__nand2_1 _3557_ (.A(_3090_),
    .B(_3065_),
    .Y(_3091_));
 sky130_fd_sc_hd__clkbuf_4 _3558_ (.A(_3091_),
    .X(_3092_));
 sky130_fd_sc_hd__o22ai_1 _3559_ (.A1(_3077_),
    .A2(_3084_),
    .B1(_3086_),
    .B2(_3092_),
    .Y(_3093_));
 sky130_fd_sc_hd__a221oi_1 _3560_ (.A1(_3057_),
    .A2(_3068_),
    .B1(_3069_),
    .B2(_3075_),
    .C1(_3093_),
    .Y(_3094_));
 sky130_fd_sc_hd__clkbuf_4 _3561_ (.A(\egd_top.BitStream_buffer.BS_buffer[66] ),
    .X(_3095_));
 sky130_fd_sc_hd__inv_2 _3562_ (.A(\egd_top.BitStream_buffer.pc[3] ),
    .Y(_3096_));
 sky130_fd_sc_hd__nand2_4 _3563_ (.A(_3060_),
    .B(_3096_),
    .Y(_3097_));
 sky130_fd_sc_hd__nor2_4 _3564_ (.A(_3097_),
    .B(_3058_),
    .Y(_3098_));
 sky130_fd_sc_hd__and2_1 _3565_ (.A(_3098_),
    .B(_3064_),
    .X(_3099_));
 sky130_fd_sc_hd__buf_1 _3566_ (.A(_3099_),
    .X(_3100_));
 sky130_fd_sc_hd__clkbuf_4 _3567_ (.A(_3100_),
    .X(_3101_));
 sky130_fd_sc_hd__clkbuf_4 _3568_ (.A(\egd_top.BitStream_buffer.BS_buffer[67] ),
    .X(_3102_));
 sky130_fd_sc_hd__nor2_4 _3569_ (.A(_3097_),
    .B(_2963_),
    .Y(_3103_));
 sky130_fd_sc_hd__and2_1 _3570_ (.A(_3103_),
    .B(_3065_),
    .X(_3104_));
 sky130_fd_sc_hd__buf_1 _3571_ (.A(_3104_),
    .X(_3105_));
 sky130_fd_sc_hd__clkbuf_4 _3572_ (.A(_3105_),
    .X(_3106_));
 sky130_fd_sc_hd__clkbuf_4 _3573_ (.A(\egd_top.BitStream_buffer.BS_buffer[64] ),
    .X(_3107_));
 sky130_fd_sc_hd__inv_2 _3574_ (.A(_3107_),
    .Y(_3108_));
 sky130_fd_sc_hd__nor2_4 _3575_ (.A(_3097_),
    .B(_3079_),
    .Y(_3109_));
 sky130_fd_sc_hd__nand2_1 _3576_ (.A(_3109_),
    .B(_3065_),
    .Y(_3110_));
 sky130_fd_sc_hd__clkbuf_4 _3577_ (.A(_3110_),
    .X(_3111_));
 sky130_fd_sc_hd__nor2_2 _3578_ (.A(_3097_),
    .B(_3087_),
    .Y(_3112_));
 sky130_fd_sc_hd__and2_1 _3579_ (.A(_3112_),
    .B(_3065_),
    .X(_3113_));
 sky130_fd_sc_hd__clkbuf_4 _3580_ (.A(_3113_),
    .X(_3114_));
 sky130_fd_sc_hd__clkbuf_4 _3581_ (.A(\egd_top.BitStream_buffer.BS_buffer[65] ),
    .X(_3115_));
 sky130_fd_sc_hd__nand2_1 _3582_ (.A(_3114_),
    .B(_3115_),
    .Y(_3116_));
 sky130_fd_sc_hd__o21ai_1 _3583_ (.A1(_3108_),
    .A2(_3111_),
    .B1(_3116_),
    .Y(_3117_));
 sky130_fd_sc_hd__a221oi_1 _3584_ (.A1(_3095_),
    .A2(_3101_),
    .B1(_3102_),
    .B2(_3106_),
    .C1(_3117_),
    .Y(_3118_));
 sky130_fd_sc_hd__clkbuf_4 _3585_ (.A(\egd_top.BitStream_buffer.BS_buffer[71] ),
    .X(_3119_));
 sky130_fd_sc_hd__inv_2 _3586_ (.A(_3119_),
    .Y(_3120_));
 sky130_fd_sc_hd__and3_1 _3587_ (.A(_3070_),
    .B(\egd_top.BitStream_buffer.pc[2] ),
    .C(_3096_),
    .X(_3121_));
 sky130_fd_sc_hd__clkbuf_4 _3588_ (.A(_3121_),
    .X(_3122_));
 sky130_fd_sc_hd__nand2_1 _3589_ (.A(_3122_),
    .B(_3065_),
    .Y(_3123_));
 sky130_fd_sc_hd__clkbuf_4 _3590_ (.A(_3123_),
    .X(_3124_));
 sky130_fd_sc_hd__and3_1 _3591_ (.A(_3080_),
    .B(\egd_top.BitStream_buffer.pc[2] ),
    .C(_3096_),
    .X(_3125_));
 sky130_fd_sc_hd__clkbuf_4 _3592_ (.A(_3125_),
    .X(_3126_));
 sky130_fd_sc_hd__and2_1 _3593_ (.A(_3126_),
    .B(_3065_),
    .X(_3127_));
 sky130_fd_sc_hd__clkbuf_4 _3594_ (.A(_3127_),
    .X(_3128_));
 sky130_fd_sc_hd__clkbuf_4 _3595_ (.A(\egd_top.BitStream_buffer.BS_buffer[68] ),
    .X(_3129_));
 sky130_fd_sc_hd__nand2_1 _3596_ (.A(_3128_),
    .B(_3129_),
    .Y(_3130_));
 sky130_fd_sc_hd__and3_4 _3597_ (.A(_3059_),
    .B(\egd_top.BitStream_buffer.pc[2] ),
    .C(_3096_),
    .X(_3131_));
 sky130_fd_sc_hd__and2_1 _3598_ (.A(_3131_),
    .B(_3065_),
    .X(_3132_));
 sky130_fd_sc_hd__clkbuf_4 _3599_ (.A(_3132_),
    .X(_3133_));
 sky130_fd_sc_hd__clkbuf_4 _3600_ (.A(\egd_top.BitStream_buffer.BS_buffer[70] ),
    .X(_3134_));
 sky130_fd_sc_hd__nand2_1 _3601_ (.A(_3133_),
    .B(_3134_),
    .Y(_3135_));
 sky130_fd_sc_hd__clkbuf_4 _3602_ (.A(\egd_top.BitStream_buffer.BS_buffer[69] ),
    .X(_3136_));
 sky130_fd_sc_hd__inv_2 _3603_ (.A(_3136_),
    .Y(_3137_));
 sky130_fd_sc_hd__and3_1 _3604_ (.A(_3088_),
    .B(\egd_top.BitStream_buffer.pc[2] ),
    .C(_3096_),
    .X(_3138_));
 sky130_fd_sc_hd__clkbuf_4 _3605_ (.A(_3138_),
    .X(_3139_));
 sky130_fd_sc_hd__nand2_1 _3606_ (.A(_3139_),
    .B(_3064_),
    .Y(_3140_));
 sky130_fd_sc_hd__buf_2 _3607_ (.A(_3140_),
    .X(_3141_));
 sky130_fd_sc_hd__or2_1 _3608_ (.A(_3137_),
    .B(_3141_),
    .X(_3142_));
 sky130_fd_sc_hd__o2111a_1 _3609_ (.A1(_3120_),
    .A2(_3124_),
    .B1(_3130_),
    .C1(_3135_),
    .D1(_3142_),
    .X(_3143_));
 sky130_fd_sc_hd__clkbuf_4 _3610_ (.A(\egd_top.BitStream_buffer.BS_buffer[78] ),
    .X(_3144_));
 sky130_fd_sc_hd__nor2_2 _3611_ (.A(_2954_),
    .B(_3058_),
    .Y(_3145_));
 sky130_fd_sc_hd__and2_1 _3612_ (.A(_3145_),
    .B(_3064_),
    .X(_3146_));
 sky130_fd_sc_hd__clkbuf_2 _3613_ (.A(_3146_),
    .X(_3147_));
 sky130_fd_sc_hd__buf_4 _3614_ (.A(_3147_),
    .X(_3148_));
 sky130_fd_sc_hd__clkbuf_4 _3615_ (.A(\egd_top.BitStream_buffer.BS_buffer[79] ),
    .X(_3149_));
 sky130_fd_sc_hd__and2_1 _3616_ (.A(_2964_),
    .B(_3064_),
    .X(_3150_));
 sky130_fd_sc_hd__clkbuf_2 _3617_ (.A(_3150_),
    .X(_3151_));
 sky130_fd_sc_hd__buf_4 _3618_ (.A(_3151_),
    .X(_3152_));
 sky130_fd_sc_hd__nor2_4 _3619_ (.A(_2954_),
    .B(_3087_),
    .Y(_3153_));
 sky130_fd_sc_hd__and2_1 _3620_ (.A(_3153_),
    .B(_3065_),
    .X(_3154_));
 sky130_fd_sc_hd__clkbuf_4 _3621_ (.A(_3154_),
    .X(_3155_));
 sky130_fd_sc_hd__clkbuf_4 _3622_ (.A(\egd_top.BitStream_buffer.BS_buffer[77] ),
    .X(_3156_));
 sky130_fd_sc_hd__nand2_1 _3623_ (.A(_3155_),
    .B(_3156_),
    .Y(_3157_));
 sky130_fd_sc_hd__nor2_4 _3624_ (.A(_2954_),
    .B(_3079_),
    .Y(_3158_));
 sky130_fd_sc_hd__and2_1 _3625_ (.A(_3158_),
    .B(_3065_),
    .X(_3159_));
 sky130_fd_sc_hd__clkbuf_4 _3626_ (.A(_3159_),
    .X(_3160_));
 sky130_fd_sc_hd__clkbuf_4 _3627_ (.A(\egd_top.BitStream_buffer.BS_buffer[76] ),
    .X(_3161_));
 sky130_fd_sc_hd__nand2_1 _3628_ (.A(_3160_),
    .B(_3161_),
    .Y(_3162_));
 sky130_fd_sc_hd__nand2_1 _3629_ (.A(_3157_),
    .B(_3162_),
    .Y(_3163_));
 sky130_fd_sc_hd__a221oi_1 _3630_ (.A1(_3144_),
    .A2(_3148_),
    .B1(_3149_),
    .B2(_3152_),
    .C1(_3163_),
    .Y(_3164_));
 sky130_fd_sc_hd__and4_1 _3631_ (.A(_3094_),
    .B(_3118_),
    .C(_3143_),
    .D(_3164_),
    .X(_3165_));
 sky130_fd_sc_hd__and3_1 _3632_ (.A(\egd_top.BitStream_buffer.pc[6] ),
    .B(\egd_top.BitStream_buffer.pc[4] ),
    .C(\egd_top.BitStream_buffer.pc[5] ),
    .X(_3166_));
 sky130_fd_sc_hd__buf_2 _3633_ (.A(_3166_),
    .X(_3167_));
 sky130_fd_sc_hd__and2_1 _3634_ (.A(_3131_),
    .B(_3167_),
    .X(_3168_));
 sky130_fd_sc_hd__buf_1 _3635_ (.A(_3168_),
    .X(_3169_));
 sky130_fd_sc_hd__clkbuf_4 _3636_ (.A(_3169_),
    .X(_3170_));
 sky130_fd_sc_hd__and2_1 _3637_ (.A(_3122_),
    .B(_3167_),
    .X(_3171_));
 sky130_fd_sc_hd__clkbuf_2 _3638_ (.A(_3171_),
    .X(_3172_));
 sky130_fd_sc_hd__buf_6 _3639_ (.A(_3172_),
    .X(_3173_));
 sky130_fd_sc_hd__inv_2 _3640_ (.A(\egd_top.BitStream_buffer.BS_buffer[116] ),
    .Y(_3174_));
 sky130_fd_sc_hd__nand2_1 _3641_ (.A(_3126_),
    .B(_3167_),
    .Y(_3175_));
 sky130_fd_sc_hd__clkbuf_4 _3642_ (.A(_3175_),
    .X(_3176_));
 sky130_fd_sc_hd__inv_2 _3643_ (.A(_3022_),
    .Y(_3177_));
 sky130_fd_sc_hd__nand2_1 _3644_ (.A(_3139_),
    .B(_3167_),
    .Y(_3178_));
 sky130_fd_sc_hd__clkbuf_4 _3645_ (.A(_3178_),
    .X(_3179_));
 sky130_fd_sc_hd__o22ai_1 _3646_ (.A1(_3174_),
    .A2(_3176_),
    .B1(_3177_),
    .B2(_3179_),
    .Y(_3180_));
 sky130_fd_sc_hd__a221oi_1 _3647_ (.A1(_3025_),
    .A2(_3170_),
    .B1(_3028_),
    .B2(_3173_),
    .C1(_3180_),
    .Y(_3181_));
 sky130_fd_sc_hd__and2_1 _3648_ (.A(_3082_),
    .B(_3166_),
    .X(_3182_));
 sky130_fd_sc_hd__buf_1 _3649_ (.A(_3182_),
    .X(_3183_));
 sky130_fd_sc_hd__buf_4 _3650_ (.A(_3183_),
    .X(_3184_));
 sky130_fd_sc_hd__and2_1 _3651_ (.A(_3090_),
    .B(_3167_),
    .X(_3185_));
 sky130_fd_sc_hd__clkbuf_2 _3652_ (.A(_3185_),
    .X(_3186_));
 sky130_fd_sc_hd__buf_6 _3653_ (.A(_3186_),
    .X(_3187_));
 sky130_fd_sc_hd__inv_2 _3654_ (.A(_3040_),
    .Y(_3188_));
 sky130_fd_sc_hd__nand2_1 _3655_ (.A(_3072_),
    .B(_3167_),
    .Y(_3189_));
 sky130_fd_sc_hd__clkbuf_4 _3656_ (.A(_3189_),
    .X(_3190_));
 sky130_fd_sc_hd__and2_1 _3657_ (.A(_3061_),
    .B(_3167_),
    .X(_3191_));
 sky130_fd_sc_hd__clkbuf_4 _3658_ (.A(_3191_),
    .X(_3192_));
 sky130_fd_sc_hd__nand2_1 _3659_ (.A(_3192_),
    .B(_3037_),
    .Y(_3193_));
 sky130_fd_sc_hd__o21ai_1 _3660_ (.A1(_3188_),
    .A2(_3190_),
    .B1(_3193_),
    .Y(_3194_));
 sky130_fd_sc_hd__a221oi_1 _3661_ (.A1(_3031_),
    .A2(_3184_),
    .B1(_3034_),
    .B2(_3187_),
    .C1(_3194_),
    .Y(_3195_));
 sky130_fd_sc_hd__and2_1 _3662_ (.A(_3098_),
    .B(_3166_),
    .X(_3196_));
 sky130_fd_sc_hd__buf_1 _3663_ (.A(_3196_),
    .X(_3197_));
 sky130_fd_sc_hd__buf_4 _3664_ (.A(_3197_),
    .X(_3198_));
 sky130_fd_sc_hd__and2_1 _3665_ (.A(_3103_),
    .B(_3167_),
    .X(_3199_));
 sky130_fd_sc_hd__buf_1 _3666_ (.A(_3199_),
    .X(_3200_));
 sky130_fd_sc_hd__buf_4 _3667_ (.A(_3200_),
    .X(_3201_));
 sky130_fd_sc_hd__inv_2 _3668_ (.A(\egd_top.BitStream_buffer.BS_buffer[112] ),
    .Y(_3202_));
 sky130_fd_sc_hd__nand2_1 _3669_ (.A(_3109_),
    .B(_3167_),
    .Y(_3203_));
 sky130_fd_sc_hd__clkbuf_4 _3670_ (.A(_3203_),
    .X(_3204_));
 sky130_fd_sc_hd__and2_1 _3671_ (.A(_3112_),
    .B(_3167_),
    .X(_3205_));
 sky130_fd_sc_hd__clkbuf_4 _3672_ (.A(_3205_),
    .X(_3206_));
 sky130_fd_sc_hd__nand2_1 _3673_ (.A(_3206_),
    .B(_3010_),
    .Y(_3207_));
 sky130_fd_sc_hd__o21ai_1 _3674_ (.A1(_3202_),
    .A2(_3204_),
    .B1(_3207_),
    .Y(_3208_));
 sky130_fd_sc_hd__a221oi_1 _3675_ (.A1(_3013_),
    .A2(_3198_),
    .B1(_3016_),
    .B2(_3201_),
    .C1(_3208_),
    .Y(_3209_));
 sky130_fd_sc_hd__and2_1 _3676_ (.A(_3145_),
    .B(_3166_),
    .X(_3210_));
 sky130_fd_sc_hd__buf_1 _3677_ (.A(_3210_),
    .X(_3211_));
 sky130_fd_sc_hd__clkbuf_4 _3678_ (.A(_3211_),
    .X(_3212_));
 sky130_fd_sc_hd__and2_1 _3679_ (.A(_2964_),
    .B(_3166_),
    .X(_3213_));
 sky130_fd_sc_hd__buf_1 _3680_ (.A(_3213_),
    .X(_3214_));
 sky130_fd_sc_hd__clkbuf_4 _3681_ (.A(_3214_),
    .X(_3215_));
 sky130_fd_sc_hd__inv_2 _3682_ (.A(_3044_),
    .Y(_3216_));
 sky130_fd_sc_hd__nand2_1 _3683_ (.A(_3158_),
    .B(_3167_),
    .Y(_3217_));
 sky130_fd_sc_hd__clkbuf_4 _3684_ (.A(_3217_),
    .X(_3218_));
 sky130_fd_sc_hd__inv_2 _3685_ (.A(_3047_),
    .Y(_3219_));
 sky130_fd_sc_hd__nand2_1 _3686_ (.A(_3153_),
    .B(_3167_),
    .Y(_3220_));
 sky130_fd_sc_hd__clkbuf_4 _3687_ (.A(_3220_),
    .X(_3221_));
 sky130_fd_sc_hd__o22ai_1 _3688_ (.A1(_3216_),
    .A2(_3218_),
    .B1(_3219_),
    .B2(_3221_),
    .Y(_3222_));
 sky130_fd_sc_hd__a221oi_1 _3689_ (.A1(_3050_),
    .A2(_3212_),
    .B1(_3053_),
    .B2(_3215_),
    .C1(_3222_),
    .Y(_3223_));
 sky130_fd_sc_hd__and4_1 _3690_ (.A(_3181_),
    .B(_3195_),
    .C(_3209_),
    .D(_3223_),
    .X(_3224_));
 sky130_fd_sc_hd__buf_4 _3691_ (.A(\egd_top.BitStream_buffer.BS_buffer[90] ),
    .X(_3225_));
 sky130_fd_sc_hd__or3_1 _3692_ (.A(\egd_top.BitStream_buffer.pc[5] ),
    .B(_2965_),
    .C(_3062_),
    .X(_3226_));
 sky130_fd_sc_hd__inv_2 _3693_ (.A(_3226_),
    .Y(_3227_));
 sky130_fd_sc_hd__buf_2 _3694_ (.A(_3227_),
    .X(_3228_));
 sky130_fd_sc_hd__and2_1 _3695_ (.A(_3061_),
    .B(_3228_),
    .X(_3229_));
 sky130_fd_sc_hd__buf_1 _3696_ (.A(_3229_),
    .X(_3230_));
 sky130_fd_sc_hd__clkbuf_4 _3697_ (.A(_3230_),
    .X(_3231_));
 sky130_fd_sc_hd__clkbuf_4 _3698_ (.A(\egd_top.BitStream_buffer.BS_buffer[91] ),
    .X(_3232_));
 sky130_fd_sc_hd__and2_1 _3699_ (.A(_3072_),
    .B(_3228_),
    .X(_3233_));
 sky130_fd_sc_hd__clkbuf_2 _3700_ (.A(_3233_),
    .X(_3234_));
 sky130_fd_sc_hd__buf_4 _3701_ (.A(_3234_),
    .X(_3235_));
 sky130_fd_sc_hd__inv_2 _3702_ (.A(\egd_top.BitStream_buffer.BS_buffer[88] ),
    .Y(_3236_));
 sky130_fd_sc_hd__nand2_1 _3703_ (.A(_3082_),
    .B(_3228_),
    .Y(_3237_));
 sky130_fd_sc_hd__clkbuf_4 _3704_ (.A(_3237_),
    .X(_3238_));
 sky130_fd_sc_hd__inv_2 _3705_ (.A(\egd_top.BitStream_buffer.BS_buffer[89] ),
    .Y(_3239_));
 sky130_fd_sc_hd__nand2_1 _3706_ (.A(_3090_),
    .B(_3228_),
    .Y(_3240_));
 sky130_fd_sc_hd__clkbuf_4 _3707_ (.A(_3240_),
    .X(_3241_));
 sky130_fd_sc_hd__o22ai_1 _3708_ (.A1(_3236_),
    .A2(_3238_),
    .B1(_3239_),
    .B2(_3241_),
    .Y(_3242_));
 sky130_fd_sc_hd__a221oi_1 _3709_ (.A1(_3225_),
    .A2(_3231_),
    .B1(_3232_),
    .B2(_3235_),
    .C1(_3242_),
    .Y(_3243_));
 sky130_fd_sc_hd__inv_2 _3710_ (.A(_3112_),
    .Y(_3244_));
 sky130_fd_sc_hd__nor2_1 _3711_ (.A(_3226_),
    .B(_3244_),
    .Y(_3245_));
 sky130_fd_sc_hd__clkbuf_4 _3712_ (.A(_3245_),
    .X(_3246_));
 sky130_fd_sc_hd__clkbuf_4 _3713_ (.A(\egd_top.BitStream_buffer.BS_buffer[81] ),
    .X(_3247_));
 sky130_fd_sc_hd__nand2_1 _3714_ (.A(_3246_),
    .B(_3247_),
    .Y(_3248_));
 sky130_fd_sc_hd__and2_1 _3715_ (.A(_3103_),
    .B(_3228_),
    .X(_3249_));
 sky130_fd_sc_hd__clkbuf_4 _3716_ (.A(_3249_),
    .X(_3250_));
 sky130_fd_sc_hd__buf_4 _3717_ (.A(\egd_top.BitStream_buffer.BS_buffer[83] ),
    .X(_3251_));
 sky130_fd_sc_hd__nand2_1 _3718_ (.A(_3250_),
    .B(_3251_),
    .Y(_3252_));
 sky130_fd_sc_hd__and2_1 _3719_ (.A(_3109_),
    .B(_3228_),
    .X(_3253_));
 sky130_fd_sc_hd__clkbuf_4 _3720_ (.A(_3253_),
    .X(_3254_));
 sky130_fd_sc_hd__clkbuf_4 _3721_ (.A(\egd_top.BitStream_buffer.BS_buffer[80] ),
    .X(_3255_));
 sky130_fd_sc_hd__nand2_1 _3722_ (.A(_3254_),
    .B(_3255_),
    .Y(_3256_));
 sky130_fd_sc_hd__and2_1 _3723_ (.A(_3098_),
    .B(_3227_),
    .X(_3257_));
 sky130_fd_sc_hd__clkbuf_4 _3724_ (.A(_3257_),
    .X(_3258_));
 sky130_fd_sc_hd__clkbuf_4 _3725_ (.A(\egd_top.BitStream_buffer.BS_buffer[82] ),
    .X(_3259_));
 sky130_fd_sc_hd__nand2_1 _3726_ (.A(_3258_),
    .B(_3259_),
    .Y(_3260_));
 sky130_fd_sc_hd__and4_1 _3727_ (.A(_3248_),
    .B(_3252_),
    .C(_3256_),
    .D(_3260_),
    .X(_3261_));
 sky130_fd_sc_hd__inv_2 _3728_ (.A(\egd_top.BitStream_buffer.BS_buffer[84] ),
    .Y(_3262_));
 sky130_fd_sc_hd__nand2_2 _3729_ (.A(_3126_),
    .B(_3228_),
    .Y(_3263_));
 sky130_fd_sc_hd__clkbuf_4 _3730_ (.A(_3263_),
    .X(_3264_));
 sky130_fd_sc_hd__buf_4 _3731_ (.A(\egd_top.BitStream_buffer.BS_buffer[85] ),
    .X(_3265_));
 sky130_fd_sc_hd__inv_2 _3732_ (.A(_3265_),
    .Y(_3266_));
 sky130_fd_sc_hd__nand2_1 _3733_ (.A(_3139_),
    .B(_3228_),
    .Y(_3267_));
 sky130_fd_sc_hd__clkbuf_4 _3734_ (.A(_3267_),
    .X(_3268_));
 sky130_fd_sc_hd__o22ai_1 _3735_ (.A1(_3262_),
    .A2(_3264_),
    .B1(_3266_),
    .B2(_3268_),
    .Y(_3269_));
 sky130_fd_sc_hd__and2_1 _3736_ (.A(_3131_),
    .B(_3228_),
    .X(_3270_));
 sky130_fd_sc_hd__clkbuf_4 _3737_ (.A(_3270_),
    .X(_3271_));
 sky130_fd_sc_hd__clkbuf_4 _3738_ (.A(\egd_top.BitStream_buffer.BS_buffer[86] ),
    .X(_3272_));
 sky130_fd_sc_hd__and2_1 _3739_ (.A(_3122_),
    .B(_3228_),
    .X(_3273_));
 sky130_fd_sc_hd__clkbuf_4 _3740_ (.A(_3273_),
    .X(_3274_));
 sky130_fd_sc_hd__clkbuf_4 _3741_ (.A(\egd_top.BitStream_buffer.BS_buffer[87] ),
    .X(_3275_));
 sky130_fd_sc_hd__a22o_1 _3742_ (.A1(_3271_),
    .A2(_3272_),
    .B1(_3274_),
    .B2(_3275_),
    .X(_3276_));
 sky130_fd_sc_hd__nor2_1 _3743_ (.A(_3269_),
    .B(_3276_),
    .Y(_3277_));
 sky130_fd_sc_hd__clkbuf_4 _3744_ (.A(\egd_top.BitStream_buffer.BS_buffer[94] ),
    .X(_3278_));
 sky130_fd_sc_hd__and2_1 _3745_ (.A(_3145_),
    .B(_3227_),
    .X(_3279_));
 sky130_fd_sc_hd__buf_1 _3746_ (.A(_3279_),
    .X(_3280_));
 sky130_fd_sc_hd__clkbuf_4 _3747_ (.A(_3280_),
    .X(_3281_));
 sky130_fd_sc_hd__clkbuf_4 _3748_ (.A(\egd_top.BitStream_buffer.BS_buffer[95] ),
    .X(_3282_));
 sky130_fd_sc_hd__and2_1 _3749_ (.A(_2964_),
    .B(_3227_),
    .X(_3283_));
 sky130_fd_sc_hd__buf_1 _3750_ (.A(_3283_),
    .X(_3284_));
 sky130_fd_sc_hd__clkbuf_4 _3751_ (.A(_3284_),
    .X(_3285_));
 sky130_fd_sc_hd__buf_4 _3752_ (.A(\egd_top.BitStream_buffer.BS_buffer[92] ),
    .X(_3286_));
 sky130_fd_sc_hd__inv_2 _3753_ (.A(_3286_),
    .Y(_3287_));
 sky130_fd_sc_hd__nand2_1 _3754_ (.A(_3158_),
    .B(_3228_),
    .Y(_3288_));
 sky130_fd_sc_hd__clkbuf_4 _3755_ (.A(_3288_),
    .X(_3289_));
 sky130_fd_sc_hd__clkbuf_4 _3756_ (.A(\egd_top.BitStream_buffer.BS_buffer[93] ),
    .X(_3290_));
 sky130_fd_sc_hd__inv_2 _3757_ (.A(_3290_),
    .Y(_3291_));
 sky130_fd_sc_hd__nand2_1 _3758_ (.A(_3153_),
    .B(_3228_),
    .Y(_3292_));
 sky130_fd_sc_hd__clkbuf_4 _3759_ (.A(_3292_),
    .X(_3293_));
 sky130_fd_sc_hd__o22ai_1 _3760_ (.A1(_3287_),
    .A2(_3289_),
    .B1(_3291_),
    .B2(_3293_),
    .Y(_3294_));
 sky130_fd_sc_hd__a221oi_1 _3761_ (.A1(_3278_),
    .A2(_3281_),
    .B1(_3282_),
    .B2(_3285_),
    .C1(_3294_),
    .Y(_3295_));
 sky130_fd_sc_hd__and4_1 _3762_ (.A(_3243_),
    .B(_3261_),
    .C(_3277_),
    .D(_3295_),
    .X(_3296_));
 sky130_fd_sc_hd__clkbuf_4 _3763_ (.A(\egd_top.BitStream_buffer.BS_buffer[106] ),
    .X(_3297_));
 sky130_fd_sc_hd__or3_1 _3764_ (.A(\egd_top.BitStream_buffer.pc[4] ),
    .B(_2965_),
    .C(_3063_),
    .X(_3298_));
 sky130_fd_sc_hd__inv_2 _3765_ (.A(_3298_),
    .Y(_3299_));
 sky130_fd_sc_hd__buf_2 _3766_ (.A(_3299_),
    .X(_3300_));
 sky130_fd_sc_hd__and2_1 _3767_ (.A(_3061_),
    .B(_3300_),
    .X(_3301_));
 sky130_fd_sc_hd__buf_1 _3768_ (.A(_3301_),
    .X(_3302_));
 sky130_fd_sc_hd__clkbuf_4 _3769_ (.A(_3302_),
    .X(_3303_));
 sky130_fd_sc_hd__clkbuf_4 _3770_ (.A(\egd_top.BitStream_buffer.BS_buffer[107] ),
    .X(_3304_));
 sky130_fd_sc_hd__and2_1 _3771_ (.A(_3072_),
    .B(_3300_),
    .X(_3305_));
 sky130_fd_sc_hd__buf_1 _3772_ (.A(_3305_),
    .X(_3306_));
 sky130_fd_sc_hd__buf_4 _3773_ (.A(_3306_),
    .X(_3307_));
 sky130_fd_sc_hd__and2_1 _3774_ (.A(_3090_),
    .B(_3300_),
    .X(_3308_));
 sky130_fd_sc_hd__buf_4 _3775_ (.A(_3308_),
    .X(_3309_));
 sky130_fd_sc_hd__clkbuf_4 _3776_ (.A(\egd_top.BitStream_buffer.BS_buffer[105] ),
    .X(_3310_));
 sky130_fd_sc_hd__nand2_1 _3777_ (.A(_3309_),
    .B(_3310_),
    .Y(_3311_));
 sky130_fd_sc_hd__and2_1 _3778_ (.A(_3082_),
    .B(_3300_),
    .X(_3312_));
 sky130_fd_sc_hd__clkbuf_4 _3779_ (.A(_3312_),
    .X(_3313_));
 sky130_fd_sc_hd__clkbuf_4 _3780_ (.A(\egd_top.BitStream_buffer.BS_buffer[104] ),
    .X(_3314_));
 sky130_fd_sc_hd__nand2_1 _3781_ (.A(_3313_),
    .B(_3314_),
    .Y(_3315_));
 sky130_fd_sc_hd__nand2_1 _3782_ (.A(_3311_),
    .B(_3315_),
    .Y(_3316_));
 sky130_fd_sc_hd__a221oi_1 _3783_ (.A1(_3297_),
    .A2(_3303_),
    .B1(_3304_),
    .B2(_3307_),
    .C1(_3316_),
    .Y(_3317_));
 sky130_fd_sc_hd__clkbuf_4 _3784_ (.A(\egd_top.BitStream_buffer.BS_buffer[96] ),
    .X(_3318_));
 sky130_fd_sc_hd__and2_1 _3785_ (.A(_3109_),
    .B(_3300_),
    .X(_3319_));
 sky130_fd_sc_hd__buf_1 _3786_ (.A(_3319_),
    .X(_3320_));
 sky130_fd_sc_hd__clkbuf_4 _3787_ (.A(_3320_),
    .X(_3321_));
 sky130_fd_sc_hd__buf_4 _3788_ (.A(\egd_top.BitStream_buffer.BS_buffer[97] ),
    .X(_3322_));
 sky130_fd_sc_hd__nor2_1 _3789_ (.A(_3298_),
    .B(_3244_),
    .Y(_3323_));
 sky130_fd_sc_hd__clkbuf_4 _3790_ (.A(_3323_),
    .X(_3324_));
 sky130_fd_sc_hd__and2_1 _3791_ (.A(_3103_),
    .B(_3300_),
    .X(_3325_));
 sky130_fd_sc_hd__clkbuf_4 _3792_ (.A(_3325_),
    .X(_3326_));
 sky130_fd_sc_hd__clkbuf_4 _3793_ (.A(\egd_top.BitStream_buffer.BS_buffer[99] ),
    .X(_3327_));
 sky130_fd_sc_hd__nand2_1 _3794_ (.A(_3326_),
    .B(_3327_),
    .Y(_3328_));
 sky130_fd_sc_hd__and2_1 _3795_ (.A(_3098_),
    .B(_3300_),
    .X(_3329_));
 sky130_fd_sc_hd__clkbuf_4 _3796_ (.A(_3329_),
    .X(_3330_));
 sky130_fd_sc_hd__clkbuf_4 _3797_ (.A(\egd_top.BitStream_buffer.BS_buffer[98] ),
    .X(_3331_));
 sky130_fd_sc_hd__nand2_1 _3798_ (.A(_3330_),
    .B(_3331_),
    .Y(_3332_));
 sky130_fd_sc_hd__nand2_1 _3799_ (.A(_3328_),
    .B(_3332_),
    .Y(_3333_));
 sky130_fd_sc_hd__a221oi_1 _3800_ (.A1(_3318_),
    .A2(_3321_),
    .B1(_3322_),
    .B2(_3324_),
    .C1(_3333_),
    .Y(_3334_));
 sky130_fd_sc_hd__buf_4 _3801_ (.A(\egd_top.BitStream_buffer.BS_buffer[103] ),
    .X(_3335_));
 sky130_fd_sc_hd__inv_2 _3802_ (.A(_3335_),
    .Y(_3336_));
 sky130_fd_sc_hd__nand2_1 _3803_ (.A(_3122_),
    .B(_3300_),
    .Y(_3337_));
 sky130_fd_sc_hd__clkbuf_4 _3804_ (.A(_3337_),
    .X(_3338_));
 sky130_fd_sc_hd__and2_1 _3805_ (.A(_3126_),
    .B(_3300_),
    .X(_3339_));
 sky130_fd_sc_hd__clkbuf_4 _3806_ (.A(_3339_),
    .X(_3340_));
 sky130_fd_sc_hd__clkbuf_4 _3807_ (.A(\egd_top.BitStream_buffer.BS_buffer[100] ),
    .X(_3341_));
 sky130_fd_sc_hd__nand2_1 _3808_ (.A(_3340_),
    .B(_3341_),
    .Y(_3342_));
 sky130_fd_sc_hd__and2_1 _3809_ (.A(_3131_),
    .B(_3300_),
    .X(_3343_));
 sky130_fd_sc_hd__clkbuf_4 _3810_ (.A(_3343_),
    .X(_3344_));
 sky130_fd_sc_hd__clkbuf_4 _3811_ (.A(\egd_top.BitStream_buffer.BS_buffer[102] ),
    .X(_3345_));
 sky130_fd_sc_hd__nand2_1 _3812_ (.A(_3344_),
    .B(_3345_),
    .Y(_3346_));
 sky130_fd_sc_hd__clkbuf_4 _3813_ (.A(\egd_top.BitStream_buffer.BS_buffer[101] ),
    .X(_3347_));
 sky130_fd_sc_hd__inv_2 _3814_ (.A(_3347_),
    .Y(_3348_));
 sky130_fd_sc_hd__nand2_1 _3815_ (.A(_3139_),
    .B(_3299_),
    .Y(_3349_));
 sky130_fd_sc_hd__buf_2 _3816_ (.A(_3349_),
    .X(_3350_));
 sky130_fd_sc_hd__or2_1 _3817_ (.A(_3348_),
    .B(_3350_),
    .X(_3351_));
 sky130_fd_sc_hd__o2111a_1 _3818_ (.A1(_3336_),
    .A2(_3338_),
    .B1(_3342_),
    .C1(_3346_),
    .D1(_3351_),
    .X(_3352_));
 sky130_fd_sc_hd__clkbuf_4 _3819_ (.A(\egd_top.BitStream_buffer.BS_buffer[108] ),
    .X(_3353_));
 sky130_fd_sc_hd__and2_1 _3820_ (.A(_3158_),
    .B(_3299_),
    .X(_3354_));
 sky130_fd_sc_hd__buf_1 _3821_ (.A(_3354_),
    .X(_3355_));
 sky130_fd_sc_hd__clkbuf_4 _3822_ (.A(_3355_),
    .X(_3356_));
 sky130_fd_sc_hd__clkbuf_4 _3823_ (.A(\egd_top.BitStream_buffer.BS_buffer[109] ),
    .X(_3357_));
 sky130_fd_sc_hd__and2_1 _3824_ (.A(_3153_),
    .B(_3299_),
    .X(_3358_));
 sky130_fd_sc_hd__buf_1 _3825_ (.A(_3358_),
    .X(_3359_));
 sky130_fd_sc_hd__buf_4 _3826_ (.A(_3359_),
    .X(_3360_));
 sky130_fd_sc_hd__inv_2 _3827_ (.A(\egd_top.BitStream_buffer.BS_buffer[111] ),
    .Y(_3361_));
 sky130_fd_sc_hd__nand2_1 _3828_ (.A(_2964_),
    .B(_3300_),
    .Y(_3362_));
 sky130_fd_sc_hd__clkbuf_4 _3829_ (.A(_3362_),
    .X(_3363_));
 sky130_fd_sc_hd__and2_1 _3830_ (.A(_3145_),
    .B(_3300_),
    .X(_3364_));
 sky130_fd_sc_hd__clkbuf_4 _3831_ (.A(_3364_),
    .X(_3365_));
 sky130_fd_sc_hd__nand2_1 _3832_ (.A(_3365_),
    .B(\egd_top.BitStream_buffer.BS_buffer[110] ),
    .Y(_3366_));
 sky130_fd_sc_hd__o21ai_1 _3833_ (.A1(_3361_),
    .A2(_3363_),
    .B1(_3366_),
    .Y(_3367_));
 sky130_fd_sc_hd__a221oi_1 _3834_ (.A1(_3353_),
    .A2(_3356_),
    .B1(_3357_),
    .B2(_3360_),
    .C1(_3367_),
    .Y(_3368_));
 sky130_fd_sc_hd__and4_1 _3835_ (.A(_3317_),
    .B(_3334_),
    .C(_3352_),
    .D(_3368_),
    .X(_3369_));
 sky130_fd_sc_hd__and4_1 _3836_ (.A(_3165_),
    .B(_3224_),
    .C(_3296_),
    .D(_3369_),
    .X(_0322_));
 sky130_fd_sc_hd__buf_4 _3837_ (.A(\egd_top.BitStream_buffer.BS_buffer[42] ),
    .X(_0323_));
 sky130_fd_sc_hd__and3_2 _3838_ (.A(_2965_),
    .B(_3062_),
    .C(\egd_top.BitStream_buffer.pc[5] ),
    .X(_0324_));
 sky130_fd_sc_hd__buf_2 _3839_ (.A(_0324_),
    .X(_0325_));
 sky130_fd_sc_hd__and2_1 _3840_ (.A(_3061_),
    .B(_0325_),
    .X(_0326_));
 sky130_fd_sc_hd__buf_1 _3841_ (.A(_0326_),
    .X(_0327_));
 sky130_fd_sc_hd__clkbuf_4 _3842_ (.A(_0327_),
    .X(_0328_));
 sky130_fd_sc_hd__clkbuf_4 _3843_ (.A(\egd_top.BitStream_buffer.BS_buffer[43] ),
    .X(_0329_));
 sky130_fd_sc_hd__and2_1 _3844_ (.A(_3072_),
    .B(_0325_),
    .X(_0330_));
 sky130_fd_sc_hd__clkbuf_2 _3845_ (.A(_0330_),
    .X(_0331_));
 sky130_fd_sc_hd__buf_6 _3846_ (.A(_0331_),
    .X(_0332_));
 sky130_fd_sc_hd__and2_1 _3847_ (.A(_3090_),
    .B(_0325_),
    .X(_0333_));
 sky130_fd_sc_hd__buf_4 _3848_ (.A(_0333_),
    .X(_0334_));
 sky130_fd_sc_hd__buf_4 _3849_ (.A(\egd_top.BitStream_buffer.BS_buffer[41] ),
    .X(_0335_));
 sky130_fd_sc_hd__nand2_1 _3850_ (.A(_0334_),
    .B(_0335_),
    .Y(_0336_));
 sky130_fd_sc_hd__and2_1 _3851_ (.A(_3082_),
    .B(_0325_),
    .X(_0337_));
 sky130_fd_sc_hd__buf_4 _3852_ (.A(_0337_),
    .X(_0338_));
 sky130_fd_sc_hd__clkbuf_4 _3853_ (.A(\egd_top.BitStream_buffer.BS_buffer[40] ),
    .X(_0339_));
 sky130_fd_sc_hd__nand2_1 _3854_ (.A(_0338_),
    .B(_0339_),
    .Y(_0340_));
 sky130_fd_sc_hd__nand2_1 _3855_ (.A(_0336_),
    .B(_0340_),
    .Y(_0341_));
 sky130_fd_sc_hd__a221oi_1 _3856_ (.A1(_0323_),
    .A2(_0328_),
    .B1(_0329_),
    .B2(_0332_),
    .C1(_0341_),
    .Y(_0342_));
 sky130_fd_sc_hd__inv_2 _3857_ (.A(\egd_top.BitStream_buffer.BS_buffer[36] ),
    .Y(_0343_));
 sky130_fd_sc_hd__nand2_1 _3858_ (.A(_3126_),
    .B(_0325_),
    .Y(_0344_));
 sky130_fd_sc_hd__clkbuf_4 _3859_ (.A(_0344_),
    .X(_0345_));
 sky130_fd_sc_hd__clkbuf_4 _3860_ (.A(\egd_top.BitStream_buffer.BS_buffer[37] ),
    .X(_0346_));
 sky130_fd_sc_hd__inv_2 _3861_ (.A(_0346_),
    .Y(_0347_));
 sky130_fd_sc_hd__nand2_1 _3862_ (.A(_3139_),
    .B(_0325_),
    .Y(_0348_));
 sky130_fd_sc_hd__clkbuf_4 _3863_ (.A(_0348_),
    .X(_0349_));
 sky130_fd_sc_hd__o22ai_1 _3864_ (.A1(_0343_),
    .A2(_0345_),
    .B1(_0347_),
    .B2(_0349_),
    .Y(_0350_));
 sky130_fd_sc_hd__and2_1 _3865_ (.A(_3131_),
    .B(_0325_),
    .X(_0351_));
 sky130_fd_sc_hd__clkbuf_4 _3866_ (.A(_0351_),
    .X(_0352_));
 sky130_fd_sc_hd__clkbuf_4 _3867_ (.A(\egd_top.BitStream_buffer.BS_buffer[38] ),
    .X(_0353_));
 sky130_fd_sc_hd__and2_1 _3868_ (.A(_3122_),
    .B(_0325_),
    .X(_0354_));
 sky130_fd_sc_hd__clkbuf_4 _3869_ (.A(_0354_),
    .X(_0355_));
 sky130_fd_sc_hd__clkbuf_4 _3870_ (.A(\egd_top.BitStream_buffer.BS_buffer[39] ),
    .X(_0356_));
 sky130_fd_sc_hd__a22o_1 _3871_ (.A1(_0352_),
    .A2(_0353_),
    .B1(_0355_),
    .B2(_0356_),
    .X(_0357_));
 sky130_fd_sc_hd__nor2_1 _3872_ (.A(_0350_),
    .B(_0357_),
    .Y(_0358_));
 sky130_fd_sc_hd__buf_4 _3873_ (.A(\egd_top.BitStream_buffer.BS_buffer[32] ),
    .X(_0359_));
 sky130_fd_sc_hd__and2_1 _3874_ (.A(_3109_),
    .B(_0324_),
    .X(_0360_));
 sky130_fd_sc_hd__buf_1 _3875_ (.A(_0360_),
    .X(_0361_));
 sky130_fd_sc_hd__clkbuf_4 _3876_ (.A(_0361_),
    .X(_0362_));
 sky130_fd_sc_hd__buf_4 _3877_ (.A(\egd_top.BitStream_buffer.BS_buffer[33] ),
    .X(_0363_));
 sky130_fd_sc_hd__and2_1 _3878_ (.A(_3112_),
    .B(_0324_),
    .X(_0364_));
 sky130_fd_sc_hd__buf_1 _3879_ (.A(_0364_),
    .X(_0365_));
 sky130_fd_sc_hd__clkbuf_4 _3880_ (.A(_0365_),
    .X(_0366_));
 sky130_fd_sc_hd__inv_2 _3881_ (.A(\egd_top.BitStream_buffer.BS_buffer[34] ),
    .Y(_0367_));
 sky130_fd_sc_hd__nand2_1 _3882_ (.A(_3098_),
    .B(_0325_),
    .Y(_0368_));
 sky130_fd_sc_hd__clkbuf_4 _3883_ (.A(_0368_),
    .X(_0369_));
 sky130_fd_sc_hd__and2_1 _3884_ (.A(_3103_),
    .B(_0325_),
    .X(_0370_));
 sky130_fd_sc_hd__clkbuf_4 _3885_ (.A(_0370_),
    .X(_0371_));
 sky130_fd_sc_hd__clkbuf_4 _3886_ (.A(\egd_top.BitStream_buffer.BS_buffer[35] ),
    .X(_0372_));
 sky130_fd_sc_hd__nand2_1 _3887_ (.A(_0371_),
    .B(_0372_),
    .Y(_0373_));
 sky130_fd_sc_hd__o21ai_1 _3888_ (.A1(_0367_),
    .A2(_0369_),
    .B1(_0373_),
    .Y(_0374_));
 sky130_fd_sc_hd__a221oi_1 _3889_ (.A1(_0359_),
    .A2(_0362_),
    .B1(_0363_),
    .B2(_0366_),
    .C1(_0374_),
    .Y(_0375_));
 sky130_fd_sc_hd__clkbuf_4 _3890_ (.A(\egd_top.BitStream_buffer.BS_buffer[44] ),
    .X(_0376_));
 sky130_fd_sc_hd__and2_1 _3891_ (.A(_3158_),
    .B(_0324_),
    .X(_0377_));
 sky130_fd_sc_hd__buf_1 _3892_ (.A(_0377_),
    .X(_0378_));
 sky130_fd_sc_hd__clkbuf_4 _3893_ (.A(_0378_),
    .X(_0379_));
 sky130_fd_sc_hd__clkbuf_4 _3894_ (.A(\egd_top.BitStream_buffer.BS_buffer[45] ),
    .X(_0380_));
 sky130_fd_sc_hd__and2_1 _3895_ (.A(_3153_),
    .B(_0324_),
    .X(_0381_));
 sky130_fd_sc_hd__buf_1 _3896_ (.A(_0381_),
    .X(_0382_));
 sky130_fd_sc_hd__clkbuf_4 _3897_ (.A(_0382_),
    .X(_0383_));
 sky130_fd_sc_hd__inv_2 _3898_ (.A(\egd_top.BitStream_buffer.BS_buffer[47] ),
    .Y(_0384_));
 sky130_fd_sc_hd__nand2_1 _3899_ (.A(_2964_),
    .B(_0325_),
    .Y(_0385_));
 sky130_fd_sc_hd__clkbuf_4 _3900_ (.A(_0385_),
    .X(_0386_));
 sky130_fd_sc_hd__and2_1 _3901_ (.A(_3145_),
    .B(_0325_),
    .X(_0387_));
 sky130_fd_sc_hd__clkbuf_4 _3902_ (.A(_0387_),
    .X(_0388_));
 sky130_fd_sc_hd__clkbuf_4 _3903_ (.A(\egd_top.BitStream_buffer.BS_buffer[46] ),
    .X(_0389_));
 sky130_fd_sc_hd__nand2_1 _3904_ (.A(_0388_),
    .B(_0389_),
    .Y(_0390_));
 sky130_fd_sc_hd__o21ai_1 _3905_ (.A1(_0384_),
    .A2(_0386_),
    .B1(_0390_),
    .Y(_0391_));
 sky130_fd_sc_hd__a221oi_1 _3906_ (.A1(_0376_),
    .A2(_0379_),
    .B1(_0380_),
    .B2(_0383_),
    .C1(_0391_),
    .Y(_0392_));
 sky130_fd_sc_hd__and4_1 _3907_ (.A(_0342_),
    .B(_0358_),
    .C(_0375_),
    .D(_0392_),
    .X(_0393_));
 sky130_fd_sc_hd__inv_2 _3908_ (.A(\egd_top.BitStream_buffer.BS_buffer[53] ),
    .Y(_0394_));
 sky130_fd_sc_hd__buf_2 _3909_ (.A(_2966_),
    .X(_0395_));
 sky130_fd_sc_hd__nand2_1 _3910_ (.A(_3139_),
    .B(_0395_),
    .Y(_0396_));
 sky130_fd_sc_hd__clkbuf_4 _3911_ (.A(_0396_),
    .X(_0397_));
 sky130_fd_sc_hd__and2_1 _3912_ (.A(_3131_),
    .B(_0395_),
    .X(_0398_));
 sky130_fd_sc_hd__clkbuf_4 _3913_ (.A(_0398_),
    .X(_0399_));
 sky130_fd_sc_hd__clkbuf_4 _3914_ (.A(\egd_top.BitStream_buffer.BS_buffer[54] ),
    .X(_0400_));
 sky130_fd_sc_hd__nand2_1 _3915_ (.A(_0399_),
    .B(_0400_),
    .Y(_0401_));
 sky130_fd_sc_hd__and2_1 _3916_ (.A(_3126_),
    .B(_0395_),
    .X(_0402_));
 sky130_fd_sc_hd__clkbuf_4 _3917_ (.A(_0402_),
    .X(_0403_));
 sky130_fd_sc_hd__clkbuf_4 _3918_ (.A(\egd_top.BitStream_buffer.BS_buffer[52] ),
    .X(_0404_));
 sky130_fd_sc_hd__nand2_1 _3919_ (.A(_0403_),
    .B(_0404_),
    .Y(_0405_));
 sky130_fd_sc_hd__inv_2 _3920_ (.A(\egd_top.BitStream_buffer.BS_buffer[55] ),
    .Y(_0406_));
 sky130_fd_sc_hd__nand2_1 _3921_ (.A(_3122_),
    .B(_0395_),
    .Y(_0407_));
 sky130_fd_sc_hd__clkbuf_4 _3922_ (.A(_0407_),
    .X(_0408_));
 sky130_fd_sc_hd__or2_1 _3923_ (.A(_0406_),
    .B(_0408_),
    .X(_0409_));
 sky130_fd_sc_hd__o2111a_1 _3924_ (.A1(_0394_),
    .A2(_0397_),
    .B1(_0401_),
    .C1(_0405_),
    .D1(_0409_),
    .X(_0410_));
 sky130_fd_sc_hd__clkbuf_4 _3925_ (.A(\egd_top.BitStream_buffer.BS_buffer[59] ),
    .X(_0411_));
 sky130_fd_sc_hd__inv_2 _3926_ (.A(_0411_),
    .Y(_0412_));
 sky130_fd_sc_hd__nand2_1 _3927_ (.A(_3072_),
    .B(_0395_),
    .Y(_0413_));
 sky130_fd_sc_hd__clkbuf_4 _3928_ (.A(_0413_),
    .X(_0414_));
 sky130_fd_sc_hd__and2_1 _3929_ (.A(_3082_),
    .B(_0395_),
    .X(_0415_));
 sky130_fd_sc_hd__buf_4 _3930_ (.A(_0415_),
    .X(_0416_));
 sky130_fd_sc_hd__clkbuf_4 _3931_ (.A(\egd_top.BitStream_buffer.BS_buffer[56] ),
    .X(_0417_));
 sky130_fd_sc_hd__nand2_1 _3932_ (.A(_0416_),
    .B(_0417_),
    .Y(_0418_));
 sky130_fd_sc_hd__and2_1 _3933_ (.A(_3061_),
    .B(_0395_),
    .X(_0419_));
 sky130_fd_sc_hd__clkbuf_4 _3934_ (.A(_0419_),
    .X(_0420_));
 sky130_fd_sc_hd__clkbuf_4 _3935_ (.A(\egd_top.BitStream_buffer.BS_buffer[58] ),
    .X(_0421_));
 sky130_fd_sc_hd__nand2_1 _3936_ (.A(_0420_),
    .B(_0421_),
    .Y(_0422_));
 sky130_fd_sc_hd__clkbuf_4 _3937_ (.A(\egd_top.BitStream_buffer.BS_buffer[57] ),
    .X(_0423_));
 sky130_fd_sc_hd__inv_2 _3938_ (.A(_0423_),
    .Y(_0424_));
 sky130_fd_sc_hd__nand2_1 _3939_ (.A(_3090_),
    .B(_0395_),
    .Y(_0425_));
 sky130_fd_sc_hd__buf_2 _3940_ (.A(_0425_),
    .X(_0426_));
 sky130_fd_sc_hd__or2_1 _3941_ (.A(_0424_),
    .B(_0426_),
    .X(_0427_));
 sky130_fd_sc_hd__o2111a_1 _3942_ (.A1(_0412_),
    .A2(_0414_),
    .B1(_0418_),
    .C1(_0422_),
    .D1(_0427_),
    .X(_0428_));
 sky130_fd_sc_hd__clkbuf_4 _3943_ (.A(\egd_top.BitStream_buffer.BS_buffer[50] ),
    .X(_0429_));
 sky130_fd_sc_hd__and2_1 _3944_ (.A(_3098_),
    .B(_2966_),
    .X(_0430_));
 sky130_fd_sc_hd__buf_1 _3945_ (.A(_0430_),
    .X(_0431_));
 sky130_fd_sc_hd__clkbuf_4 _3946_ (.A(_0431_),
    .X(_0432_));
 sky130_fd_sc_hd__clkbuf_4 _3947_ (.A(\egd_top.BitStream_buffer.BS_buffer[51] ),
    .X(_0433_));
 sky130_fd_sc_hd__and2_1 _3948_ (.A(_3103_),
    .B(_0395_),
    .X(_0434_));
 sky130_fd_sc_hd__buf_1 _3949_ (.A(_0434_),
    .X(_0435_));
 sky130_fd_sc_hd__clkbuf_4 _3950_ (.A(_0435_),
    .X(_0436_));
 sky130_fd_sc_hd__buf_4 _3951_ (.A(\egd_top.BitStream_buffer.BS_buffer[48] ),
    .X(_0437_));
 sky130_fd_sc_hd__inv_2 _3952_ (.A(_0437_),
    .Y(_0438_));
 sky130_fd_sc_hd__nand2_1 _3953_ (.A(_3109_),
    .B(_0395_),
    .Y(_0439_));
 sky130_fd_sc_hd__clkbuf_4 _3954_ (.A(_0439_),
    .X(_0440_));
 sky130_fd_sc_hd__and2_1 _3955_ (.A(_3112_),
    .B(_0395_),
    .X(_0441_));
 sky130_fd_sc_hd__clkbuf_4 _3956_ (.A(_0441_),
    .X(_0442_));
 sky130_fd_sc_hd__clkbuf_4 _3957_ (.A(\egd_top.BitStream_buffer.BS_buffer[49] ),
    .X(_0443_));
 sky130_fd_sc_hd__nand2_1 _3958_ (.A(_0442_),
    .B(_0443_),
    .Y(_0444_));
 sky130_fd_sc_hd__o21ai_1 _3959_ (.A1(_0438_),
    .A2(_0440_),
    .B1(_0444_),
    .Y(_0445_));
 sky130_fd_sc_hd__a221oi_1 _3960_ (.A1(_0429_),
    .A2(_0432_),
    .B1(_0433_),
    .B2(_0436_),
    .C1(_0445_),
    .Y(_0446_));
 sky130_fd_sc_hd__clkbuf_4 _3961_ (.A(\egd_top.BitStream_buffer.BS_buffer[60] ),
    .X(_0447_));
 sky130_fd_sc_hd__and2_1 _3962_ (.A(_3158_),
    .B(_2966_),
    .X(_0448_));
 sky130_fd_sc_hd__buf_1 _3963_ (.A(_0448_),
    .X(_0449_));
 sky130_fd_sc_hd__clkbuf_4 _3964_ (.A(_0449_),
    .X(_0450_));
 sky130_fd_sc_hd__clkbuf_4 _3965_ (.A(\egd_top.BitStream_buffer.BS_buffer[61] ),
    .X(_0451_));
 sky130_fd_sc_hd__and2_1 _3966_ (.A(_3153_),
    .B(_2966_),
    .X(_0452_));
 sky130_fd_sc_hd__buf_1 _3967_ (.A(_0452_),
    .X(_0453_));
 sky130_fd_sc_hd__clkbuf_4 _3968_ (.A(_0453_),
    .X(_0454_));
 sky130_fd_sc_hd__clkbuf_4 _3969_ (.A(\egd_top.BitStream_buffer.BS_buffer[63] ),
    .X(_0455_));
 sky130_fd_sc_hd__inv_2 _3970_ (.A(_0455_),
    .Y(_0456_));
 sky130_fd_sc_hd__inv_2 _3971_ (.A(_2967_),
    .Y(_0457_));
 sky130_fd_sc_hd__clkbuf_4 _3972_ (.A(_0457_),
    .X(_0458_));
 sky130_fd_sc_hd__and2_1 _3973_ (.A(_3145_),
    .B(_0395_),
    .X(_0459_));
 sky130_fd_sc_hd__clkbuf_4 _3974_ (.A(_0459_),
    .X(_0460_));
 sky130_fd_sc_hd__clkbuf_4 _3975_ (.A(\egd_top.BitStream_buffer.BS_buffer[62] ),
    .X(_0461_));
 sky130_fd_sc_hd__nand2_1 _3976_ (.A(_0460_),
    .B(_0461_),
    .Y(_0462_));
 sky130_fd_sc_hd__o21ai_1 _3977_ (.A1(_0456_),
    .A2(_0458_),
    .B1(_0462_),
    .Y(_0463_));
 sky130_fd_sc_hd__a221oi_1 _3978_ (.A1(_0447_),
    .A2(_0450_),
    .B1(_0451_),
    .B2(_0454_),
    .C1(_0463_),
    .Y(_0464_));
 sky130_fd_sc_hd__and4_1 _3979_ (.A(_0410_),
    .B(_0428_),
    .C(_0446_),
    .D(_0464_),
    .X(_0465_));
 sky130_fd_sc_hd__and2_1 _3980_ (.A(_0393_),
    .B(_0465_),
    .X(_0466_));
 sky130_fd_sc_hd__clkbuf_4 _3981_ (.A(\egd_top.BitStream_buffer.BS_buffer[24] ),
    .X(_0467_));
 sky130_fd_sc_hd__inv_2 _3982_ (.A(_0467_),
    .Y(_0468_));
 sky130_fd_sc_hd__and3_1 _3983_ (.A(_2965_),
    .B(_3063_),
    .C(\egd_top.BitStream_buffer.pc[4] ),
    .X(_0469_));
 sky130_fd_sc_hd__buf_2 _3984_ (.A(_0469_),
    .X(_0470_));
 sky130_fd_sc_hd__nand2_1 _3985_ (.A(_3082_),
    .B(_0470_),
    .Y(_0471_));
 sky130_fd_sc_hd__clkbuf_4 _3986_ (.A(_0471_),
    .X(_0472_));
 sky130_fd_sc_hd__and2_1 _3987_ (.A(_3090_),
    .B(_0470_),
    .X(_0473_));
 sky130_fd_sc_hd__buf_4 _3988_ (.A(_0473_),
    .X(_0474_));
 sky130_fd_sc_hd__clkbuf_4 _3989_ (.A(\egd_top.BitStream_buffer.BS_buffer[25] ),
    .X(_0475_));
 sky130_fd_sc_hd__nand2_1 _3990_ (.A(_0474_),
    .B(_0475_),
    .Y(_0476_));
 sky130_fd_sc_hd__and2_2 _3991_ (.A(_3061_),
    .B(_0469_),
    .X(_0477_));
 sky130_fd_sc_hd__clkbuf_4 _3992_ (.A(_0477_),
    .X(_0478_));
 sky130_fd_sc_hd__clkbuf_4 _3993_ (.A(\egd_top.BitStream_buffer.BS_buffer[26] ),
    .X(_0479_));
 sky130_fd_sc_hd__and2_1 _3994_ (.A(_3072_),
    .B(_0469_),
    .X(_0480_));
 sky130_fd_sc_hd__clkbuf_4 _3995_ (.A(_0480_),
    .X(_0481_));
 sky130_fd_sc_hd__clkbuf_4 _3996_ (.A(\egd_top.BitStream_buffer.BS_buffer[27] ),
    .X(_0482_));
 sky130_fd_sc_hd__a22o_1 _3997_ (.A1(_0478_),
    .A2(_0479_),
    .B1(_0481_),
    .B2(_0482_),
    .X(_0483_));
 sky130_fd_sc_hd__inv_2 _3998_ (.A(_0483_),
    .Y(_0484_));
 sky130_fd_sc_hd__o211a_1 _3999_ (.A1(_0468_),
    .A2(_0472_),
    .B1(_0476_),
    .C1(_0484_),
    .X(_0485_));
 sky130_fd_sc_hd__and2_1 _4000_ (.A(_3109_),
    .B(_0470_),
    .X(_0486_));
 sky130_fd_sc_hd__buf_1 _4001_ (.A(_0486_),
    .X(_0487_));
 sky130_fd_sc_hd__clkbuf_4 _4002_ (.A(_0487_),
    .X(_0488_));
 sky130_fd_sc_hd__clkbuf_4 _4003_ (.A(\egd_top.BitStream_buffer.BS_buffer[17] ),
    .X(_0489_));
 sky130_fd_sc_hd__and2_1 _4004_ (.A(_3112_),
    .B(_0470_),
    .X(_0490_));
 sky130_fd_sc_hd__buf_1 _4005_ (.A(_0490_),
    .X(_0491_));
 sky130_fd_sc_hd__clkbuf_4 _4006_ (.A(_0491_),
    .X(_0492_));
 sky130_fd_sc_hd__clkbuf_4 _4007_ (.A(\egd_top.BitStream_buffer.BS_buffer[18] ),
    .X(_0493_));
 sky130_fd_sc_hd__inv_2 _4008_ (.A(_0493_),
    .Y(_0494_));
 sky130_fd_sc_hd__nand2_1 _4009_ (.A(_3098_),
    .B(_0470_),
    .Y(_0495_));
 sky130_fd_sc_hd__clkbuf_4 _4010_ (.A(_0495_),
    .X(_0496_));
 sky130_fd_sc_hd__and2_1 _4011_ (.A(_3103_),
    .B(_0470_),
    .X(_0497_));
 sky130_fd_sc_hd__clkbuf_4 _4012_ (.A(_0497_),
    .X(_0498_));
 sky130_fd_sc_hd__clkbuf_4 _4013_ (.A(\egd_top.BitStream_buffer.BS_buffer[19] ),
    .X(_0499_));
 sky130_fd_sc_hd__nand2_1 _4014_ (.A(_0498_),
    .B(_0499_),
    .Y(_0500_));
 sky130_fd_sc_hd__o21ai_1 _4015_ (.A1(_0494_),
    .A2(_0496_),
    .B1(_0500_),
    .Y(_0501_));
 sky130_fd_sc_hd__a221oi_1 _4016_ (.A1(\egd_top.BitStream_buffer.BS_buffer[16] ),
    .A2(_0488_),
    .B1(_0489_),
    .B2(_0492_),
    .C1(_0501_),
    .Y(_0502_));
 sky130_fd_sc_hd__clkbuf_4 _4017_ (.A(\egd_top.BitStream_buffer.BS_buffer[23] ),
    .X(_0503_));
 sky130_fd_sc_hd__inv_2 _4018_ (.A(_0503_),
    .Y(_0504_));
 sky130_fd_sc_hd__nand2_1 _4019_ (.A(_3122_),
    .B(_0470_),
    .Y(_0505_));
 sky130_fd_sc_hd__clkbuf_4 _4020_ (.A(_0505_),
    .X(_0506_));
 sky130_fd_sc_hd__and2_1 _4021_ (.A(_3131_),
    .B(_0470_),
    .X(_0507_));
 sky130_fd_sc_hd__clkbuf_4 _4022_ (.A(_0507_),
    .X(_0508_));
 sky130_fd_sc_hd__clkbuf_4 _4023_ (.A(\egd_top.BitStream_buffer.BS_buffer[22] ),
    .X(_0509_));
 sky130_fd_sc_hd__nand2_1 _4024_ (.A(_0508_),
    .B(_0509_),
    .Y(_0510_));
 sky130_fd_sc_hd__and2_1 _4025_ (.A(_3126_),
    .B(_0470_),
    .X(_0511_));
 sky130_fd_sc_hd__clkbuf_4 _4026_ (.A(_0511_),
    .X(_0512_));
 sky130_fd_sc_hd__clkbuf_4 _4027_ (.A(\egd_top.BitStream_buffer.BS_buffer[20] ),
    .X(_0513_));
 sky130_fd_sc_hd__nand2_1 _4028_ (.A(_0512_),
    .B(_0513_),
    .Y(_0514_));
 sky130_fd_sc_hd__clkbuf_4 _4029_ (.A(\egd_top.BitStream_buffer.BS_buffer[21] ),
    .X(_0515_));
 sky130_fd_sc_hd__inv_2 _4030_ (.A(_0515_),
    .Y(_0516_));
 sky130_fd_sc_hd__nand2_1 _4031_ (.A(_3139_),
    .B(_0470_),
    .Y(_0517_));
 sky130_fd_sc_hd__buf_2 _4032_ (.A(_0517_),
    .X(_0518_));
 sky130_fd_sc_hd__or2_1 _4033_ (.A(_0516_),
    .B(_0518_),
    .X(_0519_));
 sky130_fd_sc_hd__o2111a_1 _4034_ (.A1(_0504_),
    .A2(_0506_),
    .B1(_0510_),
    .C1(_0514_),
    .D1(_0519_),
    .X(_0520_));
 sky130_fd_sc_hd__clkbuf_4 _4035_ (.A(\egd_top.BitStream_buffer.BS_buffer[30] ),
    .X(_0521_));
 sky130_fd_sc_hd__and2_1 _4036_ (.A(_3145_),
    .B(_0469_),
    .X(_0522_));
 sky130_fd_sc_hd__buf_1 _4037_ (.A(_0522_),
    .X(_0523_));
 sky130_fd_sc_hd__clkbuf_4 _4038_ (.A(_0523_),
    .X(_0524_));
 sky130_fd_sc_hd__clkbuf_4 _4039_ (.A(\egd_top.BitStream_buffer.BS_buffer[31] ),
    .X(_0525_));
 sky130_fd_sc_hd__and2_1 _4040_ (.A(_2964_),
    .B(_0469_),
    .X(_0526_));
 sky130_fd_sc_hd__buf_1 _4041_ (.A(_0526_),
    .X(_0527_));
 sky130_fd_sc_hd__clkbuf_4 _4042_ (.A(_0527_),
    .X(_0528_));
 sky130_fd_sc_hd__and2_1 _4043_ (.A(_3153_),
    .B(_0470_),
    .X(_0529_));
 sky130_fd_sc_hd__clkbuf_4 _4044_ (.A(_0529_),
    .X(_0530_));
 sky130_fd_sc_hd__clkbuf_4 _4045_ (.A(\egd_top.BitStream_buffer.BS_buffer[29] ),
    .X(_0531_));
 sky130_fd_sc_hd__nand2_1 _4046_ (.A(_0530_),
    .B(_0531_),
    .Y(_0532_));
 sky130_fd_sc_hd__and2_1 _4047_ (.A(_3158_),
    .B(_0470_),
    .X(_0533_));
 sky130_fd_sc_hd__clkbuf_4 _4048_ (.A(_0533_),
    .X(_0534_));
 sky130_fd_sc_hd__clkbuf_4 _4049_ (.A(\egd_top.BitStream_buffer.BS_buffer[28] ),
    .X(_0535_));
 sky130_fd_sc_hd__nand2_1 _4050_ (.A(_0534_),
    .B(_0535_),
    .Y(_0536_));
 sky130_fd_sc_hd__nand2_1 _4051_ (.A(_0532_),
    .B(_0536_),
    .Y(_0537_));
 sky130_fd_sc_hd__a221oi_1 _4052_ (.A1(_0521_),
    .A2(_0524_),
    .B1(_0525_),
    .B2(_0528_),
    .C1(_0537_),
    .Y(_0538_));
 sky130_fd_sc_hd__and4_1 _4053_ (.A(_0485_),
    .B(_0502_),
    .C(_0520_),
    .D(_0538_),
    .X(_0539_));
 sky130_fd_sc_hd__clkbuf_4 _4054_ (.A(\egd_top.BitStream_buffer.BS_buffer[5] ),
    .X(_0540_));
 sky130_fd_sc_hd__inv_2 _4055_ (.A(_0540_),
    .Y(_0541_));
 sky130_fd_sc_hd__and3_1 _4056_ (.A(_2965_),
    .B(_3062_),
    .C(_3063_),
    .X(_0542_));
 sky130_fd_sc_hd__clkbuf_4 _4057_ (.A(_0542_),
    .X(_0543_));
 sky130_fd_sc_hd__nand2_1 _4058_ (.A(_3139_),
    .B(_0543_),
    .Y(_0544_));
 sky130_fd_sc_hd__clkbuf_4 _4059_ (.A(_0544_),
    .X(_0545_));
 sky130_fd_sc_hd__and2_1 _4060_ (.A(_3131_),
    .B(_0543_),
    .X(_0546_));
 sky130_fd_sc_hd__clkbuf_4 _4061_ (.A(_0546_),
    .X(_0547_));
 sky130_fd_sc_hd__clkbuf_4 _4062_ (.A(\egd_top.BitStream_buffer.BS_buffer[6] ),
    .X(_0548_));
 sky130_fd_sc_hd__nand2_1 _4063_ (.A(_0547_),
    .B(_0548_),
    .Y(_0549_));
 sky130_fd_sc_hd__and2_1 _4064_ (.A(_3126_),
    .B(_0543_),
    .X(_0550_));
 sky130_fd_sc_hd__clkbuf_4 _4065_ (.A(_0550_),
    .X(_0551_));
 sky130_fd_sc_hd__clkbuf_4 _4066_ (.A(\egd_top.BitStream_buffer.BS_buffer[4] ),
    .X(_0552_));
 sky130_fd_sc_hd__nand2_1 _4067_ (.A(_0551_),
    .B(_0552_),
    .Y(_0553_));
 sky130_fd_sc_hd__inv_2 _4068_ (.A(\egd_top.BitStream_buffer.BS_buffer[7] ),
    .Y(_0554_));
 sky130_fd_sc_hd__nand2_1 _4069_ (.A(_3122_),
    .B(_0543_),
    .Y(_0555_));
 sky130_fd_sc_hd__clkbuf_4 _4070_ (.A(_0555_),
    .X(_0556_));
 sky130_fd_sc_hd__or2_1 _4071_ (.A(_0554_),
    .B(_0556_),
    .X(_0557_));
 sky130_fd_sc_hd__o2111a_1 _4072_ (.A1(_0541_),
    .A2(_0545_),
    .B1(_0549_),
    .C1(_0553_),
    .D1(_0557_),
    .X(_0558_));
 sky130_fd_sc_hd__inv_2 _4073_ (.A(\egd_top.BitStream_buffer.BS_buffer[11] ),
    .Y(_0559_));
 sky130_fd_sc_hd__nand2_1 _4074_ (.A(_3072_),
    .B(_0543_),
    .Y(_0560_));
 sky130_fd_sc_hd__clkbuf_4 _4075_ (.A(_0560_),
    .X(_0561_));
 sky130_fd_sc_hd__and2_1 _4076_ (.A(_3061_),
    .B(_0543_),
    .X(_0562_));
 sky130_fd_sc_hd__clkbuf_4 _4077_ (.A(_0562_),
    .X(_0563_));
 sky130_fd_sc_hd__nand2_1 _4078_ (.A(_0563_),
    .B(\egd_top.BitStream_buffer.BS_buffer[10] ),
    .Y(_0564_));
 sky130_fd_sc_hd__and2_1 _4079_ (.A(_3082_),
    .B(_0543_),
    .X(_0565_));
 sky130_fd_sc_hd__buf_4 _4080_ (.A(_0565_),
    .X(_0566_));
 sky130_fd_sc_hd__nand2_1 _4081_ (.A(_0566_),
    .B(\egd_top.BitStream_buffer.BS_buffer[8] ),
    .Y(_0567_));
 sky130_fd_sc_hd__inv_2 _4082_ (.A(\egd_top.BitStream_buffer.BS_buffer[9] ),
    .Y(_0568_));
 sky130_fd_sc_hd__nand2_1 _4083_ (.A(_3090_),
    .B(_0542_),
    .Y(_0569_));
 sky130_fd_sc_hd__buf_2 _4084_ (.A(_0569_),
    .X(_0570_));
 sky130_fd_sc_hd__or2_1 _4085_ (.A(_0568_),
    .B(_0570_),
    .X(_0571_));
 sky130_fd_sc_hd__o2111a_1 _4086_ (.A1(_0559_),
    .A2(_0561_),
    .B1(_0564_),
    .C1(_0567_),
    .D1(_0571_),
    .X(_0572_));
 sky130_fd_sc_hd__clkbuf_4 _4087_ (.A(\egd_top.BitStream_buffer.BS_buffer[2] ),
    .X(_0573_));
 sky130_fd_sc_hd__inv_2 _4088_ (.A(_0573_),
    .Y(_0574_));
 sky130_fd_sc_hd__nand2_1 _4089_ (.A(_3098_),
    .B(_0543_),
    .Y(_0575_));
 sky130_fd_sc_hd__clkbuf_4 _4090_ (.A(_0575_),
    .X(_0576_));
 sky130_fd_sc_hd__clkbuf_4 _4091_ (.A(\egd_top.BitStream_buffer.BS_buffer[1] ),
    .X(_0577_));
 sky130_fd_sc_hd__inv_2 _4092_ (.A(_0577_),
    .Y(_0578_));
 sky130_fd_sc_hd__nand2_1 _4093_ (.A(_3112_),
    .B(_0543_),
    .Y(_0579_));
 sky130_fd_sc_hd__clkbuf_4 _4094_ (.A(_0579_),
    .X(_0580_));
 sky130_fd_sc_hd__clkbuf_4 _4095_ (.A(\egd_top.BitStream_buffer.BS_buffer[3] ),
    .X(_0581_));
 sky130_fd_sc_hd__inv_2 _4096_ (.A(_0581_),
    .Y(_0582_));
 sky130_fd_sc_hd__nand2_1 _4097_ (.A(_3103_),
    .B(_0542_),
    .Y(_0583_));
 sky130_fd_sc_hd__buf_2 _4098_ (.A(_0583_),
    .X(_0584_));
 sky130_fd_sc_hd__or2_1 _4099_ (.A(_0582_),
    .B(_0584_),
    .X(_0585_));
 sky130_fd_sc_hd__o221a_1 _4100_ (.A1(_0574_),
    .A2(_0576_),
    .B1(_0578_),
    .B2(_0580_),
    .C1(_0585_),
    .X(_0586_));
 sky130_fd_sc_hd__and2_1 _4101_ (.A(_3145_),
    .B(_0542_),
    .X(_0587_));
 sky130_fd_sc_hd__buf_1 _4102_ (.A(_0587_),
    .X(_0588_));
 sky130_fd_sc_hd__clkbuf_4 _4103_ (.A(_0588_),
    .X(_0589_));
 sky130_fd_sc_hd__and2_1 _4104_ (.A(_2964_),
    .B(_0542_),
    .X(_0590_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _4105_ (.A(_0590_),
    .X(_0591_));
 sky130_fd_sc_hd__clkbuf_4 _4106_ (.A(_0591_),
    .X(_0592_));
 sky130_fd_sc_hd__inv_2 _4107_ (.A(\egd_top.BitStream_buffer.BS_buffer[12] ),
    .Y(_0593_));
 sky130_fd_sc_hd__nand2_1 _4108_ (.A(_3158_),
    .B(_0543_),
    .Y(_0594_));
 sky130_fd_sc_hd__clkbuf_4 _4109_ (.A(_0594_),
    .X(_0595_));
 sky130_fd_sc_hd__inv_2 _4110_ (.A(\egd_top.BitStream_buffer.BS_buffer[13] ),
    .Y(_0596_));
 sky130_fd_sc_hd__nand2_1 _4111_ (.A(_3153_),
    .B(_0543_),
    .Y(_0597_));
 sky130_fd_sc_hd__clkbuf_4 _4112_ (.A(_0597_),
    .X(_0598_));
 sky130_fd_sc_hd__o22ai_1 _4113_ (.A1(_0593_),
    .A2(_0595_),
    .B1(_0596_),
    .B2(_0598_),
    .Y(_0599_));
 sky130_fd_sc_hd__a221oi_1 _4114_ (.A1(\egd_top.BitStream_buffer.BS_buffer[14] ),
    .A2(_0589_),
    .B1(\egd_top.BitStream_buffer.BS_buffer[15] ),
    .B2(_0592_),
    .C1(_0599_),
    .Y(_0600_));
 sky130_fd_sc_hd__and4_1 _4115_ (.A(_0558_),
    .B(_0572_),
    .C(_0586_),
    .D(_0600_),
    .X(_0601_));
 sky130_fd_sc_hd__and3_1 _4116_ (.A(_0466_),
    .B(_0539_),
    .C(_0601_),
    .X(_0602_));
 sky130_fd_sc_hd__o41a_1 _4117_ (.A1(\egd_top.BitStream_buffer.pc[2] ),
    .A2(\egd_top.BitStream_buffer.pc[3] ),
    .A3(\egd_top.BitStream_buffer.pc[1] ),
    .A4(_2962_),
    .B1(_0543_),
    .X(_0603_));
 sky130_fd_sc_hd__and4b_1 _4118_ (.A_N(_0603_),
    .B(_2965_),
    .C(_3062_),
    .D(_3063_),
    .X(_0604_));
 sky130_fd_sc_hd__buf_1 _4119_ (.A(_0604_),
    .X(_0605_));
 sky130_fd_sc_hd__clkbuf_4 _4120_ (.A(_0605_),
    .X(_0606_));
 sky130_fd_sc_hd__clkbuf_4 _4121_ (.A(\egd_top.BitStream_buffer.BS_buffer[0] ),
    .X(_0607_));
 sky130_fd_sc_hd__nand2_1 _4122_ (.A(_0606_),
    .B(_0607_),
    .Y(_0608_));
 sky130_fd_sc_hd__nand3_1 _4123_ (.A(_0322_),
    .B(_0602_),
    .C(_0608_),
    .Y(_0609_));
 sky130_fd_sc_hd__o21a_1 _4124_ (.A1(\egd_top.BitStream_buffer.BitStream_buffer_output[15] ),
    .A2(_2997_),
    .B1(_2989_),
    .X(_0610_));
 sky130_fd_sc_hd__o21a_1 _4125_ (.A1(_3056_),
    .A2(_0609_),
    .B1(_0610_),
    .X(_0297_));
 sky130_fd_sc_hd__inv_2 _4126_ (.A(_3057_),
    .Y(_0611_));
 sky130_fd_sc_hd__o22ai_1 _4127_ (.A1(_3086_),
    .A2(_3084_),
    .B1(_0611_),
    .B2(_3092_),
    .Y(_0612_));
 sky130_fd_sc_hd__a221oi_1 _4128_ (.A1(_3069_),
    .A2(_3068_),
    .B1(_3161_),
    .B2(_3075_),
    .C1(_0612_),
    .Y(_0613_));
 sky130_fd_sc_hd__inv_2 _4129_ (.A(_3115_),
    .Y(_0614_));
 sky130_fd_sc_hd__nand2_1 _4130_ (.A(_3114_),
    .B(_3095_),
    .Y(_0615_));
 sky130_fd_sc_hd__o21ai_1 _4131_ (.A1(_0614_),
    .A2(_3111_),
    .B1(_0615_),
    .Y(_0616_));
 sky130_fd_sc_hd__a221oi_1 _4132_ (.A1(_3102_),
    .A2(_3101_),
    .B1(_3129_),
    .B2(_3106_),
    .C1(_0616_),
    .Y(_0617_));
 sky130_fd_sc_hd__nand2_1 _4133_ (.A(_3128_),
    .B(_3136_),
    .Y(_0618_));
 sky130_fd_sc_hd__nand2_1 _4134_ (.A(_3133_),
    .B(_3119_),
    .Y(_0619_));
 sky130_fd_sc_hd__inv_2 _4135_ (.A(_3134_),
    .Y(_0620_));
 sky130_fd_sc_hd__or2_1 _4136_ (.A(_0620_),
    .B(_3141_),
    .X(_0621_));
 sky130_fd_sc_hd__o2111a_1 _4137_ (.A1(_3077_),
    .A2(_3124_),
    .B1(_0618_),
    .C1(_0619_),
    .D1(_0621_),
    .X(_0622_));
 sky130_fd_sc_hd__nand2_1 _4138_ (.A(_3155_),
    .B(_3144_),
    .Y(_0623_));
 sky130_fd_sc_hd__nand2_1 _4139_ (.A(_3160_),
    .B(_3156_),
    .Y(_0624_));
 sky130_fd_sc_hd__nand2_1 _4140_ (.A(_0623_),
    .B(_0624_),
    .Y(_0625_));
 sky130_fd_sc_hd__a221oi_1 _4141_ (.A1(_3149_),
    .A2(_3148_),
    .B1(_3255_),
    .B2(_3152_),
    .C1(_0625_),
    .Y(_0626_));
 sky130_fd_sc_hd__and4_1 _4142_ (.A(_0613_),
    .B(_0617_),
    .C(_0622_),
    .D(_0626_),
    .X(_0627_));
 sky130_fd_sc_hd__inv_2 _4143_ (.A(\egd_top.BitStream_buffer.BS_buffer[118] ),
    .Y(_0628_));
 sky130_fd_sc_hd__o22ai_1 _4144_ (.A1(_3177_),
    .A2(_3176_),
    .B1(_0628_),
    .B2(_3179_),
    .Y(_0629_));
 sky130_fd_sc_hd__a221oi_1 _4145_ (.A1(_3028_),
    .A2(_3170_),
    .B1(_3031_),
    .B2(_3173_),
    .C1(_0629_),
    .Y(_0630_));
 sky130_fd_sc_hd__nand2_1 _4146_ (.A(_3192_),
    .B(_3040_),
    .Y(_0631_));
 sky130_fd_sc_hd__o21ai_1 _4147_ (.A1(_3216_),
    .A2(_3190_),
    .B1(_0631_),
    .Y(_0632_));
 sky130_fd_sc_hd__a221oi_1 _4148_ (.A1(_3034_),
    .A2(_3184_),
    .B1(_3037_),
    .B2(_3187_),
    .C1(_0632_),
    .Y(_0633_));
 sky130_fd_sc_hd__inv_2 _4149_ (.A(\egd_top.BitStream_buffer.BS_buffer[113] ),
    .Y(_0634_));
 sky130_fd_sc_hd__nand2_1 _4150_ (.A(_3206_),
    .B(_3013_),
    .Y(_0635_));
 sky130_fd_sc_hd__o21ai_1 _4151_ (.A1(_0634_),
    .A2(_3204_),
    .B1(_0635_),
    .Y(_0636_));
 sky130_fd_sc_hd__a221oi_1 _4152_ (.A1(_3016_),
    .A2(_3198_),
    .B1(_3019_),
    .B2(_3201_),
    .C1(_0636_),
    .Y(_0637_));
 sky130_fd_sc_hd__inv_2 _4153_ (.A(_3050_),
    .Y(_0638_));
 sky130_fd_sc_hd__o22ai_1 _4154_ (.A1(_3219_),
    .A2(_3218_),
    .B1(_0638_),
    .B2(_3221_),
    .Y(_0639_));
 sky130_fd_sc_hd__a221oi_1 _4155_ (.A1(_3053_),
    .A2(_3212_),
    .B1(_0607_),
    .B2(_3215_),
    .C1(_0639_),
    .Y(_0640_));
 sky130_fd_sc_hd__and4_1 _4156_ (.A(_0630_),
    .B(_0633_),
    .C(_0637_),
    .D(_0640_),
    .X(_0641_));
 sky130_fd_sc_hd__inv_2 _4157_ (.A(\egd_top.BitStream_buffer.BS_buffer[90] ),
    .Y(_0642_));
 sky130_fd_sc_hd__o22ai_1 _4158_ (.A1(_3239_),
    .A2(_3238_),
    .B1(_0642_),
    .B2(_3241_),
    .Y(_0643_));
 sky130_fd_sc_hd__a221oi_1 _4159_ (.A1(_3232_),
    .A2(_3231_),
    .B1(_3286_),
    .B2(_3235_),
    .C1(_0643_),
    .Y(_0644_));
 sky130_fd_sc_hd__nand2_1 _4160_ (.A(_3246_),
    .B(_3259_),
    .Y(_0645_));
 sky130_fd_sc_hd__clkbuf_4 _4161_ (.A(\egd_top.BitStream_buffer.BS_buffer[84] ),
    .X(_0646_));
 sky130_fd_sc_hd__nand2_1 _4162_ (.A(_3250_),
    .B(_0646_),
    .Y(_0647_));
 sky130_fd_sc_hd__nand2_1 _4163_ (.A(_3254_),
    .B(_3247_),
    .Y(_0648_));
 sky130_fd_sc_hd__nand2_1 _4164_ (.A(_3258_),
    .B(_3251_),
    .Y(_0649_));
 sky130_fd_sc_hd__and4_1 _4165_ (.A(_0645_),
    .B(_0647_),
    .C(_0648_),
    .D(_0649_),
    .X(_0650_));
 sky130_fd_sc_hd__inv_2 _4166_ (.A(\egd_top.BitStream_buffer.BS_buffer[86] ),
    .Y(_0651_));
 sky130_fd_sc_hd__o22ai_1 _4167_ (.A1(_3266_),
    .A2(_3264_),
    .B1(_0651_),
    .B2(_3268_),
    .Y(_0652_));
 sky130_fd_sc_hd__clkbuf_4 _4168_ (.A(\egd_top.BitStream_buffer.BS_buffer[88] ),
    .X(_0653_));
 sky130_fd_sc_hd__a22o_1 _4169_ (.A1(_3271_),
    .A2(_3275_),
    .B1(_3274_),
    .B2(_0653_),
    .X(_0654_));
 sky130_fd_sc_hd__nor2_1 _4170_ (.A(_0652_),
    .B(_0654_),
    .Y(_0655_));
 sky130_fd_sc_hd__inv_2 _4171_ (.A(_3278_),
    .Y(_0656_));
 sky130_fd_sc_hd__o22ai_1 _4172_ (.A1(_3291_),
    .A2(_3289_),
    .B1(_0656_),
    .B2(_3293_),
    .Y(_0657_));
 sky130_fd_sc_hd__a221oi_1 _4173_ (.A1(_3282_),
    .A2(_3281_),
    .B1(_3318_),
    .B2(_3285_),
    .C1(_0657_),
    .Y(_0658_));
 sky130_fd_sc_hd__and4_1 _4174_ (.A(_0644_),
    .B(_0650_),
    .C(_0655_),
    .D(_0658_),
    .X(_0659_));
 sky130_fd_sc_hd__nand2_1 _4175_ (.A(_3309_),
    .B(_3297_),
    .Y(_0660_));
 sky130_fd_sc_hd__nand2_1 _4176_ (.A(_3313_),
    .B(_3310_),
    .Y(_0661_));
 sky130_fd_sc_hd__nand2_1 _4177_ (.A(_0660_),
    .B(_0661_),
    .Y(_0662_));
 sky130_fd_sc_hd__a221oi_1 _4178_ (.A1(_3304_),
    .A2(_3303_),
    .B1(_3353_),
    .B2(_3307_),
    .C1(_0662_),
    .Y(_0663_));
 sky130_fd_sc_hd__nand2_1 _4179_ (.A(_3326_),
    .B(_3341_),
    .Y(_0664_));
 sky130_fd_sc_hd__nand2_1 _4180_ (.A(_3330_),
    .B(_3327_),
    .Y(_0665_));
 sky130_fd_sc_hd__nand2_1 _4181_ (.A(_0664_),
    .B(_0665_),
    .Y(_0666_));
 sky130_fd_sc_hd__a221oi_1 _4182_ (.A1(_3322_),
    .A2(_3321_),
    .B1(_3331_),
    .B2(_3324_),
    .C1(_0666_),
    .Y(_0667_));
 sky130_fd_sc_hd__inv_2 _4183_ (.A(\egd_top.BitStream_buffer.BS_buffer[104] ),
    .Y(_0668_));
 sky130_fd_sc_hd__nand2_1 _4184_ (.A(_3340_),
    .B(_3347_),
    .Y(_0669_));
 sky130_fd_sc_hd__nand2_1 _4185_ (.A(_3344_),
    .B(_3335_),
    .Y(_0670_));
 sky130_fd_sc_hd__inv_2 _4186_ (.A(_3345_),
    .Y(_0671_));
 sky130_fd_sc_hd__or2_1 _4187_ (.A(_0671_),
    .B(_3350_),
    .X(_0672_));
 sky130_fd_sc_hd__o2111a_1 _4188_ (.A1(_0668_),
    .A2(_3338_),
    .B1(_0669_),
    .C1(_0670_),
    .D1(_0672_),
    .X(_0673_));
 sky130_fd_sc_hd__clkbuf_4 _4189_ (.A(\egd_top.BitStream_buffer.BS_buffer[110] ),
    .X(_0674_));
 sky130_fd_sc_hd__clkbuf_4 _4190_ (.A(\egd_top.BitStream_buffer.BS_buffer[111] ),
    .X(_0675_));
 sky130_fd_sc_hd__nand2_1 _4191_ (.A(_3365_),
    .B(_0675_),
    .Y(_0676_));
 sky130_fd_sc_hd__o21ai_1 _4192_ (.A1(_3202_),
    .A2(_3363_),
    .B1(_0676_),
    .Y(_0677_));
 sky130_fd_sc_hd__a221oi_1 _4193_ (.A1(_3357_),
    .A2(_3356_),
    .B1(_0674_),
    .B2(_3360_),
    .C1(_0677_),
    .Y(_0678_));
 sky130_fd_sc_hd__and4_1 _4194_ (.A(_0663_),
    .B(_0667_),
    .C(_0673_),
    .D(_0678_),
    .X(_0679_));
 sky130_fd_sc_hd__and4_1 _4195_ (.A(_0627_),
    .B(_0641_),
    .C(_0659_),
    .D(_0679_),
    .X(_0680_));
 sky130_fd_sc_hd__nand2_1 _4196_ (.A(_0334_),
    .B(_0323_),
    .Y(_0681_));
 sky130_fd_sc_hd__nand2_1 _4197_ (.A(_0338_),
    .B(_0335_),
    .Y(_0682_));
 sky130_fd_sc_hd__nand2_1 _4198_ (.A(_0681_),
    .B(_0682_),
    .Y(_0683_));
 sky130_fd_sc_hd__a221oi_1 _4199_ (.A1(_0329_),
    .A2(_0328_),
    .B1(_0376_),
    .B2(_0332_),
    .C1(_0683_),
    .Y(_0684_));
 sky130_fd_sc_hd__inv_2 _4200_ (.A(\egd_top.BitStream_buffer.BS_buffer[38] ),
    .Y(_0685_));
 sky130_fd_sc_hd__o22ai_1 _4201_ (.A1(_0347_),
    .A2(_0345_),
    .B1(_0685_),
    .B2(_0349_),
    .Y(_0686_));
 sky130_fd_sc_hd__a22o_1 _4202_ (.A1(_0352_),
    .A2(_0356_),
    .B1(_0355_),
    .B2(_0339_),
    .X(_0687_));
 sky130_fd_sc_hd__nor2_1 _4203_ (.A(_0686_),
    .B(_0687_),
    .Y(_0688_));
 sky130_fd_sc_hd__clkbuf_4 _4204_ (.A(\egd_top.BitStream_buffer.BS_buffer[34] ),
    .X(_0689_));
 sky130_fd_sc_hd__inv_2 _4205_ (.A(\egd_top.BitStream_buffer.BS_buffer[35] ),
    .Y(_0690_));
 sky130_fd_sc_hd__clkbuf_4 _4206_ (.A(\egd_top.BitStream_buffer.BS_buffer[36] ),
    .X(_0691_));
 sky130_fd_sc_hd__nand2_1 _4207_ (.A(_0371_),
    .B(_0691_),
    .Y(_0692_));
 sky130_fd_sc_hd__o21ai_1 _4208_ (.A1(_0690_),
    .A2(_0369_),
    .B1(_0692_),
    .Y(_0693_));
 sky130_fd_sc_hd__a221oi_1 _4209_ (.A1(_0363_),
    .A2(_0362_),
    .B1(_0689_),
    .B2(_0366_),
    .C1(_0693_),
    .Y(_0694_));
 sky130_fd_sc_hd__clkbuf_4 _4210_ (.A(\egd_top.BitStream_buffer.BS_buffer[47] ),
    .X(_0695_));
 sky130_fd_sc_hd__nand2_1 _4211_ (.A(_0388_),
    .B(_0695_),
    .Y(_0696_));
 sky130_fd_sc_hd__o21ai_1 _4212_ (.A1(_0438_),
    .A2(_0386_),
    .B1(_0696_),
    .Y(_0697_));
 sky130_fd_sc_hd__a221oi_1 _4213_ (.A1(_0380_),
    .A2(_0379_),
    .B1(_0389_),
    .B2(_0383_),
    .C1(_0697_),
    .Y(_0698_));
 sky130_fd_sc_hd__and4_1 _4214_ (.A(_0684_),
    .B(_0688_),
    .C(_0694_),
    .D(_0698_),
    .X(_0699_));
 sky130_fd_sc_hd__inv_2 _4215_ (.A(\egd_top.BitStream_buffer.BS_buffer[54] ),
    .Y(_0700_));
 sky130_fd_sc_hd__clkbuf_4 _4216_ (.A(\egd_top.BitStream_buffer.BS_buffer[55] ),
    .X(_0701_));
 sky130_fd_sc_hd__nand2_1 _4217_ (.A(_0399_),
    .B(_0701_),
    .Y(_0702_));
 sky130_fd_sc_hd__clkbuf_4 _4218_ (.A(\egd_top.BitStream_buffer.BS_buffer[53] ),
    .X(_0703_));
 sky130_fd_sc_hd__nand2_1 _4219_ (.A(_0403_),
    .B(_0703_),
    .Y(_0704_));
 sky130_fd_sc_hd__inv_2 _4220_ (.A(\egd_top.BitStream_buffer.BS_buffer[56] ),
    .Y(_0705_));
 sky130_fd_sc_hd__or2_1 _4221_ (.A(_0705_),
    .B(_0408_),
    .X(_0706_));
 sky130_fd_sc_hd__o2111a_1 _4222_ (.A1(_0700_),
    .A2(_0397_),
    .B1(_0702_),
    .C1(_0704_),
    .D1(_0706_),
    .X(_0707_));
 sky130_fd_sc_hd__inv_2 _4223_ (.A(_0447_),
    .Y(_0708_));
 sky130_fd_sc_hd__nand2_1 _4224_ (.A(_0416_),
    .B(_0423_),
    .Y(_0709_));
 sky130_fd_sc_hd__nand2_1 _4225_ (.A(_0420_),
    .B(_0411_),
    .Y(_0710_));
 sky130_fd_sc_hd__inv_2 _4226_ (.A(_0421_),
    .Y(_0711_));
 sky130_fd_sc_hd__or2_1 _4227_ (.A(_0711_),
    .B(_0426_),
    .X(_0712_));
 sky130_fd_sc_hd__o2111a_1 _4228_ (.A1(_0708_),
    .A2(_0414_),
    .B1(_0709_),
    .C1(_0710_),
    .D1(_0712_),
    .X(_0713_));
 sky130_fd_sc_hd__inv_2 _4229_ (.A(\egd_top.BitStream_buffer.BS_buffer[49] ),
    .Y(_0714_));
 sky130_fd_sc_hd__nand2_1 _4230_ (.A(_0442_),
    .B(_0429_),
    .Y(_0715_));
 sky130_fd_sc_hd__o21ai_1 _4231_ (.A1(_0714_),
    .A2(_0440_),
    .B1(_0715_),
    .Y(_0716_));
 sky130_fd_sc_hd__a221oi_1 _4232_ (.A1(_0433_),
    .A2(_0432_),
    .B1(_0404_),
    .B2(_0436_),
    .C1(_0716_),
    .Y(_0717_));
 sky130_fd_sc_hd__nand2_1 _4233_ (.A(_0460_),
    .B(_0455_),
    .Y(_0718_));
 sky130_fd_sc_hd__o21ai_1 _4234_ (.A1(_3108_),
    .A2(_0458_),
    .B1(_0718_),
    .Y(_0719_));
 sky130_fd_sc_hd__a221oi_1 _4235_ (.A1(_0451_),
    .A2(_0450_),
    .B1(_0461_),
    .B2(_0454_),
    .C1(_0719_),
    .Y(_0720_));
 sky130_fd_sc_hd__and4_1 _4236_ (.A(_0707_),
    .B(_0713_),
    .C(_0717_),
    .D(_0720_),
    .X(_0721_));
 sky130_fd_sc_hd__and2_1 _4237_ (.A(_0699_),
    .B(_0721_),
    .X(_0722_));
 sky130_fd_sc_hd__inv_2 _4238_ (.A(_0475_),
    .Y(_0723_));
 sky130_fd_sc_hd__nand2_1 _4239_ (.A(_0474_),
    .B(_0479_),
    .Y(_0724_));
 sky130_fd_sc_hd__a22o_1 _4240_ (.A1(_0478_),
    .A2(_0482_),
    .B1(_0481_),
    .B2(_0535_),
    .X(_0725_));
 sky130_fd_sc_hd__inv_2 _4241_ (.A(_0725_),
    .Y(_0726_));
 sky130_fd_sc_hd__o211a_1 _4242_ (.A1(_0723_),
    .A2(_0472_),
    .B1(_0724_),
    .C1(_0726_),
    .X(_0727_));
 sky130_fd_sc_hd__inv_2 _4243_ (.A(_0499_),
    .Y(_0728_));
 sky130_fd_sc_hd__nand2_1 _4244_ (.A(_0498_),
    .B(_0513_),
    .Y(_0729_));
 sky130_fd_sc_hd__o21ai_1 _4245_ (.A1(_0728_),
    .A2(_0496_),
    .B1(_0729_),
    .Y(_0730_));
 sky130_fd_sc_hd__a221oi_1 _4246_ (.A1(_0489_),
    .A2(_0488_),
    .B1(_0493_),
    .B2(_0492_),
    .C1(_0730_),
    .Y(_0731_));
 sky130_fd_sc_hd__nand2_1 _4247_ (.A(_0508_),
    .B(_0503_),
    .Y(_0732_));
 sky130_fd_sc_hd__nand2_1 _4248_ (.A(_0512_),
    .B(_0515_),
    .Y(_0733_));
 sky130_fd_sc_hd__inv_2 _4249_ (.A(_0509_),
    .Y(_0734_));
 sky130_fd_sc_hd__or2_1 _4250_ (.A(_0734_),
    .B(_0518_),
    .X(_0735_));
 sky130_fd_sc_hd__o2111a_1 _4251_ (.A1(_0468_),
    .A2(_0506_),
    .B1(_0732_),
    .C1(_0733_),
    .D1(_0735_),
    .X(_0736_));
 sky130_fd_sc_hd__nand2_1 _4252_ (.A(_0530_),
    .B(_0521_),
    .Y(_0737_));
 sky130_fd_sc_hd__nand2_1 _4253_ (.A(_0534_),
    .B(_0531_),
    .Y(_0738_));
 sky130_fd_sc_hd__nand2_1 _4254_ (.A(_0737_),
    .B(_0738_),
    .Y(_0739_));
 sky130_fd_sc_hd__a221oi_1 _4255_ (.A1(_0525_),
    .A2(_0524_),
    .B1(_0359_),
    .B2(_0528_),
    .C1(_0739_),
    .Y(_0740_));
 sky130_fd_sc_hd__and4_1 _4256_ (.A(_0727_),
    .B(_0731_),
    .C(_0736_),
    .D(_0740_),
    .X(_0741_));
 sky130_fd_sc_hd__inv_2 _4257_ (.A(_0548_),
    .Y(_0742_));
 sky130_fd_sc_hd__nand2_1 _4258_ (.A(_0547_),
    .B(\egd_top.BitStream_buffer.BS_buffer[7] ),
    .Y(_0743_));
 sky130_fd_sc_hd__nand2_1 _4259_ (.A(_0551_),
    .B(_0540_),
    .Y(_0744_));
 sky130_fd_sc_hd__inv_2 _4260_ (.A(\egd_top.BitStream_buffer.BS_buffer[8] ),
    .Y(_0745_));
 sky130_fd_sc_hd__or2_1 _4261_ (.A(_0745_),
    .B(_0556_),
    .X(_0746_));
 sky130_fd_sc_hd__o2111a_1 _4262_ (.A1(_0742_),
    .A2(_0545_),
    .B1(_0743_),
    .C1(_0744_),
    .D1(_0746_),
    .X(_0747_));
 sky130_fd_sc_hd__nand2_1 _4263_ (.A(_0563_),
    .B(\egd_top.BitStream_buffer.BS_buffer[11] ),
    .Y(_0748_));
 sky130_fd_sc_hd__nand2_1 _4264_ (.A(_0566_),
    .B(\egd_top.BitStream_buffer.BS_buffer[9] ),
    .Y(_0749_));
 sky130_fd_sc_hd__inv_2 _4265_ (.A(\egd_top.BitStream_buffer.BS_buffer[10] ),
    .Y(_0750_));
 sky130_fd_sc_hd__or2_1 _4266_ (.A(_0750_),
    .B(_0570_),
    .X(_0751_));
 sky130_fd_sc_hd__o2111a_1 _4267_ (.A1(_0593_),
    .A2(_0561_),
    .B1(_0748_),
    .C1(_0749_),
    .D1(_0751_),
    .X(_0752_));
 sky130_fd_sc_hd__inv_2 _4268_ (.A(_0552_),
    .Y(_0753_));
 sky130_fd_sc_hd__or2_1 _4269_ (.A(_0753_),
    .B(_0584_),
    .X(_0754_));
 sky130_fd_sc_hd__o221a_1 _4270_ (.A1(_0582_),
    .A2(_0576_),
    .B1(_0574_),
    .B2(_0580_),
    .C1(_0754_),
    .X(_0755_));
 sky130_fd_sc_hd__inv_2 _4271_ (.A(\egd_top.BitStream_buffer.BS_buffer[14] ),
    .Y(_0756_));
 sky130_fd_sc_hd__o22ai_1 _4272_ (.A1(_0596_),
    .A2(_0595_),
    .B1(_0756_),
    .B2(_0598_),
    .Y(_0757_));
 sky130_fd_sc_hd__a221oi_1 _4273_ (.A1(\egd_top.BitStream_buffer.BS_buffer[15] ),
    .A2(_0589_),
    .B1(\egd_top.BitStream_buffer.BS_buffer[16] ),
    .B2(_0592_),
    .C1(_0757_),
    .Y(_0758_));
 sky130_fd_sc_hd__and4_1 _4274_ (.A(_0747_),
    .B(_0752_),
    .C(_0755_),
    .D(_0758_),
    .X(_0759_));
 sky130_fd_sc_hd__and3_1 _4275_ (.A(_0722_),
    .B(_0741_),
    .C(_0759_),
    .X(_0760_));
 sky130_fd_sc_hd__nand2_1 _4276_ (.A(_0606_),
    .B(_0577_),
    .Y(_0761_));
 sky130_fd_sc_hd__nand3_1 _4277_ (.A(_0680_),
    .B(_0760_),
    .C(_0761_),
    .Y(_0762_));
 sky130_fd_sc_hd__o21a_1 _4278_ (.A1(\egd_top.BitStream_buffer.BitStream_buffer_output[14] ),
    .A2(_2997_),
    .B1(_2989_),
    .X(_0763_));
 sky130_fd_sc_hd__o21a_1 _4279_ (.A1(_3056_),
    .A2(_0762_),
    .B1(_0763_),
    .X(_0296_));
 sky130_fd_sc_hd__inv_2 _4280_ (.A(_3069_),
    .Y(_0764_));
 sky130_fd_sc_hd__o22ai_1 _4281_ (.A1(_0611_),
    .A2(_3084_),
    .B1(_0764_),
    .B2(_3092_),
    .Y(_0765_));
 sky130_fd_sc_hd__a221oi_1 _4282_ (.A1(_3161_),
    .A2(_3068_),
    .B1(_3156_),
    .B2(_3075_),
    .C1(_0765_),
    .Y(_0766_));
 sky130_fd_sc_hd__inv_2 _4283_ (.A(_3095_),
    .Y(_0767_));
 sky130_fd_sc_hd__nand2_1 _4284_ (.A(_3114_),
    .B(_3102_),
    .Y(_0768_));
 sky130_fd_sc_hd__o21ai_1 _4285_ (.A1(_0767_),
    .A2(_3111_),
    .B1(_0768_),
    .Y(_0769_));
 sky130_fd_sc_hd__a221oi_1 _4286_ (.A1(_3129_),
    .A2(_3101_),
    .B1(_3136_),
    .B2(_3106_),
    .C1(_0769_),
    .Y(_0770_));
 sky130_fd_sc_hd__nand2_1 _4287_ (.A(_3128_),
    .B(_3134_),
    .Y(_0771_));
 sky130_fd_sc_hd__nand2_1 _4288_ (.A(_3133_),
    .B(_3076_),
    .Y(_0772_));
 sky130_fd_sc_hd__or2_1 _4289_ (.A(_3120_),
    .B(_3141_),
    .X(_0773_));
 sky130_fd_sc_hd__o2111a_1 _4290_ (.A1(_3086_),
    .A2(_3124_),
    .B1(_0771_),
    .C1(_0772_),
    .D1(_0773_),
    .X(_0774_));
 sky130_fd_sc_hd__nand2_1 _4291_ (.A(_3155_),
    .B(_3149_),
    .Y(_0775_));
 sky130_fd_sc_hd__nand2_1 _4292_ (.A(_3160_),
    .B(_3144_),
    .Y(_0776_));
 sky130_fd_sc_hd__nand2_1 _4293_ (.A(_0775_),
    .B(_0776_),
    .Y(_0777_));
 sky130_fd_sc_hd__a221oi_1 _4294_ (.A1(_3255_),
    .A2(_3148_),
    .B1(_3247_),
    .B2(_3152_),
    .C1(_0777_),
    .Y(_0778_));
 sky130_fd_sc_hd__and4_1 _4295_ (.A(_0766_),
    .B(_0770_),
    .C(_0774_),
    .D(_0778_),
    .X(_0779_));
 sky130_fd_sc_hd__inv_2 _4296_ (.A(\egd_top.BitStream_buffer.BS_buffer[119] ),
    .Y(_0780_));
 sky130_fd_sc_hd__o22ai_1 _4297_ (.A1(_0628_),
    .A2(_3176_),
    .B1(_0780_),
    .B2(_3179_),
    .Y(_0781_));
 sky130_fd_sc_hd__a221oi_1 _4298_ (.A1(_3031_),
    .A2(_3170_),
    .B1(_3034_),
    .B2(_3173_),
    .C1(_0781_),
    .Y(_0782_));
 sky130_fd_sc_hd__nand2_1 _4299_ (.A(_3192_),
    .B(_3044_),
    .Y(_0783_));
 sky130_fd_sc_hd__o21ai_1 _4300_ (.A1(_3219_),
    .A2(_3190_),
    .B1(_0783_),
    .Y(_0784_));
 sky130_fd_sc_hd__a221oi_1 _4301_ (.A1(_3037_),
    .A2(_3184_),
    .B1(_3040_),
    .B2(_3187_),
    .C1(_0784_),
    .Y(_0785_));
 sky130_fd_sc_hd__inv_2 _4302_ (.A(\egd_top.BitStream_buffer.BS_buffer[114] ),
    .Y(_0786_));
 sky130_fd_sc_hd__nand2_1 _4303_ (.A(_3206_),
    .B(_3016_),
    .Y(_0787_));
 sky130_fd_sc_hd__o21ai_1 _4304_ (.A1(_0786_),
    .A2(_3204_),
    .B1(_0787_),
    .Y(_0788_));
 sky130_fd_sc_hd__a221oi_1 _4305_ (.A1(_3019_),
    .A2(_3198_),
    .B1(_3022_),
    .B2(_3201_),
    .C1(_0788_),
    .Y(_0789_));
 sky130_fd_sc_hd__inv_2 _4306_ (.A(_3053_),
    .Y(_0790_));
 sky130_fd_sc_hd__o22ai_1 _4307_ (.A1(_0638_),
    .A2(_3218_),
    .B1(_0790_),
    .B2(_3221_),
    .Y(_0791_));
 sky130_fd_sc_hd__a221oi_1 _4308_ (.A1(_0607_),
    .A2(_3212_),
    .B1(_0577_),
    .B2(_3215_),
    .C1(_0791_),
    .Y(_0792_));
 sky130_fd_sc_hd__and4_1 _4309_ (.A(_0782_),
    .B(_0785_),
    .C(_0789_),
    .D(_0792_),
    .X(_0793_));
 sky130_fd_sc_hd__inv_2 _4310_ (.A(\egd_top.BitStream_buffer.BS_buffer[91] ),
    .Y(_0794_));
 sky130_fd_sc_hd__o22ai_1 _4311_ (.A1(_0642_),
    .A2(_3238_),
    .B1(_0794_),
    .B2(_3241_),
    .Y(_0795_));
 sky130_fd_sc_hd__a221oi_1 _4312_ (.A1(_3286_),
    .A2(_3231_),
    .B1(_3290_),
    .B2(_3235_),
    .C1(_0795_),
    .Y(_0796_));
 sky130_fd_sc_hd__nand2_1 _4313_ (.A(_3246_),
    .B(_3251_),
    .Y(_0797_));
 sky130_fd_sc_hd__nand2_1 _4314_ (.A(_3250_),
    .B(_3265_),
    .Y(_0798_));
 sky130_fd_sc_hd__nand2_1 _4315_ (.A(_3254_),
    .B(_3259_),
    .Y(_0799_));
 sky130_fd_sc_hd__nand2_1 _4316_ (.A(_3258_),
    .B(_0646_),
    .Y(_0800_));
 sky130_fd_sc_hd__and4_1 _4317_ (.A(_0797_),
    .B(_0798_),
    .C(_0799_),
    .D(_0800_),
    .X(_0801_));
 sky130_fd_sc_hd__inv_2 _4318_ (.A(\egd_top.BitStream_buffer.BS_buffer[87] ),
    .Y(_0802_));
 sky130_fd_sc_hd__o22ai_1 _4319_ (.A1(_0651_),
    .A2(_3264_),
    .B1(_0802_),
    .B2(_3268_),
    .Y(_0803_));
 sky130_fd_sc_hd__buf_4 _4320_ (.A(\egd_top.BitStream_buffer.BS_buffer[89] ),
    .X(_0804_));
 sky130_fd_sc_hd__a22o_1 _4321_ (.A1(_3271_),
    .A2(_0653_),
    .B1(_3274_),
    .B2(_0804_),
    .X(_0805_));
 sky130_fd_sc_hd__nor2_1 _4322_ (.A(_0803_),
    .B(_0805_),
    .Y(_0806_));
 sky130_fd_sc_hd__inv_2 _4323_ (.A(_3282_),
    .Y(_0807_));
 sky130_fd_sc_hd__o22ai_1 _4324_ (.A1(_0656_),
    .A2(_3289_),
    .B1(_0807_),
    .B2(_3293_),
    .Y(_0808_));
 sky130_fd_sc_hd__a221oi_1 _4325_ (.A1(_3318_),
    .A2(_3281_),
    .B1(_3322_),
    .B2(_3285_),
    .C1(_0808_),
    .Y(_0809_));
 sky130_fd_sc_hd__and4_1 _4326_ (.A(_0796_),
    .B(_0801_),
    .C(_0806_),
    .D(_0809_),
    .X(_0810_));
 sky130_fd_sc_hd__nand2_1 _4327_ (.A(_3309_),
    .B(_3304_),
    .Y(_0811_));
 sky130_fd_sc_hd__nand2_1 _4328_ (.A(_3313_),
    .B(_3297_),
    .Y(_0812_));
 sky130_fd_sc_hd__nand2_1 _4329_ (.A(_0811_),
    .B(_0812_),
    .Y(_0813_));
 sky130_fd_sc_hd__a221oi_1 _4330_ (.A1(_3353_),
    .A2(_3303_),
    .B1(_3357_),
    .B2(_3307_),
    .C1(_0813_),
    .Y(_0814_));
 sky130_fd_sc_hd__nand2_1 _4331_ (.A(_3326_),
    .B(_3347_),
    .Y(_0815_));
 sky130_fd_sc_hd__nand2_1 _4332_ (.A(_3330_),
    .B(_3341_),
    .Y(_0816_));
 sky130_fd_sc_hd__nand2_1 _4333_ (.A(_0815_),
    .B(_0816_),
    .Y(_0817_));
 sky130_fd_sc_hd__a221oi_1 _4334_ (.A1(_3331_),
    .A2(_3321_),
    .B1(_3327_),
    .B2(_3324_),
    .C1(_0817_),
    .Y(_0818_));
 sky130_fd_sc_hd__inv_2 _4335_ (.A(\egd_top.BitStream_buffer.BS_buffer[105] ),
    .Y(_0819_));
 sky130_fd_sc_hd__nand2_1 _4336_ (.A(_3340_),
    .B(_3345_),
    .Y(_0820_));
 sky130_fd_sc_hd__nand2_1 _4337_ (.A(_3344_),
    .B(_3314_),
    .Y(_0821_));
 sky130_fd_sc_hd__or2_1 _4338_ (.A(_3336_),
    .B(_3350_),
    .X(_0822_));
 sky130_fd_sc_hd__o2111a_1 _4339_ (.A1(_0819_),
    .A2(_3338_),
    .B1(_0820_),
    .C1(_0821_),
    .D1(_0822_),
    .X(_0823_));
 sky130_fd_sc_hd__nand2_1 _4340_ (.A(_3365_),
    .B(_2998_),
    .Y(_0824_));
 sky130_fd_sc_hd__o21ai_1 _4341_ (.A1(_0634_),
    .A2(_3363_),
    .B1(_0824_),
    .Y(_0825_));
 sky130_fd_sc_hd__a221oi_1 _4342_ (.A1(_0674_),
    .A2(_3356_),
    .B1(_0675_),
    .B2(_3360_),
    .C1(_0825_),
    .Y(_0826_));
 sky130_fd_sc_hd__and4_1 _4343_ (.A(_0814_),
    .B(_0818_),
    .C(_0823_),
    .D(_0826_),
    .X(_0827_));
 sky130_fd_sc_hd__and4_1 _4344_ (.A(_0779_),
    .B(_0793_),
    .C(_0810_),
    .D(_0827_),
    .X(_0828_));
 sky130_fd_sc_hd__nand2_1 _4345_ (.A(_0334_),
    .B(_0329_),
    .Y(_0829_));
 sky130_fd_sc_hd__nand2_1 _4346_ (.A(_0338_),
    .B(_0323_),
    .Y(_0830_));
 sky130_fd_sc_hd__nand2_1 _4347_ (.A(_0829_),
    .B(_0830_),
    .Y(_0831_));
 sky130_fd_sc_hd__a221oi_1 _4348_ (.A1(_0376_),
    .A2(_0328_),
    .B1(_0380_),
    .B2(_0332_),
    .C1(_0831_),
    .Y(_0832_));
 sky130_fd_sc_hd__inv_2 _4349_ (.A(\egd_top.BitStream_buffer.BS_buffer[39] ),
    .Y(_0833_));
 sky130_fd_sc_hd__o22ai_1 _4350_ (.A1(_0685_),
    .A2(_0345_),
    .B1(_0833_),
    .B2(_0349_),
    .Y(_0834_));
 sky130_fd_sc_hd__a22o_1 _4351_ (.A1(_0352_),
    .A2(_0339_),
    .B1(_0355_),
    .B2(_0335_),
    .X(_0835_));
 sky130_fd_sc_hd__nor2_1 _4352_ (.A(_0834_),
    .B(_0835_),
    .Y(_0836_));
 sky130_fd_sc_hd__nand2_1 _4353_ (.A(_0371_),
    .B(_0346_),
    .Y(_0837_));
 sky130_fd_sc_hd__o21ai_1 _4354_ (.A1(_0343_),
    .A2(_0369_),
    .B1(_0837_),
    .Y(_0838_));
 sky130_fd_sc_hd__a221oi_1 _4355_ (.A1(_0689_),
    .A2(_0362_),
    .B1(_0372_),
    .B2(_0366_),
    .C1(_0838_),
    .Y(_0839_));
 sky130_fd_sc_hd__nand2_1 _4356_ (.A(_0388_),
    .B(_0437_),
    .Y(_0840_));
 sky130_fd_sc_hd__o21ai_1 _4357_ (.A1(_0714_),
    .A2(_0386_),
    .B1(_0840_),
    .Y(_0841_));
 sky130_fd_sc_hd__a221oi_1 _4358_ (.A1(_0389_),
    .A2(_0379_),
    .B1(_0695_),
    .B2(_0383_),
    .C1(_0841_),
    .Y(_0842_));
 sky130_fd_sc_hd__and4_1 _4359_ (.A(_0832_),
    .B(_0836_),
    .C(_0839_),
    .D(_0842_),
    .X(_0843_));
 sky130_fd_sc_hd__nand2_1 _4360_ (.A(_0399_),
    .B(_0417_),
    .Y(_0844_));
 sky130_fd_sc_hd__nand2_1 _4361_ (.A(_0403_),
    .B(_0400_),
    .Y(_0845_));
 sky130_fd_sc_hd__or2_1 _4362_ (.A(_0424_),
    .B(_0408_),
    .X(_0846_));
 sky130_fd_sc_hd__o2111a_1 _4363_ (.A1(_0406_),
    .A2(_0397_),
    .B1(_0844_),
    .C1(_0845_),
    .D1(_0846_),
    .X(_0847_));
 sky130_fd_sc_hd__inv_2 _4364_ (.A(_0451_),
    .Y(_0848_));
 sky130_fd_sc_hd__nand2_1 _4365_ (.A(_0416_),
    .B(_0421_),
    .Y(_0849_));
 sky130_fd_sc_hd__nand2_1 _4366_ (.A(_0420_),
    .B(_0447_),
    .Y(_0850_));
 sky130_fd_sc_hd__or2_1 _4367_ (.A(_0412_),
    .B(_0426_),
    .X(_0851_));
 sky130_fd_sc_hd__o2111a_1 _4368_ (.A1(_0848_),
    .A2(_0414_),
    .B1(_0849_),
    .C1(_0850_),
    .D1(_0851_),
    .X(_0852_));
 sky130_fd_sc_hd__inv_2 _4369_ (.A(\egd_top.BitStream_buffer.BS_buffer[50] ),
    .Y(_0853_));
 sky130_fd_sc_hd__nand2_1 _4370_ (.A(_0442_),
    .B(_0433_),
    .Y(_0854_));
 sky130_fd_sc_hd__o21ai_1 _4371_ (.A1(_0853_),
    .A2(_0440_),
    .B1(_0854_),
    .Y(_0855_));
 sky130_fd_sc_hd__a221oi_1 _4372_ (.A1(_0404_),
    .A2(_0432_),
    .B1(_0703_),
    .B2(_0436_),
    .C1(_0855_),
    .Y(_0856_));
 sky130_fd_sc_hd__nand2_1 _4373_ (.A(_0460_),
    .B(_3107_),
    .Y(_0857_));
 sky130_fd_sc_hd__o21ai_1 _4374_ (.A1(_0614_),
    .A2(_0458_),
    .B1(_0857_),
    .Y(_0858_));
 sky130_fd_sc_hd__a221oi_1 _4375_ (.A1(_0461_),
    .A2(_0450_),
    .B1(_0455_),
    .B2(_0454_),
    .C1(_0858_),
    .Y(_0859_));
 sky130_fd_sc_hd__and4_1 _4376_ (.A(_0847_),
    .B(_0852_),
    .C(_0856_),
    .D(_0859_),
    .X(_0860_));
 sky130_fd_sc_hd__and2_1 _4377_ (.A(_0843_),
    .B(_0860_),
    .X(_0861_));
 sky130_fd_sc_hd__inv_2 _4378_ (.A(_0479_),
    .Y(_0862_));
 sky130_fd_sc_hd__nand2_1 _4379_ (.A(_0474_),
    .B(_0482_),
    .Y(_0863_));
 sky130_fd_sc_hd__a22o_1 _4380_ (.A1(_0478_),
    .A2(_0535_),
    .B1(_0481_),
    .B2(_0531_),
    .X(_0864_));
 sky130_fd_sc_hd__inv_2 _4381_ (.A(_0864_),
    .Y(_0865_));
 sky130_fd_sc_hd__o211a_1 _4382_ (.A1(_0862_),
    .A2(_0472_),
    .B1(_0863_),
    .C1(_0865_),
    .X(_0866_));
 sky130_fd_sc_hd__inv_2 _4383_ (.A(_0513_),
    .Y(_0867_));
 sky130_fd_sc_hd__nand2_1 _4384_ (.A(_0498_),
    .B(_0515_),
    .Y(_0868_));
 sky130_fd_sc_hd__o21ai_1 _4385_ (.A1(_0867_),
    .A2(_0496_),
    .B1(_0868_),
    .Y(_0869_));
 sky130_fd_sc_hd__a221oi_1 _4386_ (.A1(_0493_),
    .A2(_0488_),
    .B1(_0499_),
    .B2(_0492_),
    .C1(_0869_),
    .Y(_0870_));
 sky130_fd_sc_hd__nand2_1 _4387_ (.A(_0508_),
    .B(_0467_),
    .Y(_0871_));
 sky130_fd_sc_hd__nand2_1 _4388_ (.A(_0512_),
    .B(_0509_),
    .Y(_0872_));
 sky130_fd_sc_hd__or2_1 _4389_ (.A(_0504_),
    .B(_0518_),
    .X(_0873_));
 sky130_fd_sc_hd__o2111a_1 _4390_ (.A1(_0723_),
    .A2(_0506_),
    .B1(_0871_),
    .C1(_0872_),
    .D1(_0873_),
    .X(_0874_));
 sky130_fd_sc_hd__nand2_1 _4391_ (.A(_0530_),
    .B(_0525_),
    .Y(_0875_));
 sky130_fd_sc_hd__nand2_1 _4392_ (.A(_0534_),
    .B(_0521_),
    .Y(_0876_));
 sky130_fd_sc_hd__nand2_1 _4393_ (.A(_0875_),
    .B(_0876_),
    .Y(_0877_));
 sky130_fd_sc_hd__a221oi_1 _4394_ (.A1(_0359_),
    .A2(_0524_),
    .B1(_0363_),
    .B2(_0528_),
    .C1(_0877_),
    .Y(_0878_));
 sky130_fd_sc_hd__and4_1 _4395_ (.A(_0866_),
    .B(_0870_),
    .C(_0874_),
    .D(_0878_),
    .X(_0879_));
 sky130_fd_sc_hd__nand2_1 _4396_ (.A(_0547_),
    .B(\egd_top.BitStream_buffer.BS_buffer[8] ),
    .Y(_0880_));
 sky130_fd_sc_hd__nand2_1 _4397_ (.A(_0551_),
    .B(_0548_),
    .Y(_0881_));
 sky130_fd_sc_hd__or2_1 _4398_ (.A(_0568_),
    .B(_0556_),
    .X(_0882_));
 sky130_fd_sc_hd__o2111a_1 _4399_ (.A1(_0554_),
    .A2(_0545_),
    .B1(_0880_),
    .C1(_0881_),
    .D1(_0882_),
    .X(_0883_));
 sky130_fd_sc_hd__nand2_1 _4400_ (.A(_0563_),
    .B(\egd_top.BitStream_buffer.BS_buffer[12] ),
    .Y(_0884_));
 sky130_fd_sc_hd__nand2_1 _4401_ (.A(_0566_),
    .B(\egd_top.BitStream_buffer.BS_buffer[10] ),
    .Y(_0885_));
 sky130_fd_sc_hd__or2_1 _4402_ (.A(_0559_),
    .B(_0570_),
    .X(_0886_));
 sky130_fd_sc_hd__o2111a_1 _4403_ (.A1(_0596_),
    .A2(_0561_),
    .B1(_0884_),
    .C1(_0885_),
    .D1(_0886_),
    .X(_0887_));
 sky130_fd_sc_hd__or2_1 _4404_ (.A(_0541_),
    .B(_0584_),
    .X(_0888_));
 sky130_fd_sc_hd__o221a_1 _4405_ (.A1(_0753_),
    .A2(_0576_),
    .B1(_0582_),
    .B2(_0580_),
    .C1(_0888_),
    .X(_0889_));
 sky130_fd_sc_hd__inv_2 _4406_ (.A(\egd_top.BitStream_buffer.BS_buffer[15] ),
    .Y(_0890_));
 sky130_fd_sc_hd__o22ai_1 _4407_ (.A1(_0756_),
    .A2(_0595_),
    .B1(_0890_),
    .B2(_0598_),
    .Y(_0891_));
 sky130_fd_sc_hd__a221oi_1 _4408_ (.A1(\egd_top.BitStream_buffer.BS_buffer[16] ),
    .A2(_0589_),
    .B1(_0489_),
    .B2(_0592_),
    .C1(_0891_),
    .Y(_0892_));
 sky130_fd_sc_hd__and4_1 _4409_ (.A(_0883_),
    .B(_0887_),
    .C(_0889_),
    .D(_0892_),
    .X(_0893_));
 sky130_fd_sc_hd__and3_1 _4410_ (.A(_0861_),
    .B(_0879_),
    .C(_0893_),
    .X(_0894_));
 sky130_fd_sc_hd__nand2_1 _4411_ (.A(_0606_),
    .B(_0573_),
    .Y(_0895_));
 sky130_fd_sc_hd__nand3_1 _4412_ (.A(_0828_),
    .B(_0894_),
    .C(_0895_),
    .Y(_0896_));
 sky130_fd_sc_hd__inv_2 _4413_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[13] ),
    .Y(_0897_));
 sky130_fd_sc_hd__clkbuf_4 _4414_ (.A(_2996_),
    .X(_0898_));
 sky130_fd_sc_hd__a21oi_1 _4415_ (.A1(_0897_),
    .A2(_0898_),
    .B1(_2938_),
    .Y(_0899_));
 sky130_fd_sc_hd__o21a_1 _4416_ (.A1(_3056_),
    .A2(_0896_),
    .B1(_0899_),
    .X(_0295_));
 sky130_fd_sc_hd__inv_2 _4417_ (.A(_3161_),
    .Y(_0900_));
 sky130_fd_sc_hd__o22ai_1 _4418_ (.A1(_0764_),
    .A2(_3084_),
    .B1(_0900_),
    .B2(_3092_),
    .Y(_0901_));
 sky130_fd_sc_hd__a221oi_1 _4419_ (.A1(_3156_),
    .A2(_3068_),
    .B1(_3144_),
    .B2(_3075_),
    .C1(_0901_),
    .Y(_0902_));
 sky130_fd_sc_hd__inv_2 _4420_ (.A(_3102_),
    .Y(_0903_));
 sky130_fd_sc_hd__nand2_1 _4421_ (.A(_3114_),
    .B(_3129_),
    .Y(_0904_));
 sky130_fd_sc_hd__o21ai_1 _4422_ (.A1(_0903_),
    .A2(_3111_),
    .B1(_0904_),
    .Y(_0905_));
 sky130_fd_sc_hd__a221oi_1 _4423_ (.A1(_3136_),
    .A2(_3101_),
    .B1(_3134_),
    .B2(_3106_),
    .C1(_0905_),
    .Y(_0906_));
 sky130_fd_sc_hd__nand2_1 _4424_ (.A(_3128_),
    .B(_3119_),
    .Y(_0907_));
 sky130_fd_sc_hd__nand2_1 _4425_ (.A(_3133_),
    .B(_3085_),
    .Y(_0908_));
 sky130_fd_sc_hd__or2_1 _4426_ (.A(_3077_),
    .B(_3141_),
    .X(_0909_));
 sky130_fd_sc_hd__o2111a_1 _4427_ (.A1(_0611_),
    .A2(_3124_),
    .B1(_0907_),
    .C1(_0908_),
    .D1(_0909_),
    .X(_0910_));
 sky130_fd_sc_hd__nand2_1 _4428_ (.A(_3155_),
    .B(_3255_),
    .Y(_0911_));
 sky130_fd_sc_hd__nand2_1 _4429_ (.A(_3160_),
    .B(_3149_),
    .Y(_0912_));
 sky130_fd_sc_hd__nand2_1 _4430_ (.A(_0911_),
    .B(_0912_),
    .Y(_0913_));
 sky130_fd_sc_hd__a221oi_1 _4431_ (.A1(_3247_),
    .A2(_3148_),
    .B1(_3259_),
    .B2(_3152_),
    .C1(_0913_),
    .Y(_0914_));
 sky130_fd_sc_hd__and4_1 _4432_ (.A(_0902_),
    .B(_0906_),
    .C(_0910_),
    .D(_0914_),
    .X(_0915_));
 sky130_fd_sc_hd__inv_2 _4433_ (.A(\egd_top.BitStream_buffer.BS_buffer[120] ),
    .Y(_0916_));
 sky130_fd_sc_hd__o22ai_1 _4434_ (.A1(_0780_),
    .A2(_3176_),
    .B1(_0916_),
    .B2(_3179_),
    .Y(_0917_));
 sky130_fd_sc_hd__a221oi_1 _4435_ (.A1(_3034_),
    .A2(_3170_),
    .B1(_3037_),
    .B2(_3173_),
    .C1(_0917_),
    .Y(_0918_));
 sky130_fd_sc_hd__nand2_1 _4436_ (.A(_3192_),
    .B(_3047_),
    .Y(_0919_));
 sky130_fd_sc_hd__o21ai_1 _4437_ (.A1(_0638_),
    .A2(_3190_),
    .B1(_0919_),
    .Y(_0920_));
 sky130_fd_sc_hd__a221oi_1 _4438_ (.A1(_3040_),
    .A2(_3184_),
    .B1(_3044_),
    .B2(_3187_),
    .C1(_0920_),
    .Y(_0921_));
 sky130_fd_sc_hd__inv_2 _4439_ (.A(\egd_top.BitStream_buffer.BS_buffer[115] ),
    .Y(_0922_));
 sky130_fd_sc_hd__nand2_1 _4440_ (.A(_3206_),
    .B(_3019_),
    .Y(_0923_));
 sky130_fd_sc_hd__o21ai_1 _4441_ (.A1(_0922_),
    .A2(_3204_),
    .B1(_0923_),
    .Y(_0924_));
 sky130_fd_sc_hd__a221oi_1 _4442_ (.A1(_3022_),
    .A2(_3198_),
    .B1(_3025_),
    .B2(_3201_),
    .C1(_0924_),
    .Y(_0925_));
 sky130_fd_sc_hd__inv_2 _4443_ (.A(_0607_),
    .Y(_0926_));
 sky130_fd_sc_hd__o22ai_1 _4444_ (.A1(_0790_),
    .A2(_3218_),
    .B1(_0926_),
    .B2(_3221_),
    .Y(_0927_));
 sky130_fd_sc_hd__a221oi_1 _4445_ (.A1(_0577_),
    .A2(_3212_),
    .B1(_0573_),
    .B2(_3215_),
    .C1(_0927_),
    .Y(_0928_));
 sky130_fd_sc_hd__and4_1 _4446_ (.A(_0918_),
    .B(_0921_),
    .C(_0925_),
    .D(_0928_),
    .X(_0929_));
 sky130_fd_sc_hd__o22ai_1 _4447_ (.A1(_0794_),
    .A2(_3238_),
    .B1(_3287_),
    .B2(_3241_),
    .Y(_0930_));
 sky130_fd_sc_hd__a221oi_1 _4448_ (.A1(_3290_),
    .A2(_3231_),
    .B1(_3278_),
    .B2(_3235_),
    .C1(_0930_),
    .Y(_0931_));
 sky130_fd_sc_hd__nand2_1 _4449_ (.A(_3246_),
    .B(_0646_),
    .Y(_0932_));
 sky130_fd_sc_hd__nand2_1 _4450_ (.A(_3250_),
    .B(_3272_),
    .Y(_0933_));
 sky130_fd_sc_hd__nand2_1 _4451_ (.A(_3254_),
    .B(_3251_),
    .Y(_0934_));
 sky130_fd_sc_hd__nand2_1 _4452_ (.A(_3258_),
    .B(_3265_),
    .Y(_0935_));
 sky130_fd_sc_hd__and4_1 _4453_ (.A(_0932_),
    .B(_0933_),
    .C(_0934_),
    .D(_0935_),
    .X(_0936_));
 sky130_fd_sc_hd__o22ai_1 _4454_ (.A1(_0802_),
    .A2(_3264_),
    .B1(_3236_),
    .B2(_3268_),
    .Y(_0937_));
 sky130_fd_sc_hd__a22o_1 _4455_ (.A1(_3271_),
    .A2(_0804_),
    .B1(_3274_),
    .B2(_3225_),
    .X(_0938_));
 sky130_fd_sc_hd__nor2_1 _4456_ (.A(_0937_),
    .B(_0938_),
    .Y(_0939_));
 sky130_fd_sc_hd__inv_2 _4457_ (.A(_3318_),
    .Y(_0940_));
 sky130_fd_sc_hd__o22ai_1 _4458_ (.A1(_0807_),
    .A2(_3289_),
    .B1(_0940_),
    .B2(_3293_),
    .Y(_0941_));
 sky130_fd_sc_hd__a221oi_1 _4459_ (.A1(_3322_),
    .A2(_3281_),
    .B1(_3331_),
    .B2(_3285_),
    .C1(_0941_),
    .Y(_0942_));
 sky130_fd_sc_hd__and4_1 _4460_ (.A(_0931_),
    .B(_0936_),
    .C(_0939_),
    .D(_0942_),
    .X(_0943_));
 sky130_fd_sc_hd__nand2_1 _4461_ (.A(_3309_),
    .B(_3353_),
    .Y(_0944_));
 sky130_fd_sc_hd__nand2_1 _4462_ (.A(_3313_),
    .B(_3304_),
    .Y(_0945_));
 sky130_fd_sc_hd__nand2_1 _4463_ (.A(_0944_),
    .B(_0945_),
    .Y(_0946_));
 sky130_fd_sc_hd__a221oi_1 _4464_ (.A1(_3357_),
    .A2(_3303_),
    .B1(_0674_),
    .B2(_3307_),
    .C1(_0946_),
    .Y(_0947_));
 sky130_fd_sc_hd__nand2_1 _4465_ (.A(_3326_),
    .B(_3345_),
    .Y(_0948_));
 sky130_fd_sc_hd__nand2_1 _4466_ (.A(_3330_),
    .B(_3347_),
    .Y(_0949_));
 sky130_fd_sc_hd__nand2_1 _4467_ (.A(_0948_),
    .B(_0949_),
    .Y(_0950_));
 sky130_fd_sc_hd__a221oi_1 _4468_ (.A1(_3327_),
    .A2(_3321_),
    .B1(_3341_),
    .B2(_3324_),
    .C1(_0950_),
    .Y(_0951_));
 sky130_fd_sc_hd__inv_2 _4469_ (.A(\egd_top.BitStream_buffer.BS_buffer[106] ),
    .Y(_0952_));
 sky130_fd_sc_hd__nand2_1 _4470_ (.A(_3340_),
    .B(_3335_),
    .Y(_0953_));
 sky130_fd_sc_hd__nand2_1 _4471_ (.A(_3344_),
    .B(_3310_),
    .Y(_0954_));
 sky130_fd_sc_hd__or2_1 _4472_ (.A(_0668_),
    .B(_3350_),
    .X(_0955_));
 sky130_fd_sc_hd__o2111a_1 _4473_ (.A1(_0952_),
    .A2(_3338_),
    .B1(_0953_),
    .C1(_0954_),
    .D1(_0955_),
    .X(_0956_));
 sky130_fd_sc_hd__nand2_1 _4474_ (.A(_3365_),
    .B(_3010_),
    .Y(_0957_));
 sky130_fd_sc_hd__o21ai_1 _4475_ (.A1(_0786_),
    .A2(_3363_),
    .B1(_0957_),
    .Y(_0958_));
 sky130_fd_sc_hd__a221oi_1 _4476_ (.A1(_0675_),
    .A2(_3356_),
    .B1(_2998_),
    .B2(_3360_),
    .C1(_0958_),
    .Y(_0959_));
 sky130_fd_sc_hd__and4_1 _4477_ (.A(_0947_),
    .B(_0951_),
    .C(_0956_),
    .D(_0959_),
    .X(_0960_));
 sky130_fd_sc_hd__and4_1 _4478_ (.A(_0915_),
    .B(_0929_),
    .C(_0943_),
    .D(_0960_),
    .X(_0961_));
 sky130_fd_sc_hd__nand2_1 _4479_ (.A(_0334_),
    .B(_0376_),
    .Y(_0962_));
 sky130_fd_sc_hd__nand2_1 _4480_ (.A(_0338_),
    .B(_0329_),
    .Y(_0963_));
 sky130_fd_sc_hd__nand2_1 _4481_ (.A(_0962_),
    .B(_0963_),
    .Y(_0964_));
 sky130_fd_sc_hd__a221oi_1 _4482_ (.A1(_0380_),
    .A2(_0328_),
    .B1(_0389_),
    .B2(_0332_),
    .C1(_0964_),
    .Y(_0965_));
 sky130_fd_sc_hd__inv_2 _4483_ (.A(\egd_top.BitStream_buffer.BS_buffer[40] ),
    .Y(_0966_));
 sky130_fd_sc_hd__o22ai_1 _4484_ (.A1(_0833_),
    .A2(_0345_),
    .B1(_0966_),
    .B2(_0349_),
    .Y(_0967_));
 sky130_fd_sc_hd__a22o_1 _4485_ (.A1(_0352_),
    .A2(_0335_),
    .B1(_0355_),
    .B2(_0323_),
    .X(_0968_));
 sky130_fd_sc_hd__nor2_1 _4486_ (.A(_0967_),
    .B(_0968_),
    .Y(_0969_));
 sky130_fd_sc_hd__nand2_1 _4487_ (.A(_0371_),
    .B(_0353_),
    .Y(_0970_));
 sky130_fd_sc_hd__o21ai_1 _4488_ (.A1(_0347_),
    .A2(_0369_),
    .B1(_0970_),
    .Y(_0971_));
 sky130_fd_sc_hd__a221oi_1 _4489_ (.A1(_0372_),
    .A2(_0362_),
    .B1(_0691_),
    .B2(_0366_),
    .C1(_0971_),
    .Y(_0972_));
 sky130_fd_sc_hd__nand2_1 _4490_ (.A(_0388_),
    .B(_0443_),
    .Y(_0973_));
 sky130_fd_sc_hd__o21ai_1 _4491_ (.A1(_0853_),
    .A2(_0386_),
    .B1(_0973_),
    .Y(_0974_));
 sky130_fd_sc_hd__a221oi_1 _4492_ (.A1(_0695_),
    .A2(_0379_),
    .B1(_0437_),
    .B2(_0383_),
    .C1(_0974_),
    .Y(_0975_));
 sky130_fd_sc_hd__and4_1 _4493_ (.A(_0965_),
    .B(_0969_),
    .C(_0972_),
    .D(_0975_),
    .X(_0976_));
 sky130_fd_sc_hd__nand2_1 _4494_ (.A(_0399_),
    .B(_0423_),
    .Y(_0977_));
 sky130_fd_sc_hd__nand2_1 _4495_ (.A(_0403_),
    .B(_0701_),
    .Y(_0978_));
 sky130_fd_sc_hd__or2_1 _4496_ (.A(_0711_),
    .B(_0408_),
    .X(_0979_));
 sky130_fd_sc_hd__o2111a_1 _4497_ (.A1(_0705_),
    .A2(_0397_),
    .B1(_0977_),
    .C1(_0978_),
    .D1(_0979_),
    .X(_0980_));
 sky130_fd_sc_hd__inv_2 _4498_ (.A(_0461_),
    .Y(_0981_));
 sky130_fd_sc_hd__nand2_1 _4499_ (.A(_0416_),
    .B(_0411_),
    .Y(_0982_));
 sky130_fd_sc_hd__nand2_1 _4500_ (.A(_0420_),
    .B(_0451_),
    .Y(_0983_));
 sky130_fd_sc_hd__or2_1 _4501_ (.A(_0708_),
    .B(_0426_),
    .X(_0984_));
 sky130_fd_sc_hd__o2111a_1 _4502_ (.A1(_0981_),
    .A2(_0414_),
    .B1(_0982_),
    .C1(_0983_),
    .D1(_0984_),
    .X(_0985_));
 sky130_fd_sc_hd__inv_2 _4503_ (.A(\egd_top.BitStream_buffer.BS_buffer[51] ),
    .Y(_0986_));
 sky130_fd_sc_hd__nand2_1 _4504_ (.A(_0442_),
    .B(_0404_),
    .Y(_0987_));
 sky130_fd_sc_hd__o21ai_1 _4505_ (.A1(_0986_),
    .A2(_0440_),
    .B1(_0987_),
    .Y(_0988_));
 sky130_fd_sc_hd__a221oi_1 _4506_ (.A1(_0703_),
    .A2(_0432_),
    .B1(_0400_),
    .B2(_0436_),
    .C1(_0988_),
    .Y(_0989_));
 sky130_fd_sc_hd__nand2_1 _4507_ (.A(_0460_),
    .B(_3115_),
    .Y(_0990_));
 sky130_fd_sc_hd__o21ai_1 _4508_ (.A1(_0767_),
    .A2(_0458_),
    .B1(_0990_),
    .Y(_0991_));
 sky130_fd_sc_hd__a221oi_1 _4509_ (.A1(_0455_),
    .A2(_0450_),
    .B1(_3107_),
    .B2(_0454_),
    .C1(_0991_),
    .Y(_0992_));
 sky130_fd_sc_hd__and4_1 _4510_ (.A(_0980_),
    .B(_0985_),
    .C(_0989_),
    .D(_0992_),
    .X(_0993_));
 sky130_fd_sc_hd__and2_1 _4511_ (.A(_0976_),
    .B(_0993_),
    .X(_0994_));
 sky130_fd_sc_hd__inv_2 _4512_ (.A(_0482_),
    .Y(_0995_));
 sky130_fd_sc_hd__nand2_1 _4513_ (.A(_0474_),
    .B(_0535_),
    .Y(_0996_));
 sky130_fd_sc_hd__a22o_1 _4514_ (.A1(_0478_),
    .A2(_0531_),
    .B1(_0481_),
    .B2(_0521_),
    .X(_0997_));
 sky130_fd_sc_hd__inv_2 _4515_ (.A(_0997_),
    .Y(_0998_));
 sky130_fd_sc_hd__o211a_1 _4516_ (.A1(_0995_),
    .A2(_0472_),
    .B1(_0996_),
    .C1(_0998_),
    .X(_0999_));
 sky130_fd_sc_hd__nand2_1 _4517_ (.A(_0498_),
    .B(_0509_),
    .Y(_1000_));
 sky130_fd_sc_hd__o21ai_1 _4518_ (.A1(_0516_),
    .A2(_0496_),
    .B1(_1000_),
    .Y(_1001_));
 sky130_fd_sc_hd__a221oi_1 _4519_ (.A1(_0499_),
    .A2(_0488_),
    .B1(_0513_),
    .B2(_0492_),
    .C1(_1001_),
    .Y(_1002_));
 sky130_fd_sc_hd__nand2_1 _4520_ (.A(_0508_),
    .B(_0475_),
    .Y(_1003_));
 sky130_fd_sc_hd__nand2_1 _4521_ (.A(_0512_),
    .B(_0503_),
    .Y(_1004_));
 sky130_fd_sc_hd__or2_1 _4522_ (.A(_0468_),
    .B(_0518_),
    .X(_1005_));
 sky130_fd_sc_hd__o2111a_1 _4523_ (.A1(_0862_),
    .A2(_0506_),
    .B1(_1003_),
    .C1(_1004_),
    .D1(_1005_),
    .X(_1006_));
 sky130_fd_sc_hd__nand2_1 _4524_ (.A(_0530_),
    .B(_0359_),
    .Y(_1007_));
 sky130_fd_sc_hd__nand2_1 _4525_ (.A(_0534_),
    .B(_0525_),
    .Y(_1008_));
 sky130_fd_sc_hd__nand2_1 _4526_ (.A(_1007_),
    .B(_1008_),
    .Y(_1009_));
 sky130_fd_sc_hd__a221oi_1 _4527_ (.A1(_0363_),
    .A2(_0524_),
    .B1(_0689_),
    .B2(_0528_),
    .C1(_1009_),
    .Y(_1010_));
 sky130_fd_sc_hd__and4_1 _4528_ (.A(_0999_),
    .B(_1002_),
    .C(_1006_),
    .D(_1010_),
    .X(_1011_));
 sky130_fd_sc_hd__nand2_1 _4529_ (.A(_0547_),
    .B(\egd_top.BitStream_buffer.BS_buffer[9] ),
    .Y(_1012_));
 sky130_fd_sc_hd__nand2_1 _4530_ (.A(_0551_),
    .B(\egd_top.BitStream_buffer.BS_buffer[7] ),
    .Y(_1013_));
 sky130_fd_sc_hd__or2_1 _4531_ (.A(_0750_),
    .B(_0556_),
    .X(_1014_));
 sky130_fd_sc_hd__o2111a_1 _4532_ (.A1(_0745_),
    .A2(_0545_),
    .B1(_1012_),
    .C1(_1013_),
    .D1(_1014_),
    .X(_1015_));
 sky130_fd_sc_hd__nand2_1 _4533_ (.A(_0563_),
    .B(\egd_top.BitStream_buffer.BS_buffer[13] ),
    .Y(_1016_));
 sky130_fd_sc_hd__nand2_1 _4534_ (.A(_0566_),
    .B(\egd_top.BitStream_buffer.BS_buffer[11] ),
    .Y(_1017_));
 sky130_fd_sc_hd__or2_1 _4535_ (.A(_0593_),
    .B(_0570_),
    .X(_1018_));
 sky130_fd_sc_hd__o2111a_1 _4536_ (.A1(_0756_),
    .A2(_0561_),
    .B1(_1016_),
    .C1(_1017_),
    .D1(_1018_),
    .X(_1019_));
 sky130_fd_sc_hd__or2_1 _4537_ (.A(_0742_),
    .B(_0584_),
    .X(_1020_));
 sky130_fd_sc_hd__o221a_1 _4538_ (.A1(_0541_),
    .A2(_0576_),
    .B1(_0753_),
    .B2(_0580_),
    .C1(_1020_),
    .X(_1021_));
 sky130_fd_sc_hd__inv_2 _4539_ (.A(\egd_top.BitStream_buffer.BS_buffer[16] ),
    .Y(_1022_));
 sky130_fd_sc_hd__o22ai_1 _4540_ (.A1(_0890_),
    .A2(_0595_),
    .B1(_1022_),
    .B2(_0598_),
    .Y(_1023_));
 sky130_fd_sc_hd__a221oi_1 _4541_ (.A1(_0489_),
    .A2(_0589_),
    .B1(_0493_),
    .B2(_0592_),
    .C1(_1023_),
    .Y(_1024_));
 sky130_fd_sc_hd__and4_1 _4542_ (.A(_1015_),
    .B(_1019_),
    .C(_1021_),
    .D(_1024_),
    .X(_1025_));
 sky130_fd_sc_hd__and3_1 _4543_ (.A(_0994_),
    .B(_1011_),
    .C(_1025_),
    .X(_1026_));
 sky130_fd_sc_hd__nand2_1 _4544_ (.A(_0606_),
    .B(_0581_),
    .Y(_1027_));
 sky130_fd_sc_hd__nand3_1 _4545_ (.A(_0961_),
    .B(_1026_),
    .C(_1027_),
    .Y(_1028_));
 sky130_fd_sc_hd__inv_2 _4546_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[12] ),
    .Y(_1029_));
 sky130_fd_sc_hd__a21oi_1 _4547_ (.A1(_1029_),
    .A2(_0898_),
    .B1(_2938_),
    .Y(_1030_));
 sky130_fd_sc_hd__o21a_1 _4548_ (.A1(_3056_),
    .A2(_1028_),
    .B1(_1030_),
    .X(_0294_));
 sky130_fd_sc_hd__inv_2 _4549_ (.A(_3156_),
    .Y(_1031_));
 sky130_fd_sc_hd__o22ai_1 _4550_ (.A1(_0900_),
    .A2(_3084_),
    .B1(_1031_),
    .B2(_3092_),
    .Y(_1032_));
 sky130_fd_sc_hd__a221oi_1 _4551_ (.A1(_3144_),
    .A2(_3068_),
    .B1(_3149_),
    .B2(_3075_),
    .C1(_1032_),
    .Y(_1033_));
 sky130_fd_sc_hd__inv_2 _4552_ (.A(_3129_),
    .Y(_1034_));
 sky130_fd_sc_hd__nand2_1 _4553_ (.A(_3114_),
    .B(_3136_),
    .Y(_1035_));
 sky130_fd_sc_hd__o21ai_1 _4554_ (.A1(_1034_),
    .A2(_3111_),
    .B1(_1035_),
    .Y(_1036_));
 sky130_fd_sc_hd__a221oi_1 _4555_ (.A1(_3134_),
    .A2(_3101_),
    .B1(_3119_),
    .B2(_3106_),
    .C1(_1036_),
    .Y(_1037_));
 sky130_fd_sc_hd__nand2_1 _4556_ (.A(_3128_),
    .B(_3076_),
    .Y(_1038_));
 sky130_fd_sc_hd__nand2_1 _4557_ (.A(_3133_),
    .B(_3057_),
    .Y(_1039_));
 sky130_fd_sc_hd__or2_1 _4558_ (.A(_3086_),
    .B(_3141_),
    .X(_1040_));
 sky130_fd_sc_hd__o2111a_1 _4559_ (.A1(_0764_),
    .A2(_3124_),
    .B1(_1038_),
    .C1(_1039_),
    .D1(_1040_),
    .X(_1041_));
 sky130_fd_sc_hd__nand2_1 _4560_ (.A(_3155_),
    .B(_3247_),
    .Y(_1042_));
 sky130_fd_sc_hd__nand2_1 _4561_ (.A(_3160_),
    .B(_3255_),
    .Y(_1043_));
 sky130_fd_sc_hd__nand2_1 _4562_ (.A(_1042_),
    .B(_1043_),
    .Y(_1044_));
 sky130_fd_sc_hd__a221oi_2 _4563_ (.A1(_3259_),
    .A2(_3148_),
    .B1(_3251_),
    .B2(_3152_),
    .C1(_1044_),
    .Y(_1045_));
 sky130_fd_sc_hd__and4_1 _4564_ (.A(_1033_),
    .B(_1037_),
    .C(_1041_),
    .D(_1045_),
    .X(_1046_));
 sky130_fd_sc_hd__inv_2 _4565_ (.A(\egd_top.BitStream_buffer.BS_buffer[121] ),
    .Y(_1047_));
 sky130_fd_sc_hd__o22ai_1 _4566_ (.A1(_0916_),
    .A2(_3176_),
    .B1(_1047_),
    .B2(_3179_),
    .Y(_1048_));
 sky130_fd_sc_hd__a221oi_1 _4567_ (.A1(_3037_),
    .A2(_3170_),
    .B1(_3040_),
    .B2(_3173_),
    .C1(_1048_),
    .Y(_1049_));
 sky130_fd_sc_hd__nand2_1 _4568_ (.A(_3192_),
    .B(_3050_),
    .Y(_1050_));
 sky130_fd_sc_hd__o21ai_1 _4569_ (.A1(_0790_),
    .A2(_3190_),
    .B1(_1050_),
    .Y(_1051_));
 sky130_fd_sc_hd__a221oi_1 _4570_ (.A1(_3044_),
    .A2(_3184_),
    .B1(_3047_),
    .B2(_3187_),
    .C1(_1051_),
    .Y(_1052_));
 sky130_fd_sc_hd__nand2_1 _4571_ (.A(_3206_),
    .B(_3022_),
    .Y(_1053_));
 sky130_fd_sc_hd__o21ai_1 _4572_ (.A1(_3174_),
    .A2(_3204_),
    .B1(_1053_),
    .Y(_1054_));
 sky130_fd_sc_hd__a221oi_1 _4573_ (.A1(_3025_),
    .A2(_3198_),
    .B1(_3028_),
    .B2(_3201_),
    .C1(_1054_),
    .Y(_1055_));
 sky130_fd_sc_hd__o22ai_1 _4574_ (.A1(_0926_),
    .A2(_3218_),
    .B1(_0578_),
    .B2(_3221_),
    .Y(_1056_));
 sky130_fd_sc_hd__a221oi_1 _4575_ (.A1(_0573_),
    .A2(_3212_),
    .B1(_0581_),
    .B2(_3215_),
    .C1(_1056_),
    .Y(_1057_));
 sky130_fd_sc_hd__and4_1 _4576_ (.A(_1049_),
    .B(_1052_),
    .C(_1055_),
    .D(_1057_),
    .X(_1058_));
 sky130_fd_sc_hd__o22ai_1 _4577_ (.A1(_3287_),
    .A2(_3238_),
    .B1(_3291_),
    .B2(_3241_),
    .Y(_1059_));
 sky130_fd_sc_hd__a221oi_1 _4578_ (.A1(_3278_),
    .A2(_3231_),
    .B1(_3282_),
    .B2(_3235_),
    .C1(_1059_),
    .Y(_1060_));
 sky130_fd_sc_hd__nand2_1 _4579_ (.A(_3246_),
    .B(_3265_),
    .Y(_1061_));
 sky130_fd_sc_hd__nand2_1 _4580_ (.A(_3250_),
    .B(_3275_),
    .Y(_1062_));
 sky130_fd_sc_hd__nand2_1 _4581_ (.A(_3254_),
    .B(_0646_),
    .Y(_1063_));
 sky130_fd_sc_hd__nand2_1 _4582_ (.A(_3258_),
    .B(_3272_),
    .Y(_1064_));
 sky130_fd_sc_hd__and4_1 _4583_ (.A(_1061_),
    .B(_1062_),
    .C(_1063_),
    .D(_1064_),
    .X(_1065_));
 sky130_fd_sc_hd__o22ai_1 _4584_ (.A1(_3236_),
    .A2(_3264_),
    .B1(_3239_),
    .B2(_3268_),
    .Y(_1066_));
 sky130_fd_sc_hd__a22o_1 _4585_ (.A1(_3271_),
    .A2(_3225_),
    .B1(_3274_),
    .B2(_3232_),
    .X(_1067_));
 sky130_fd_sc_hd__nor2_1 _4586_ (.A(_1066_),
    .B(_1067_),
    .Y(_1068_));
 sky130_fd_sc_hd__inv_2 _4587_ (.A(_3322_),
    .Y(_1069_));
 sky130_fd_sc_hd__o22ai_1 _4588_ (.A1(_0940_),
    .A2(_3289_),
    .B1(_1069_),
    .B2(_3293_),
    .Y(_1070_));
 sky130_fd_sc_hd__a221oi_1 _4589_ (.A1(_3331_),
    .A2(_3281_),
    .B1(_3327_),
    .B2(_3285_),
    .C1(_1070_),
    .Y(_1071_));
 sky130_fd_sc_hd__and4_1 _4590_ (.A(_1060_),
    .B(_1065_),
    .C(_1068_),
    .D(_1071_),
    .X(_1072_));
 sky130_fd_sc_hd__nand2_1 _4591_ (.A(_3309_),
    .B(_3357_),
    .Y(_1073_));
 sky130_fd_sc_hd__nand2_1 _4592_ (.A(_3313_),
    .B(_3353_),
    .Y(_1074_));
 sky130_fd_sc_hd__nand2_1 _4593_ (.A(_1073_),
    .B(_1074_),
    .Y(_1075_));
 sky130_fd_sc_hd__a221oi_1 _4594_ (.A1(_0674_),
    .A2(_3303_),
    .B1(_0675_),
    .B2(_3307_),
    .C1(_1075_),
    .Y(_1076_));
 sky130_fd_sc_hd__nand2_1 _4595_ (.A(_3326_),
    .B(_3335_),
    .Y(_1077_));
 sky130_fd_sc_hd__nand2_1 _4596_ (.A(_3330_),
    .B(_3345_),
    .Y(_1078_));
 sky130_fd_sc_hd__nand2_1 _4597_ (.A(_1077_),
    .B(_1078_),
    .Y(_1079_));
 sky130_fd_sc_hd__a221oi_1 _4598_ (.A1(_3341_),
    .A2(_3321_),
    .B1(_3347_),
    .B2(_3324_),
    .C1(_1079_),
    .Y(_1080_));
 sky130_fd_sc_hd__inv_2 _4599_ (.A(\egd_top.BitStream_buffer.BS_buffer[107] ),
    .Y(_1081_));
 sky130_fd_sc_hd__nand2_1 _4600_ (.A(_3340_),
    .B(_3314_),
    .Y(_1082_));
 sky130_fd_sc_hd__nand2_1 _4601_ (.A(_3344_),
    .B(_3297_),
    .Y(_1083_));
 sky130_fd_sc_hd__or2_1 _4602_ (.A(_0819_),
    .B(_3350_),
    .X(_1084_));
 sky130_fd_sc_hd__o2111a_1 _4603_ (.A1(_1081_),
    .A2(_3338_),
    .B1(_1082_),
    .C1(_1083_),
    .D1(_1084_),
    .X(_1085_));
 sky130_fd_sc_hd__nand2_1 _4604_ (.A(_3365_),
    .B(_3013_),
    .Y(_1086_));
 sky130_fd_sc_hd__o21ai_1 _4605_ (.A1(_0922_),
    .A2(_3363_),
    .B1(_1086_),
    .Y(_1087_));
 sky130_fd_sc_hd__a221oi_1 _4606_ (.A1(_2998_),
    .A2(_3356_),
    .B1(_3010_),
    .B2(_3360_),
    .C1(_1087_),
    .Y(_1088_));
 sky130_fd_sc_hd__and4_1 _4607_ (.A(_1076_),
    .B(_1080_),
    .C(_1085_),
    .D(_1088_),
    .X(_1089_));
 sky130_fd_sc_hd__and4_1 _4608_ (.A(_1046_),
    .B(_1058_),
    .C(_1072_),
    .D(_1089_),
    .X(_1090_));
 sky130_fd_sc_hd__nand2_1 _4609_ (.A(_0334_),
    .B(_0380_),
    .Y(_1091_));
 sky130_fd_sc_hd__nand2_1 _4610_ (.A(_0338_),
    .B(_0376_),
    .Y(_1092_));
 sky130_fd_sc_hd__nand2_1 _4611_ (.A(_1091_),
    .B(_1092_),
    .Y(_1093_));
 sky130_fd_sc_hd__a221oi_1 _4612_ (.A1(_0389_),
    .A2(_0328_),
    .B1(_0695_),
    .B2(_0332_),
    .C1(_1093_),
    .Y(_1094_));
 sky130_fd_sc_hd__inv_2 _4613_ (.A(\egd_top.BitStream_buffer.BS_buffer[41] ),
    .Y(_1095_));
 sky130_fd_sc_hd__o22ai_1 _4614_ (.A1(_0966_),
    .A2(_0345_),
    .B1(_1095_),
    .B2(_0349_),
    .Y(_1096_));
 sky130_fd_sc_hd__a22o_1 _4615_ (.A1(_0352_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[42] ),
    .B1(_0355_),
    .B2(_0329_),
    .X(_1097_));
 sky130_fd_sc_hd__nor2_1 _4616_ (.A(_1096_),
    .B(_1097_),
    .Y(_1098_));
 sky130_fd_sc_hd__nand2_1 _4617_ (.A(_0371_),
    .B(_0356_),
    .Y(_1099_));
 sky130_fd_sc_hd__o21ai_1 _4618_ (.A1(_0685_),
    .A2(_0369_),
    .B1(_1099_),
    .Y(_1100_));
 sky130_fd_sc_hd__a221oi_1 _4619_ (.A1(_0691_),
    .A2(_0362_),
    .B1(_0346_),
    .B2(_0366_),
    .C1(_1100_),
    .Y(_1101_));
 sky130_fd_sc_hd__nand2_1 _4620_ (.A(_0388_),
    .B(_0429_),
    .Y(_1102_));
 sky130_fd_sc_hd__o21ai_1 _4621_ (.A1(_0986_),
    .A2(_0386_),
    .B1(_1102_),
    .Y(_1103_));
 sky130_fd_sc_hd__a221oi_1 _4622_ (.A1(_0437_),
    .A2(_0379_),
    .B1(_0443_),
    .B2(_0383_),
    .C1(_1103_),
    .Y(_1104_));
 sky130_fd_sc_hd__and4_1 _4623_ (.A(_1094_),
    .B(_1098_),
    .C(_1101_),
    .D(_1104_),
    .X(_1105_));
 sky130_fd_sc_hd__nand2_1 _4624_ (.A(_0399_),
    .B(_0421_),
    .Y(_1106_));
 sky130_fd_sc_hd__nand2_1 _4625_ (.A(_0403_),
    .B(_0417_),
    .Y(_1107_));
 sky130_fd_sc_hd__or2_1 _4626_ (.A(_0412_),
    .B(_0408_),
    .X(_1108_));
 sky130_fd_sc_hd__o2111a_1 _4627_ (.A1(_0424_),
    .A2(_0397_),
    .B1(_1106_),
    .C1(_1107_),
    .D1(_1108_),
    .X(_1109_));
 sky130_fd_sc_hd__nand2_1 _4628_ (.A(_0416_),
    .B(_0447_),
    .Y(_1110_));
 sky130_fd_sc_hd__nand2_1 _4629_ (.A(_0420_),
    .B(_0461_),
    .Y(_1111_));
 sky130_fd_sc_hd__or2_1 _4630_ (.A(_0848_),
    .B(_0426_),
    .X(_1112_));
 sky130_fd_sc_hd__o2111a_1 _4631_ (.A1(_0456_),
    .A2(_0414_),
    .B1(_1110_),
    .C1(_1111_),
    .D1(_1112_),
    .X(_1113_));
 sky130_fd_sc_hd__inv_2 _4632_ (.A(\egd_top.BitStream_buffer.BS_buffer[52] ),
    .Y(_1114_));
 sky130_fd_sc_hd__nand2_1 _4633_ (.A(_0442_),
    .B(_0703_),
    .Y(_1115_));
 sky130_fd_sc_hd__o21ai_1 _4634_ (.A1(_1114_),
    .A2(_0440_),
    .B1(_1115_),
    .Y(_1116_));
 sky130_fd_sc_hd__a221oi_1 _4635_ (.A1(_0400_),
    .A2(_0432_),
    .B1(_0701_),
    .B2(_0436_),
    .C1(_1116_),
    .Y(_1117_));
 sky130_fd_sc_hd__nand2_1 _4636_ (.A(_0460_),
    .B(_3095_),
    .Y(_1118_));
 sky130_fd_sc_hd__o21ai_1 _4637_ (.A1(_0903_),
    .A2(_0458_),
    .B1(_1118_),
    .Y(_1119_));
 sky130_fd_sc_hd__a221oi_1 _4638_ (.A1(_3107_),
    .A2(_0450_),
    .B1(_3115_),
    .B2(_0454_),
    .C1(_1119_),
    .Y(_1120_));
 sky130_fd_sc_hd__and4_1 _4639_ (.A(_1109_),
    .B(_1113_),
    .C(_1117_),
    .D(_1120_),
    .X(_1121_));
 sky130_fd_sc_hd__and2_1 _4640_ (.A(_1105_),
    .B(_1121_),
    .X(_1122_));
 sky130_fd_sc_hd__inv_2 _4641_ (.A(\egd_top.BitStream_buffer.BS_buffer[28] ),
    .Y(_1123_));
 sky130_fd_sc_hd__nand2_1 _4642_ (.A(_0474_),
    .B(_0531_),
    .Y(_1124_));
 sky130_fd_sc_hd__a22o_1 _4643_ (.A1(_0478_),
    .A2(_0521_),
    .B1(_0481_),
    .B2(_0525_),
    .X(_1125_));
 sky130_fd_sc_hd__inv_2 _4644_ (.A(_1125_),
    .Y(_1126_));
 sky130_fd_sc_hd__o211a_1 _4645_ (.A1(_1123_),
    .A2(_0472_),
    .B1(_1124_),
    .C1(_1126_),
    .X(_1127_));
 sky130_fd_sc_hd__nand2_1 _4646_ (.A(_0498_),
    .B(_0503_),
    .Y(_1128_));
 sky130_fd_sc_hd__o21ai_1 _4647_ (.A1(_0734_),
    .A2(_0496_),
    .B1(_1128_),
    .Y(_1129_));
 sky130_fd_sc_hd__a221oi_1 _4648_ (.A1(_0513_),
    .A2(_0488_),
    .B1(_0515_),
    .B2(_0492_),
    .C1(_1129_),
    .Y(_1130_));
 sky130_fd_sc_hd__nand2_1 _4649_ (.A(_0508_),
    .B(_0479_),
    .Y(_1131_));
 sky130_fd_sc_hd__nand2_1 _4650_ (.A(_0512_),
    .B(_0467_),
    .Y(_1132_));
 sky130_fd_sc_hd__or2_1 _4651_ (.A(_0723_),
    .B(_0518_),
    .X(_1133_));
 sky130_fd_sc_hd__o2111a_1 _4652_ (.A1(_0995_),
    .A2(_0506_),
    .B1(_1131_),
    .C1(_1132_),
    .D1(_1133_),
    .X(_1134_));
 sky130_fd_sc_hd__nand2_1 _4653_ (.A(_0530_),
    .B(_0363_),
    .Y(_1135_));
 sky130_fd_sc_hd__nand2_1 _4654_ (.A(_0534_),
    .B(_0359_),
    .Y(_1136_));
 sky130_fd_sc_hd__nand2_1 _4655_ (.A(_1135_),
    .B(_1136_),
    .Y(_1137_));
 sky130_fd_sc_hd__a221oi_1 _4656_ (.A1(_0689_),
    .A2(_0524_),
    .B1(_0372_),
    .B2(_0528_),
    .C1(_1137_),
    .Y(_1138_));
 sky130_fd_sc_hd__and4_1 _4657_ (.A(_1127_),
    .B(_1130_),
    .C(_1134_),
    .D(_1138_),
    .X(_1139_));
 sky130_fd_sc_hd__nand2_1 _4658_ (.A(_0547_),
    .B(\egd_top.BitStream_buffer.BS_buffer[10] ),
    .Y(_1140_));
 sky130_fd_sc_hd__nand2_1 _4659_ (.A(_0551_),
    .B(\egd_top.BitStream_buffer.BS_buffer[8] ),
    .Y(_1141_));
 sky130_fd_sc_hd__or2_1 _4660_ (.A(_0559_),
    .B(_0556_),
    .X(_1142_));
 sky130_fd_sc_hd__o2111a_1 _4661_ (.A1(_0568_),
    .A2(_0545_),
    .B1(_1140_),
    .C1(_1141_),
    .D1(_1142_),
    .X(_1143_));
 sky130_fd_sc_hd__nand2_1 _4662_ (.A(_0563_),
    .B(\egd_top.BitStream_buffer.BS_buffer[14] ),
    .Y(_1144_));
 sky130_fd_sc_hd__nand2_1 _4663_ (.A(_0566_),
    .B(\egd_top.BitStream_buffer.BS_buffer[12] ),
    .Y(_1145_));
 sky130_fd_sc_hd__or2_1 _4664_ (.A(_0596_),
    .B(_0570_),
    .X(_1146_));
 sky130_fd_sc_hd__o2111a_1 _4665_ (.A1(_0890_),
    .A2(_0561_),
    .B1(_1144_),
    .C1(_1145_),
    .D1(_1146_),
    .X(_1147_));
 sky130_fd_sc_hd__or2_1 _4666_ (.A(_0554_),
    .B(_0584_),
    .X(_1148_));
 sky130_fd_sc_hd__o221a_1 _4667_ (.A1(_0742_),
    .A2(_0576_),
    .B1(_0541_),
    .B2(_0580_),
    .C1(_1148_),
    .X(_1149_));
 sky130_fd_sc_hd__inv_2 _4668_ (.A(_0489_),
    .Y(_1150_));
 sky130_fd_sc_hd__o22ai_1 _4669_ (.A1(_1022_),
    .A2(_0595_),
    .B1(_1150_),
    .B2(_0598_),
    .Y(_1151_));
 sky130_fd_sc_hd__a221oi_1 _4670_ (.A1(_0493_),
    .A2(_0589_),
    .B1(_0499_),
    .B2(_0592_),
    .C1(_1151_),
    .Y(_1152_));
 sky130_fd_sc_hd__and4_1 _4671_ (.A(_1143_),
    .B(_1147_),
    .C(_1149_),
    .D(_1152_),
    .X(_1153_));
 sky130_fd_sc_hd__and3_1 _4672_ (.A(_1122_),
    .B(_1139_),
    .C(_1153_),
    .X(_1154_));
 sky130_fd_sc_hd__nand2_1 _4673_ (.A(_0606_),
    .B(_0552_),
    .Y(_1155_));
 sky130_fd_sc_hd__nand3_1 _4674_ (.A(_1090_),
    .B(_1154_),
    .C(_1155_),
    .Y(_1156_));
 sky130_fd_sc_hd__inv_4 _4675_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[11] ),
    .Y(_1157_));
 sky130_fd_sc_hd__a21oi_1 _4676_ (.A1(_1157_),
    .A2(_0898_),
    .B1(_2938_),
    .Y(_1158_));
 sky130_fd_sc_hd__o21a_1 _4677_ (.A1(_3056_),
    .A2(_1156_),
    .B1(_1158_),
    .X(_0293_));
 sky130_fd_sc_hd__inv_2 _4678_ (.A(_3144_),
    .Y(_1159_));
 sky130_fd_sc_hd__o22ai_1 _4679_ (.A1(_1031_),
    .A2(_3084_),
    .B1(_1159_),
    .B2(_3092_),
    .Y(_1160_));
 sky130_fd_sc_hd__a221oi_1 _4680_ (.A1(_3149_),
    .A2(_3068_),
    .B1(_3255_),
    .B2(_3075_),
    .C1(_1160_),
    .Y(_1161_));
 sky130_fd_sc_hd__nand2_1 _4681_ (.A(_3114_),
    .B(_3134_),
    .Y(_1162_));
 sky130_fd_sc_hd__o21ai_1 _4682_ (.A1(_3137_),
    .A2(_3111_),
    .B1(_1162_),
    .Y(_1163_));
 sky130_fd_sc_hd__a221oi_1 _4683_ (.A1(_3119_),
    .A2(_3101_),
    .B1(_3076_),
    .B2(_3106_),
    .C1(_1163_),
    .Y(_1164_));
 sky130_fd_sc_hd__nand2_1 _4684_ (.A(_3128_),
    .B(_3085_),
    .Y(_1165_));
 sky130_fd_sc_hd__nand2_1 _4685_ (.A(_3133_),
    .B(_3069_),
    .Y(_1166_));
 sky130_fd_sc_hd__or2_1 _4686_ (.A(_0611_),
    .B(_3141_),
    .X(_1167_));
 sky130_fd_sc_hd__o2111a_1 _4687_ (.A1(_0900_),
    .A2(_3124_),
    .B1(_1165_),
    .C1(_1166_),
    .D1(_1167_),
    .X(_1168_));
 sky130_fd_sc_hd__nand2_1 _4688_ (.A(_3155_),
    .B(_3259_),
    .Y(_1169_));
 sky130_fd_sc_hd__nand2_1 _4689_ (.A(_3160_),
    .B(_3247_),
    .Y(_1170_));
 sky130_fd_sc_hd__nand2_1 _4690_ (.A(_1169_),
    .B(_1170_),
    .Y(_1171_));
 sky130_fd_sc_hd__a221oi_2 _4691_ (.A1(_3251_),
    .A2(_3148_),
    .B1(_0646_),
    .B2(_3152_),
    .C1(_1171_),
    .Y(_1172_));
 sky130_fd_sc_hd__and4_1 _4692_ (.A(_1161_),
    .B(_1164_),
    .C(_1168_),
    .D(_1172_),
    .X(_1173_));
 sky130_fd_sc_hd__inv_2 _4693_ (.A(\egd_top.BitStream_buffer.BS_buffer[122] ),
    .Y(_1174_));
 sky130_fd_sc_hd__o22ai_1 _4694_ (.A1(_1047_),
    .A2(_3176_),
    .B1(_1174_),
    .B2(_3179_),
    .Y(_1175_));
 sky130_fd_sc_hd__a221oi_1 _4695_ (.A1(_3040_),
    .A2(_3170_),
    .B1(_3044_),
    .B2(_3173_),
    .C1(_1175_),
    .Y(_1176_));
 sky130_fd_sc_hd__nand2_1 _4696_ (.A(_3192_),
    .B(_3053_),
    .Y(_1177_));
 sky130_fd_sc_hd__o21ai_1 _4697_ (.A1(_0926_),
    .A2(_3190_),
    .B1(_1177_),
    .Y(_1178_));
 sky130_fd_sc_hd__a221oi_1 _4698_ (.A1(_3047_),
    .A2(_3184_),
    .B1(_3050_),
    .B2(_3187_),
    .C1(_1178_),
    .Y(_1179_));
 sky130_fd_sc_hd__nand2_1 _4699_ (.A(_3206_),
    .B(_3025_),
    .Y(_1180_));
 sky130_fd_sc_hd__o21ai_1 _4700_ (.A1(_3177_),
    .A2(_3204_),
    .B1(_1180_),
    .Y(_1181_));
 sky130_fd_sc_hd__a221oi_2 _4701_ (.A1(_3028_),
    .A2(_3198_),
    .B1(_3031_),
    .B2(_3201_),
    .C1(_1181_),
    .Y(_1182_));
 sky130_fd_sc_hd__o22ai_1 _4702_ (.A1(_0578_),
    .A2(_3218_),
    .B1(_0574_),
    .B2(_3221_),
    .Y(_1183_));
 sky130_fd_sc_hd__a221oi_1 _4703_ (.A1(_0581_),
    .A2(_3212_),
    .B1(_0552_),
    .B2(_3215_),
    .C1(_1183_),
    .Y(_1184_));
 sky130_fd_sc_hd__and4_1 _4704_ (.A(_1176_),
    .B(_1179_),
    .C(_1182_),
    .D(_1184_),
    .X(_1185_));
 sky130_fd_sc_hd__o22ai_1 _4705_ (.A1(_3291_),
    .A2(_3238_),
    .B1(_0656_),
    .B2(_3241_),
    .Y(_1186_));
 sky130_fd_sc_hd__a221oi_1 _4706_ (.A1(_3282_),
    .A2(_3231_),
    .B1(_3318_),
    .B2(_3235_),
    .C1(_1186_),
    .Y(_1187_));
 sky130_fd_sc_hd__nand2_1 _4707_ (.A(_3246_),
    .B(_3272_),
    .Y(_1188_));
 sky130_fd_sc_hd__nand2_1 _4708_ (.A(_3250_),
    .B(_0653_),
    .Y(_1189_));
 sky130_fd_sc_hd__nand2_1 _4709_ (.A(_3254_),
    .B(_3265_),
    .Y(_1190_));
 sky130_fd_sc_hd__nand2_1 _4710_ (.A(_3258_),
    .B(\egd_top.BitStream_buffer.BS_buffer[87] ),
    .Y(_1191_));
 sky130_fd_sc_hd__and4_1 _4711_ (.A(_1188_),
    .B(_1189_),
    .C(_1190_),
    .D(_1191_),
    .X(_1192_));
 sky130_fd_sc_hd__o22ai_1 _4712_ (.A1(_3239_),
    .A2(_3264_),
    .B1(_0642_),
    .B2(_3268_),
    .Y(_1193_));
 sky130_fd_sc_hd__a22o_1 _4713_ (.A1(_3271_),
    .A2(_3232_),
    .B1(_3274_),
    .B2(_3286_),
    .X(_1194_));
 sky130_fd_sc_hd__nor2_1 _4714_ (.A(_1193_),
    .B(_1194_),
    .Y(_1195_));
 sky130_fd_sc_hd__inv_2 _4715_ (.A(_3331_),
    .Y(_1196_));
 sky130_fd_sc_hd__o22ai_1 _4716_ (.A1(_1069_),
    .A2(_3289_),
    .B1(_1196_),
    .B2(_3293_),
    .Y(_1197_));
 sky130_fd_sc_hd__a221oi_1 _4717_ (.A1(_3327_),
    .A2(_3281_),
    .B1(_3341_),
    .B2(_3285_),
    .C1(_1197_),
    .Y(_1198_));
 sky130_fd_sc_hd__and4_1 _4718_ (.A(_1187_),
    .B(_1192_),
    .C(_1195_),
    .D(_1198_),
    .X(_1199_));
 sky130_fd_sc_hd__nand2_1 _4719_ (.A(_3309_),
    .B(_0674_),
    .Y(_1200_));
 sky130_fd_sc_hd__nand2_1 _4720_ (.A(_3313_),
    .B(_3357_),
    .Y(_1201_));
 sky130_fd_sc_hd__nand2_1 _4721_ (.A(_1200_),
    .B(_1201_),
    .Y(_1202_));
 sky130_fd_sc_hd__a221oi_1 _4722_ (.A1(_0675_),
    .A2(_3303_),
    .B1(_2998_),
    .B2(_3307_),
    .C1(_1202_),
    .Y(_1203_));
 sky130_fd_sc_hd__nand2_1 _4723_ (.A(_3326_),
    .B(_3314_),
    .Y(_1204_));
 sky130_fd_sc_hd__nand2_1 _4724_ (.A(_3330_),
    .B(_3335_),
    .Y(_1205_));
 sky130_fd_sc_hd__nand2_1 _4725_ (.A(_1204_),
    .B(_1205_),
    .Y(_1206_));
 sky130_fd_sc_hd__a221oi_1 _4726_ (.A1(_3347_),
    .A2(_3321_),
    .B1(_3345_),
    .B2(_3324_),
    .C1(_1206_),
    .Y(_1207_));
 sky130_fd_sc_hd__inv_2 _4727_ (.A(\egd_top.BitStream_buffer.BS_buffer[108] ),
    .Y(_1208_));
 sky130_fd_sc_hd__nand2_1 _4728_ (.A(_3340_),
    .B(_3310_),
    .Y(_1209_));
 sky130_fd_sc_hd__nand2_1 _4729_ (.A(_3344_),
    .B(_3304_),
    .Y(_1210_));
 sky130_fd_sc_hd__or2_1 _4730_ (.A(_0952_),
    .B(_3350_),
    .X(_1211_));
 sky130_fd_sc_hd__o2111a_1 _4731_ (.A1(_1208_),
    .A2(_3338_),
    .B1(_1209_),
    .C1(_1210_),
    .D1(_1211_),
    .X(_1212_));
 sky130_fd_sc_hd__nand2_1 _4732_ (.A(_3365_),
    .B(_3016_),
    .Y(_1213_));
 sky130_fd_sc_hd__o21ai_1 _4733_ (.A1(_3174_),
    .A2(_3363_),
    .B1(_1213_),
    .Y(_1214_));
 sky130_fd_sc_hd__a221oi_2 _4734_ (.A1(_3010_),
    .A2(_3356_),
    .B1(_3013_),
    .B2(_3360_),
    .C1(_1214_),
    .Y(_1215_));
 sky130_fd_sc_hd__and4_1 _4735_ (.A(_1203_),
    .B(_1207_),
    .C(_1212_),
    .D(_1215_),
    .X(_1216_));
 sky130_fd_sc_hd__and4_1 _4736_ (.A(_1173_),
    .B(_1185_),
    .C(_1199_),
    .D(_1216_),
    .X(_1217_));
 sky130_fd_sc_hd__nand2_1 _4737_ (.A(_0334_),
    .B(_0389_),
    .Y(_1218_));
 sky130_fd_sc_hd__nand2_1 _4738_ (.A(_0338_),
    .B(_0380_),
    .Y(_1219_));
 sky130_fd_sc_hd__nand2_1 _4739_ (.A(_1218_),
    .B(_1219_),
    .Y(_1220_));
 sky130_fd_sc_hd__a221oi_1 _4740_ (.A1(_0695_),
    .A2(_0328_),
    .B1(_0437_),
    .B2(_0332_),
    .C1(_1220_),
    .Y(_1221_));
 sky130_fd_sc_hd__inv_2 _4741_ (.A(\egd_top.BitStream_buffer.BS_buffer[42] ),
    .Y(_1222_));
 sky130_fd_sc_hd__o22ai_1 _4742_ (.A1(_1095_),
    .A2(_0345_),
    .B1(_1222_),
    .B2(_0349_),
    .Y(_1223_));
 sky130_fd_sc_hd__a22o_1 _4743_ (.A1(_0352_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[43] ),
    .B1(_0355_),
    .B2(_0376_),
    .X(_1224_));
 sky130_fd_sc_hd__nor2_1 _4744_ (.A(_1223_),
    .B(_1224_),
    .Y(_1225_));
 sky130_fd_sc_hd__nand2_1 _4745_ (.A(_0371_),
    .B(_0339_),
    .Y(_1226_));
 sky130_fd_sc_hd__o21ai_1 _4746_ (.A1(_0833_),
    .A2(_0369_),
    .B1(_1226_),
    .Y(_1227_));
 sky130_fd_sc_hd__a221oi_1 _4747_ (.A1(_0346_),
    .A2(_0362_),
    .B1(_0353_),
    .B2(_0366_),
    .C1(_1227_),
    .Y(_1228_));
 sky130_fd_sc_hd__nand2_1 _4748_ (.A(_0388_),
    .B(_0433_),
    .Y(_1229_));
 sky130_fd_sc_hd__o21ai_1 _4749_ (.A1(_1114_),
    .A2(_0386_),
    .B1(_1229_),
    .Y(_1230_));
 sky130_fd_sc_hd__a221oi_2 _4750_ (.A1(_0443_),
    .A2(_0379_),
    .B1(_0429_),
    .B2(_0383_),
    .C1(_1230_),
    .Y(_1231_));
 sky130_fd_sc_hd__and4_1 _4751_ (.A(_1221_),
    .B(_1225_),
    .C(_1228_),
    .D(_1231_),
    .X(_1232_));
 sky130_fd_sc_hd__nand2_1 _4752_ (.A(_0399_),
    .B(_0411_),
    .Y(_1233_));
 sky130_fd_sc_hd__nand2_1 _4753_ (.A(_0403_),
    .B(_0423_),
    .Y(_1234_));
 sky130_fd_sc_hd__or2_1 _4754_ (.A(_0708_),
    .B(_0408_),
    .X(_1235_));
 sky130_fd_sc_hd__o2111a_1 _4755_ (.A1(_0711_),
    .A2(_0397_),
    .B1(_1233_),
    .C1(_1234_),
    .D1(_1235_),
    .X(_1236_));
 sky130_fd_sc_hd__nand2_1 _4756_ (.A(_0416_),
    .B(_0451_),
    .Y(_1237_));
 sky130_fd_sc_hd__nand2_1 _4757_ (.A(_0420_),
    .B(_0455_),
    .Y(_1238_));
 sky130_fd_sc_hd__or2_1 _4758_ (.A(_0981_),
    .B(_0426_),
    .X(_1239_));
 sky130_fd_sc_hd__o2111a_1 _4759_ (.A1(_3108_),
    .A2(_0414_),
    .B1(_1237_),
    .C1(_1238_),
    .D1(_1239_),
    .X(_1240_));
 sky130_fd_sc_hd__nand2_1 _4760_ (.A(_0442_),
    .B(\egd_top.BitStream_buffer.BS_buffer[54] ),
    .Y(_1241_));
 sky130_fd_sc_hd__o21ai_1 _4761_ (.A1(_0394_),
    .A2(_0440_),
    .B1(_1241_),
    .Y(_1242_));
 sky130_fd_sc_hd__a221oi_1 _4762_ (.A1(_0701_),
    .A2(_0432_),
    .B1(_0417_),
    .B2(_0436_),
    .C1(_1242_),
    .Y(_1243_));
 sky130_fd_sc_hd__nand2_1 _4763_ (.A(_0460_),
    .B(_3102_),
    .Y(_1244_));
 sky130_fd_sc_hd__o21ai_1 _4764_ (.A1(_1034_),
    .A2(_0458_),
    .B1(_1244_),
    .Y(_1245_));
 sky130_fd_sc_hd__a221oi_1 _4765_ (.A1(_3115_),
    .A2(_0450_),
    .B1(_3095_),
    .B2(_0454_),
    .C1(_1245_),
    .Y(_1246_));
 sky130_fd_sc_hd__and4_1 _4766_ (.A(_1236_),
    .B(_1240_),
    .C(_1243_),
    .D(_1246_),
    .X(_1247_));
 sky130_fd_sc_hd__and2_1 _4767_ (.A(_1232_),
    .B(_1247_),
    .X(_1248_));
 sky130_fd_sc_hd__inv_2 _4768_ (.A(\egd_top.BitStream_buffer.BS_buffer[29] ),
    .Y(_1249_));
 sky130_fd_sc_hd__nand2_1 _4769_ (.A(_0474_),
    .B(_0521_),
    .Y(_1250_));
 sky130_fd_sc_hd__a22o_1 _4770_ (.A1(_0478_),
    .A2(_0525_),
    .B1(_0481_),
    .B2(_0359_),
    .X(_1251_));
 sky130_fd_sc_hd__inv_2 _4771_ (.A(_1251_),
    .Y(_1252_));
 sky130_fd_sc_hd__o211a_1 _4772_ (.A1(_1249_),
    .A2(_0472_),
    .B1(_1250_),
    .C1(_1252_),
    .X(_1253_));
 sky130_fd_sc_hd__nand2_1 _4773_ (.A(_0498_),
    .B(_0467_),
    .Y(_1254_));
 sky130_fd_sc_hd__o21ai_1 _4774_ (.A1(_0504_),
    .A2(_0496_),
    .B1(_1254_),
    .Y(_1255_));
 sky130_fd_sc_hd__a221oi_1 _4775_ (.A1(_0515_),
    .A2(_0488_),
    .B1(_0509_),
    .B2(_0492_),
    .C1(_1255_),
    .Y(_1256_));
 sky130_fd_sc_hd__nand2_1 _4776_ (.A(_0508_),
    .B(_0482_),
    .Y(_1257_));
 sky130_fd_sc_hd__nand2_1 _4777_ (.A(_0512_),
    .B(_0475_),
    .Y(_1258_));
 sky130_fd_sc_hd__or2_1 _4778_ (.A(_0862_),
    .B(_0518_),
    .X(_1259_));
 sky130_fd_sc_hd__o2111a_1 _4779_ (.A1(_1123_),
    .A2(_0506_),
    .B1(_1257_),
    .C1(_1258_),
    .D1(_1259_),
    .X(_1260_));
 sky130_fd_sc_hd__nand2_1 _4780_ (.A(_0530_),
    .B(_0689_),
    .Y(_1261_));
 sky130_fd_sc_hd__nand2_1 _4781_ (.A(_0534_),
    .B(_0363_),
    .Y(_1262_));
 sky130_fd_sc_hd__nand2_1 _4782_ (.A(_1261_),
    .B(_1262_),
    .Y(_1263_));
 sky130_fd_sc_hd__a221oi_1 _4783_ (.A1(_0372_),
    .A2(_0524_),
    .B1(_0691_),
    .B2(_0528_),
    .C1(_1263_),
    .Y(_1264_));
 sky130_fd_sc_hd__and4_1 _4784_ (.A(_1253_),
    .B(_1256_),
    .C(_1260_),
    .D(_1264_),
    .X(_1265_));
 sky130_fd_sc_hd__nand2_1 _4785_ (.A(_0547_),
    .B(\egd_top.BitStream_buffer.BS_buffer[11] ),
    .Y(_1266_));
 sky130_fd_sc_hd__nand2_1 _4786_ (.A(_0551_),
    .B(\egd_top.BitStream_buffer.BS_buffer[9] ),
    .Y(_1267_));
 sky130_fd_sc_hd__or2_1 _4787_ (.A(_0593_),
    .B(_0556_),
    .X(_1268_));
 sky130_fd_sc_hd__o2111a_1 _4788_ (.A1(_0750_),
    .A2(_0545_),
    .B1(_1266_),
    .C1(_1267_),
    .D1(_1268_),
    .X(_1269_));
 sky130_fd_sc_hd__nand2_1 _4789_ (.A(_0563_),
    .B(\egd_top.BitStream_buffer.BS_buffer[15] ),
    .Y(_1270_));
 sky130_fd_sc_hd__nand2_1 _4790_ (.A(_0566_),
    .B(\egd_top.BitStream_buffer.BS_buffer[13] ),
    .Y(_1271_));
 sky130_fd_sc_hd__or2_1 _4791_ (.A(_0756_),
    .B(_0570_),
    .X(_1272_));
 sky130_fd_sc_hd__o2111a_1 _4792_ (.A1(_1022_),
    .A2(_0561_),
    .B1(_1270_),
    .C1(_1271_),
    .D1(_1272_),
    .X(_1273_));
 sky130_fd_sc_hd__or2_1 _4793_ (.A(_0745_),
    .B(_0584_),
    .X(_1274_));
 sky130_fd_sc_hd__o221a_1 _4794_ (.A1(_0554_),
    .A2(_0576_),
    .B1(_0742_),
    .B2(_0580_),
    .C1(_1274_),
    .X(_1275_));
 sky130_fd_sc_hd__o22ai_1 _4795_ (.A1(_1150_),
    .A2(_0595_),
    .B1(_0494_),
    .B2(_0598_),
    .Y(_1276_));
 sky130_fd_sc_hd__a221oi_1 _4796_ (.A1(_0499_),
    .A2(_0589_),
    .B1(_0513_),
    .B2(_0592_),
    .C1(_1276_),
    .Y(_1277_));
 sky130_fd_sc_hd__and4_1 _4797_ (.A(_1269_),
    .B(_1273_),
    .C(_1275_),
    .D(_1277_),
    .X(_1278_));
 sky130_fd_sc_hd__and3_1 _4798_ (.A(_1248_),
    .B(_1265_),
    .C(_1278_),
    .X(_1279_));
 sky130_fd_sc_hd__nand2_1 _4799_ (.A(_0606_),
    .B(_0540_),
    .Y(_1280_));
 sky130_fd_sc_hd__nand3_1 _4800_ (.A(_1217_),
    .B(_1279_),
    .C(_1280_),
    .Y(_1281_));
 sky130_fd_sc_hd__inv_2 _4801_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[10] ),
    .Y(_1282_));
 sky130_fd_sc_hd__a21oi_1 _4802_ (.A1(_1282_),
    .A2(_0898_),
    .B1(_2938_),
    .Y(_1283_));
 sky130_fd_sc_hd__o21a_1 _4803_ (.A1(_3056_),
    .A2(_1281_),
    .B1(_1283_),
    .X(_0292_));
 sky130_fd_sc_hd__inv_2 _4804_ (.A(\egd_top.BitStream_buffer.BS_buffer[79] ),
    .Y(_1284_));
 sky130_fd_sc_hd__o22ai_1 _4805_ (.A1(_1159_),
    .A2(_3084_),
    .B1(_1284_),
    .B2(_3092_),
    .Y(_1285_));
 sky130_fd_sc_hd__a221oi_1 _4806_ (.A1(_3255_),
    .A2(_3068_),
    .B1(_3247_),
    .B2(_3075_),
    .C1(_1285_),
    .Y(_1286_));
 sky130_fd_sc_hd__nand2_1 _4807_ (.A(_3114_),
    .B(_3119_),
    .Y(_1287_));
 sky130_fd_sc_hd__o21ai_1 _4808_ (.A1(_0620_),
    .A2(_3111_),
    .B1(_1287_),
    .Y(_1288_));
 sky130_fd_sc_hd__a221oi_1 _4809_ (.A1(_3076_),
    .A2(_3101_),
    .B1(_3085_),
    .B2(_3106_),
    .C1(_1288_),
    .Y(_1289_));
 sky130_fd_sc_hd__nand2_1 _4810_ (.A(_3128_),
    .B(_3057_),
    .Y(_1290_));
 sky130_fd_sc_hd__nand2_1 _4811_ (.A(_3133_),
    .B(_3161_),
    .Y(_1291_));
 sky130_fd_sc_hd__or2_1 _4812_ (.A(_0764_),
    .B(_3141_),
    .X(_1292_));
 sky130_fd_sc_hd__o2111a_1 _4813_ (.A1(_1031_),
    .A2(_3124_),
    .B1(_1290_),
    .C1(_1291_),
    .D1(_1292_),
    .X(_1293_));
 sky130_fd_sc_hd__nand2_1 _4814_ (.A(_3155_),
    .B(_3251_),
    .Y(_1294_));
 sky130_fd_sc_hd__nand2_1 _4815_ (.A(_3160_),
    .B(_3259_),
    .Y(_1295_));
 sky130_fd_sc_hd__nand2_1 _4816_ (.A(_1294_),
    .B(_1295_),
    .Y(_1296_));
 sky130_fd_sc_hd__a221oi_1 _4817_ (.A1(_0646_),
    .A2(_3148_),
    .B1(_3265_),
    .B2(_3152_),
    .C1(_1296_),
    .Y(_1297_));
 sky130_fd_sc_hd__and4_1 _4818_ (.A(_1286_),
    .B(_1289_),
    .C(_1293_),
    .D(_1297_),
    .X(_1298_));
 sky130_fd_sc_hd__o22ai_1 _4819_ (.A1(_1174_),
    .A2(_3176_),
    .B1(_3188_),
    .B2(_3179_),
    .Y(_1299_));
 sky130_fd_sc_hd__a221oi_1 _4820_ (.A1(_3044_),
    .A2(_3170_),
    .B1(_3047_),
    .B2(_3173_),
    .C1(_1299_),
    .Y(_1300_));
 sky130_fd_sc_hd__nand2_1 _4821_ (.A(_3192_),
    .B(_0607_),
    .Y(_1301_));
 sky130_fd_sc_hd__o21ai_1 _4822_ (.A1(_0578_),
    .A2(_3190_),
    .B1(_1301_),
    .Y(_1302_));
 sky130_fd_sc_hd__a221oi_1 _4823_ (.A1(_3050_),
    .A2(_3184_),
    .B1(_3053_),
    .B2(_3187_),
    .C1(_1302_),
    .Y(_1303_));
 sky130_fd_sc_hd__nand2_1 _4824_ (.A(_3206_),
    .B(_3028_),
    .Y(_1304_));
 sky130_fd_sc_hd__o21ai_1 _4825_ (.A1(_0628_),
    .A2(_3204_),
    .B1(_1304_),
    .Y(_1305_));
 sky130_fd_sc_hd__a221oi_1 _4826_ (.A1(_3031_),
    .A2(_3198_),
    .B1(_3034_),
    .B2(_3201_),
    .C1(_1305_),
    .Y(_1306_));
 sky130_fd_sc_hd__o22ai_1 _4827_ (.A1(_0574_),
    .A2(_3218_),
    .B1(_0582_),
    .B2(_3221_),
    .Y(_1307_));
 sky130_fd_sc_hd__a221oi_1 _4828_ (.A1(_0552_),
    .A2(_3212_),
    .B1(_0540_),
    .B2(_3215_),
    .C1(_1307_),
    .Y(_1308_));
 sky130_fd_sc_hd__and4_1 _4829_ (.A(_1300_),
    .B(_1303_),
    .C(_1306_),
    .D(_1308_),
    .X(_1309_));
 sky130_fd_sc_hd__o22ai_1 _4830_ (.A1(_0656_),
    .A2(_3238_),
    .B1(_0807_),
    .B2(_3241_),
    .Y(_1310_));
 sky130_fd_sc_hd__a221oi_1 _4831_ (.A1(_3318_),
    .A2(_3231_),
    .B1(_3322_),
    .B2(_3235_),
    .C1(_1310_),
    .Y(_1311_));
 sky130_fd_sc_hd__nand2_1 _4832_ (.A(_3246_),
    .B(_3275_),
    .Y(_1312_));
 sky130_fd_sc_hd__nand2_1 _4833_ (.A(_3250_),
    .B(_0804_),
    .Y(_1313_));
 sky130_fd_sc_hd__nand2_1 _4834_ (.A(_3254_),
    .B(_3272_),
    .Y(_1314_));
 sky130_fd_sc_hd__nand2_1 _4835_ (.A(_3258_),
    .B(\egd_top.BitStream_buffer.BS_buffer[88] ),
    .Y(_1315_));
 sky130_fd_sc_hd__and4_1 _4836_ (.A(_1312_),
    .B(_1313_),
    .C(_1314_),
    .D(_1315_),
    .X(_1316_));
 sky130_fd_sc_hd__o22ai_1 _4837_ (.A1(_0642_),
    .A2(_3264_),
    .B1(_0794_),
    .B2(_3268_),
    .Y(_1317_));
 sky130_fd_sc_hd__a22o_1 _4838_ (.A1(_3271_),
    .A2(_3286_),
    .B1(_3274_),
    .B2(_3290_),
    .X(_1318_));
 sky130_fd_sc_hd__nor2_1 _4839_ (.A(_1317_),
    .B(_1318_),
    .Y(_1319_));
 sky130_fd_sc_hd__inv_2 _4840_ (.A(_3327_),
    .Y(_1320_));
 sky130_fd_sc_hd__o22ai_1 _4841_ (.A1(_1196_),
    .A2(_3289_),
    .B1(_1320_),
    .B2(_3293_),
    .Y(_1321_));
 sky130_fd_sc_hd__a221oi_1 _4842_ (.A1(_3341_),
    .A2(_3281_),
    .B1(_3347_),
    .B2(_3285_),
    .C1(_1321_),
    .Y(_1322_));
 sky130_fd_sc_hd__and4_1 _4843_ (.A(_1311_),
    .B(_1316_),
    .C(_1319_),
    .D(_1322_),
    .X(_1323_));
 sky130_fd_sc_hd__nand2_1 _4844_ (.A(_3309_),
    .B(_0675_),
    .Y(_1324_));
 sky130_fd_sc_hd__nand2_1 _4845_ (.A(_3313_),
    .B(_0674_),
    .Y(_1325_));
 sky130_fd_sc_hd__nand2_1 _4846_ (.A(_1324_),
    .B(_1325_),
    .Y(_1326_));
 sky130_fd_sc_hd__a221oi_1 _4847_ (.A1(_2998_),
    .A2(_3303_),
    .B1(_3010_),
    .B2(_3307_),
    .C1(_1326_),
    .Y(_1327_));
 sky130_fd_sc_hd__nand2_1 _4848_ (.A(_3326_),
    .B(_3310_),
    .Y(_1328_));
 sky130_fd_sc_hd__nand2_1 _4849_ (.A(_3330_),
    .B(_3314_),
    .Y(_1329_));
 sky130_fd_sc_hd__nand2_1 _4850_ (.A(_1328_),
    .B(_1329_),
    .Y(_1330_));
 sky130_fd_sc_hd__a221oi_1 _4851_ (.A1(_3345_),
    .A2(_3321_),
    .B1(_3335_),
    .B2(_3324_),
    .C1(_1330_),
    .Y(_1331_));
 sky130_fd_sc_hd__inv_2 _4852_ (.A(\egd_top.BitStream_buffer.BS_buffer[109] ),
    .Y(_1332_));
 sky130_fd_sc_hd__nand2_1 _4853_ (.A(_3340_),
    .B(_3297_),
    .Y(_1333_));
 sky130_fd_sc_hd__nand2_1 _4854_ (.A(_3344_),
    .B(\egd_top.BitStream_buffer.BS_buffer[108] ),
    .Y(_1334_));
 sky130_fd_sc_hd__or2_1 _4855_ (.A(_1081_),
    .B(_3350_),
    .X(_1335_));
 sky130_fd_sc_hd__o2111a_1 _4856_ (.A1(_1332_),
    .A2(_3338_),
    .B1(_1333_),
    .C1(_1334_),
    .D1(_1335_),
    .X(_1336_));
 sky130_fd_sc_hd__nand2_1 _4857_ (.A(_3365_),
    .B(_3019_),
    .Y(_1337_));
 sky130_fd_sc_hd__o21ai_1 _4858_ (.A1(_3177_),
    .A2(_3363_),
    .B1(_1337_),
    .Y(_1338_));
 sky130_fd_sc_hd__a221oi_1 _4859_ (.A1(_3013_),
    .A2(_3356_),
    .B1(_3016_),
    .B2(_3360_),
    .C1(_1338_),
    .Y(_1339_));
 sky130_fd_sc_hd__and4_1 _4860_ (.A(_1327_),
    .B(_1331_),
    .C(_1336_),
    .D(_1339_),
    .X(_1340_));
 sky130_fd_sc_hd__and4_1 _4861_ (.A(_1298_),
    .B(_1309_),
    .C(_1323_),
    .D(_1340_),
    .X(_1341_));
 sky130_fd_sc_hd__nand2_1 _4862_ (.A(_0334_),
    .B(_0695_),
    .Y(_1342_));
 sky130_fd_sc_hd__nand2_1 _4863_ (.A(_0338_),
    .B(_0389_),
    .Y(_1343_));
 sky130_fd_sc_hd__nand2_1 _4864_ (.A(_1342_),
    .B(_1343_),
    .Y(_1344_));
 sky130_fd_sc_hd__a221oi_1 _4865_ (.A1(_0437_),
    .A2(_0328_),
    .B1(_0443_),
    .B2(_0332_),
    .C1(_1344_),
    .Y(_1345_));
 sky130_fd_sc_hd__inv_2 _4866_ (.A(\egd_top.BitStream_buffer.BS_buffer[43] ),
    .Y(_1346_));
 sky130_fd_sc_hd__o22ai_1 _4867_ (.A1(_1222_),
    .A2(_0345_),
    .B1(_1346_),
    .B2(_0349_),
    .Y(_1347_));
 sky130_fd_sc_hd__a22o_1 _4868_ (.A1(_0352_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[44] ),
    .B1(_0355_),
    .B2(_0380_),
    .X(_1348_));
 sky130_fd_sc_hd__nor2_1 _4869_ (.A(_1347_),
    .B(_1348_),
    .Y(_1349_));
 sky130_fd_sc_hd__nand2_1 _4870_ (.A(_0371_),
    .B(_0335_),
    .Y(_1350_));
 sky130_fd_sc_hd__o21ai_1 _4871_ (.A1(_0966_),
    .A2(_0369_),
    .B1(_1350_),
    .Y(_1351_));
 sky130_fd_sc_hd__a221oi_1 _4872_ (.A1(_0353_),
    .A2(_0362_),
    .B1(_0356_),
    .B2(_0366_),
    .C1(_1351_),
    .Y(_1352_));
 sky130_fd_sc_hd__nand2_1 _4873_ (.A(_0388_),
    .B(_0404_),
    .Y(_1353_));
 sky130_fd_sc_hd__o21ai_1 _4874_ (.A1(_0394_),
    .A2(_0386_),
    .B1(_1353_),
    .Y(_1354_));
 sky130_fd_sc_hd__a221oi_1 _4875_ (.A1(_0429_),
    .A2(_0379_),
    .B1(_0433_),
    .B2(_0383_),
    .C1(_1354_),
    .Y(_1355_));
 sky130_fd_sc_hd__and4_1 _4876_ (.A(_1345_),
    .B(_1349_),
    .C(_1352_),
    .D(_1355_),
    .X(_1356_));
 sky130_fd_sc_hd__nand2_1 _4877_ (.A(_0399_),
    .B(_0447_),
    .Y(_1357_));
 sky130_fd_sc_hd__nand2_1 _4878_ (.A(_0403_),
    .B(_0421_),
    .Y(_1358_));
 sky130_fd_sc_hd__or2_1 _4879_ (.A(_0848_),
    .B(_0408_),
    .X(_1359_));
 sky130_fd_sc_hd__o2111a_1 _4880_ (.A1(_0412_),
    .A2(_0397_),
    .B1(_1357_),
    .C1(_1358_),
    .D1(_1359_),
    .X(_1360_));
 sky130_fd_sc_hd__nand2_1 _4881_ (.A(_0416_),
    .B(_0461_),
    .Y(_1361_));
 sky130_fd_sc_hd__nand2_1 _4882_ (.A(_0420_),
    .B(_3107_),
    .Y(_1362_));
 sky130_fd_sc_hd__or2_1 _4883_ (.A(_0456_),
    .B(_0426_),
    .X(_1363_));
 sky130_fd_sc_hd__o2111a_1 _4884_ (.A1(_0614_),
    .A2(_0414_),
    .B1(_1361_),
    .C1(_1362_),
    .D1(_1363_),
    .X(_1364_));
 sky130_fd_sc_hd__nand2_1 _4885_ (.A(_0442_),
    .B(_0701_),
    .Y(_1365_));
 sky130_fd_sc_hd__o21ai_1 _4886_ (.A1(_0700_),
    .A2(_0440_),
    .B1(_1365_),
    .Y(_1366_));
 sky130_fd_sc_hd__a221oi_1 _4887_ (.A1(_0417_),
    .A2(_0432_),
    .B1(_0423_),
    .B2(_0436_),
    .C1(_1366_),
    .Y(_1367_));
 sky130_fd_sc_hd__nand2_1 _4888_ (.A(_0460_),
    .B(_3129_),
    .Y(_1368_));
 sky130_fd_sc_hd__o21ai_1 _4889_ (.A1(_3137_),
    .A2(_0458_),
    .B1(_1368_),
    .Y(_1369_));
 sky130_fd_sc_hd__a221oi_1 _4890_ (.A1(_3095_),
    .A2(_0450_),
    .B1(_3102_),
    .B2(_0454_),
    .C1(_1369_),
    .Y(_1370_));
 sky130_fd_sc_hd__and4_1 _4891_ (.A(_1360_),
    .B(_1364_),
    .C(_1367_),
    .D(_1370_),
    .X(_1371_));
 sky130_fd_sc_hd__and2_1 _4892_ (.A(_1356_),
    .B(_1371_),
    .X(_1372_));
 sky130_fd_sc_hd__inv_2 _4893_ (.A(\egd_top.BitStream_buffer.BS_buffer[30] ),
    .Y(_1373_));
 sky130_fd_sc_hd__nand2_1 _4894_ (.A(_0474_),
    .B(_0525_),
    .Y(_1374_));
 sky130_fd_sc_hd__a22o_1 _4895_ (.A1(_0478_),
    .A2(_0359_),
    .B1(_0481_),
    .B2(_0363_),
    .X(_1375_));
 sky130_fd_sc_hd__inv_2 _4896_ (.A(_1375_),
    .Y(_1376_));
 sky130_fd_sc_hd__o211a_1 _4897_ (.A1(_1373_),
    .A2(_0472_),
    .B1(_1374_),
    .C1(_1376_),
    .X(_1377_));
 sky130_fd_sc_hd__nand2_1 _4898_ (.A(_0498_),
    .B(_0475_),
    .Y(_1378_));
 sky130_fd_sc_hd__o21ai_1 _4899_ (.A1(_0468_),
    .A2(_0496_),
    .B1(_1378_),
    .Y(_1379_));
 sky130_fd_sc_hd__a221oi_1 _4900_ (.A1(_0509_),
    .A2(_0488_),
    .B1(_0503_),
    .B2(_0492_),
    .C1(_1379_),
    .Y(_1380_));
 sky130_fd_sc_hd__nand2_1 _4901_ (.A(_0508_),
    .B(_0535_),
    .Y(_1381_));
 sky130_fd_sc_hd__nand2_1 _4902_ (.A(_0512_),
    .B(_0479_),
    .Y(_1382_));
 sky130_fd_sc_hd__or2_1 _4903_ (.A(_0995_),
    .B(_0518_),
    .X(_1383_));
 sky130_fd_sc_hd__o2111a_1 _4904_ (.A1(_1249_),
    .A2(_0506_),
    .B1(_1381_),
    .C1(_1382_),
    .D1(_1383_),
    .X(_1384_));
 sky130_fd_sc_hd__nand2_1 _4905_ (.A(_0530_),
    .B(_0372_),
    .Y(_1385_));
 sky130_fd_sc_hd__nand2_1 _4906_ (.A(_0534_),
    .B(_0689_),
    .Y(_1386_));
 sky130_fd_sc_hd__nand2_1 _4907_ (.A(_1385_),
    .B(_1386_),
    .Y(_1387_));
 sky130_fd_sc_hd__a221oi_1 _4908_ (.A1(_0691_),
    .A2(_0524_),
    .B1(_0346_),
    .B2(_0528_),
    .C1(_1387_),
    .Y(_1388_));
 sky130_fd_sc_hd__and4_1 _4909_ (.A(_1377_),
    .B(_1380_),
    .C(_1384_),
    .D(_1388_),
    .X(_1389_));
 sky130_fd_sc_hd__nand2_1 _4910_ (.A(_0547_),
    .B(\egd_top.BitStream_buffer.BS_buffer[12] ),
    .Y(_1390_));
 sky130_fd_sc_hd__nand2_1 _4911_ (.A(_0551_),
    .B(\egd_top.BitStream_buffer.BS_buffer[10] ),
    .Y(_1391_));
 sky130_fd_sc_hd__or2_1 _4912_ (.A(_0596_),
    .B(_0556_),
    .X(_1392_));
 sky130_fd_sc_hd__o2111a_1 _4913_ (.A1(_0559_),
    .A2(_0545_),
    .B1(_1390_),
    .C1(_1391_),
    .D1(_1392_),
    .X(_1393_));
 sky130_fd_sc_hd__nand2_1 _4914_ (.A(_0563_),
    .B(\egd_top.BitStream_buffer.BS_buffer[16] ),
    .Y(_1394_));
 sky130_fd_sc_hd__nand2_1 _4915_ (.A(_0566_),
    .B(\egd_top.BitStream_buffer.BS_buffer[14] ),
    .Y(_1395_));
 sky130_fd_sc_hd__or2_1 _4916_ (.A(_0890_),
    .B(_0570_),
    .X(_1396_));
 sky130_fd_sc_hd__o2111a_1 _4917_ (.A1(_1150_),
    .A2(_0561_),
    .B1(_1394_),
    .C1(_1395_),
    .D1(_1396_),
    .X(_1397_));
 sky130_fd_sc_hd__or2_1 _4918_ (.A(_0568_),
    .B(_0584_),
    .X(_1398_));
 sky130_fd_sc_hd__o221a_1 _4919_ (.A1(_0745_),
    .A2(_0576_),
    .B1(_0554_),
    .B2(_0580_),
    .C1(_1398_),
    .X(_1399_));
 sky130_fd_sc_hd__o22ai_1 _4920_ (.A1(_0494_),
    .A2(_0595_),
    .B1(_0728_),
    .B2(_0598_),
    .Y(_1400_));
 sky130_fd_sc_hd__a221oi_1 _4921_ (.A1(_0513_),
    .A2(_0589_),
    .B1(_0515_),
    .B2(_0592_),
    .C1(_1400_),
    .Y(_1401_));
 sky130_fd_sc_hd__and4_1 _4922_ (.A(_1393_),
    .B(_1397_),
    .C(_1399_),
    .D(_1401_),
    .X(_1402_));
 sky130_fd_sc_hd__and3_1 _4923_ (.A(_1372_),
    .B(_1389_),
    .C(_1402_),
    .X(_1403_));
 sky130_fd_sc_hd__nand2_1 _4924_ (.A(_0606_),
    .B(_0548_),
    .Y(_1404_));
 sky130_fd_sc_hd__nand3_1 _4925_ (.A(_1341_),
    .B(_1403_),
    .C(_1404_),
    .Y(_1405_));
 sky130_fd_sc_hd__inv_2 _4926_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[9] ),
    .Y(_1406_));
 sky130_fd_sc_hd__a21oi_1 _4927_ (.A1(_1406_),
    .A2(_0898_),
    .B1(_2938_),
    .Y(_1407_));
 sky130_fd_sc_hd__o21a_1 _4928_ (.A1(_3056_),
    .A2(_1405_),
    .B1(_1407_),
    .X(_0291_));
 sky130_fd_sc_hd__inv_2 _4929_ (.A(\egd_top.BitStream_buffer.BS_buffer[80] ),
    .Y(_1408_));
 sky130_fd_sc_hd__o22ai_1 _4930_ (.A1(_1284_),
    .A2(_3084_),
    .B1(_1408_),
    .B2(_3092_),
    .Y(_1409_));
 sky130_fd_sc_hd__a221oi_1 _4931_ (.A1(_3247_),
    .A2(_3068_),
    .B1(_3259_),
    .B2(_3075_),
    .C1(_1409_),
    .Y(_1410_));
 sky130_fd_sc_hd__nand2_1 _4932_ (.A(_3114_),
    .B(_3076_),
    .Y(_1411_));
 sky130_fd_sc_hd__o21ai_1 _4933_ (.A1(_3120_),
    .A2(_3111_),
    .B1(_1411_),
    .Y(_1412_));
 sky130_fd_sc_hd__a221oi_1 _4934_ (.A1(_3085_),
    .A2(_3101_),
    .B1(_3057_),
    .B2(_3106_),
    .C1(_1412_),
    .Y(_1413_));
 sky130_fd_sc_hd__nand2_1 _4935_ (.A(_3128_),
    .B(_3069_),
    .Y(_1414_));
 sky130_fd_sc_hd__nand2_1 _4936_ (.A(_3133_),
    .B(_3156_),
    .Y(_1415_));
 sky130_fd_sc_hd__or2_1 _4937_ (.A(_0900_),
    .B(_3141_),
    .X(_1416_));
 sky130_fd_sc_hd__o2111a_1 _4938_ (.A1(_1159_),
    .A2(_3124_),
    .B1(_1414_),
    .C1(_1415_),
    .D1(_1416_),
    .X(_1417_));
 sky130_fd_sc_hd__nand2_1 _4939_ (.A(_3155_),
    .B(_0646_),
    .Y(_1418_));
 sky130_fd_sc_hd__nand2_1 _4940_ (.A(_3160_),
    .B(_3251_),
    .Y(_1419_));
 sky130_fd_sc_hd__nand2_1 _4941_ (.A(_1418_),
    .B(_1419_),
    .Y(_1420_));
 sky130_fd_sc_hd__a221oi_1 _4942_ (.A1(_3265_),
    .A2(_3148_),
    .B1(_3272_),
    .B2(_3152_),
    .C1(_1420_),
    .Y(_1421_));
 sky130_fd_sc_hd__and4_1 _4943_ (.A(_1410_),
    .B(_1413_),
    .C(_1417_),
    .D(_1421_),
    .X(_1422_));
 sky130_fd_sc_hd__o22ai_1 _4944_ (.A1(_3188_),
    .A2(_3176_),
    .B1(_3216_),
    .B2(_3179_),
    .Y(_1423_));
 sky130_fd_sc_hd__a221oi_1 _4945_ (.A1(_3047_),
    .A2(_3170_),
    .B1(_3050_),
    .B2(_3173_),
    .C1(_1423_),
    .Y(_1424_));
 sky130_fd_sc_hd__nand2_1 _4946_ (.A(_3192_),
    .B(_0577_),
    .Y(_1425_));
 sky130_fd_sc_hd__o21ai_1 _4947_ (.A1(_0574_),
    .A2(_3190_),
    .B1(_1425_),
    .Y(_1426_));
 sky130_fd_sc_hd__a221oi_1 _4948_ (.A1(_3053_),
    .A2(_3184_),
    .B1(_0607_),
    .B2(_3187_),
    .C1(_1426_),
    .Y(_1427_));
 sky130_fd_sc_hd__nand2_1 _4949_ (.A(_3206_),
    .B(_3031_),
    .Y(_1428_));
 sky130_fd_sc_hd__o21ai_1 _4950_ (.A1(_0780_),
    .A2(_3204_),
    .B1(_1428_),
    .Y(_1429_));
 sky130_fd_sc_hd__a221oi_2 _4951_ (.A1(_3034_),
    .A2(_3198_),
    .B1(_3037_),
    .B2(_3201_),
    .C1(_1429_),
    .Y(_1430_));
 sky130_fd_sc_hd__o22ai_1 _4952_ (.A1(_0582_),
    .A2(_3218_),
    .B1(_0753_),
    .B2(_3221_),
    .Y(_1431_));
 sky130_fd_sc_hd__a221oi_1 _4953_ (.A1(_0540_),
    .A2(_3212_),
    .B1(_0548_),
    .B2(_3215_),
    .C1(_1431_),
    .Y(_1432_));
 sky130_fd_sc_hd__and4_1 _4954_ (.A(_1424_),
    .B(_1427_),
    .C(_1430_),
    .D(_1432_),
    .X(_1433_));
 sky130_fd_sc_hd__o22ai_1 _4955_ (.A1(_0807_),
    .A2(_3238_),
    .B1(_0940_),
    .B2(_3241_),
    .Y(_1434_));
 sky130_fd_sc_hd__a221oi_1 _4956_ (.A1(_3322_),
    .A2(_3231_),
    .B1(_3331_),
    .B2(_3235_),
    .C1(_1434_),
    .Y(_1435_));
 sky130_fd_sc_hd__nand2_1 _4957_ (.A(_3246_),
    .B(_0653_),
    .Y(_1436_));
 sky130_fd_sc_hd__nand2_1 _4958_ (.A(_3250_),
    .B(_3225_),
    .Y(_1437_));
 sky130_fd_sc_hd__nand2_1 _4959_ (.A(_3254_),
    .B(_3275_),
    .Y(_1438_));
 sky130_fd_sc_hd__nand2_1 _4960_ (.A(_3258_),
    .B(_0804_),
    .Y(_1439_));
 sky130_fd_sc_hd__and4_1 _4961_ (.A(_1436_),
    .B(_1437_),
    .C(_1438_),
    .D(_1439_),
    .X(_1440_));
 sky130_fd_sc_hd__o22ai_1 _4962_ (.A1(_0794_),
    .A2(_3264_),
    .B1(_3287_),
    .B2(_3268_),
    .Y(_1441_));
 sky130_fd_sc_hd__a22o_1 _4963_ (.A1(_3271_),
    .A2(_3290_),
    .B1(_3274_),
    .B2(_3278_),
    .X(_1442_));
 sky130_fd_sc_hd__nor2_1 _4964_ (.A(_1441_),
    .B(_1442_),
    .Y(_1443_));
 sky130_fd_sc_hd__inv_2 _4965_ (.A(\egd_top.BitStream_buffer.BS_buffer[100] ),
    .Y(_1444_));
 sky130_fd_sc_hd__o22ai_1 _4966_ (.A1(_1320_),
    .A2(_3289_),
    .B1(_1444_),
    .B2(_3293_),
    .Y(_1445_));
 sky130_fd_sc_hd__a221oi_1 _4967_ (.A1(_3347_),
    .A2(_3281_),
    .B1(_3345_),
    .B2(_3285_),
    .C1(_1445_),
    .Y(_1446_));
 sky130_fd_sc_hd__and4_1 _4968_ (.A(_1435_),
    .B(_1440_),
    .C(_1443_),
    .D(_1446_),
    .X(_1447_));
 sky130_fd_sc_hd__nand2_1 _4969_ (.A(_3309_),
    .B(_2998_),
    .Y(_1448_));
 sky130_fd_sc_hd__nand2_1 _4970_ (.A(_3313_),
    .B(_0675_),
    .Y(_1449_));
 sky130_fd_sc_hd__nand2_1 _4971_ (.A(_1448_),
    .B(_1449_),
    .Y(_1450_));
 sky130_fd_sc_hd__a221oi_1 _4972_ (.A1(_3010_),
    .A2(_3303_),
    .B1(_3013_),
    .B2(_3307_),
    .C1(_1450_),
    .Y(_1451_));
 sky130_fd_sc_hd__nand2_1 _4973_ (.A(_3326_),
    .B(_3297_),
    .Y(_1452_));
 sky130_fd_sc_hd__nand2_1 _4974_ (.A(_3330_),
    .B(_3310_),
    .Y(_1453_));
 sky130_fd_sc_hd__nand2_1 _4975_ (.A(_1452_),
    .B(_1453_),
    .Y(_1454_));
 sky130_fd_sc_hd__a221oi_1 _4976_ (.A1(_3335_),
    .A2(_3321_),
    .B1(_3314_),
    .B2(_3324_),
    .C1(_1454_),
    .Y(_1455_));
 sky130_fd_sc_hd__inv_2 _4977_ (.A(\egd_top.BitStream_buffer.BS_buffer[110] ),
    .Y(_1456_));
 sky130_fd_sc_hd__nand2_1 _4978_ (.A(_3340_),
    .B(\egd_top.BitStream_buffer.BS_buffer[107] ),
    .Y(_1457_));
 sky130_fd_sc_hd__nand2_1 _4979_ (.A(_3344_),
    .B(\egd_top.BitStream_buffer.BS_buffer[109] ),
    .Y(_1458_));
 sky130_fd_sc_hd__or2_1 _4980_ (.A(_1208_),
    .B(_3350_),
    .X(_1459_));
 sky130_fd_sc_hd__o2111a_1 _4981_ (.A1(_1456_),
    .A2(_3338_),
    .B1(_1457_),
    .C1(_1458_),
    .D1(_1459_),
    .X(_1460_));
 sky130_fd_sc_hd__nand2_1 _4982_ (.A(_3365_),
    .B(_3022_),
    .Y(_1461_));
 sky130_fd_sc_hd__o21ai_1 _4983_ (.A1(_0628_),
    .A2(_3363_),
    .B1(_1461_),
    .Y(_1462_));
 sky130_fd_sc_hd__a221oi_2 _4984_ (.A1(_3016_),
    .A2(_3356_),
    .B1(_3019_),
    .B2(_3360_),
    .C1(_1462_),
    .Y(_1463_));
 sky130_fd_sc_hd__and4_1 _4985_ (.A(_1451_),
    .B(_1455_),
    .C(_1460_),
    .D(_1463_),
    .X(_1464_));
 sky130_fd_sc_hd__and4_1 _4986_ (.A(_1422_),
    .B(_1433_),
    .C(_1447_),
    .D(_1464_),
    .X(_1465_));
 sky130_fd_sc_hd__nand2_1 _4987_ (.A(_0334_),
    .B(_0437_),
    .Y(_1466_));
 sky130_fd_sc_hd__nand2_1 _4988_ (.A(_0338_),
    .B(_0695_),
    .Y(_1467_));
 sky130_fd_sc_hd__nand2_1 _4989_ (.A(_1466_),
    .B(_1467_),
    .Y(_1468_));
 sky130_fd_sc_hd__a221oi_1 _4990_ (.A1(_0443_),
    .A2(_0328_),
    .B1(_0429_),
    .B2(_0332_),
    .C1(_1468_),
    .Y(_1469_));
 sky130_fd_sc_hd__inv_2 _4991_ (.A(\egd_top.BitStream_buffer.BS_buffer[44] ),
    .Y(_1470_));
 sky130_fd_sc_hd__o22ai_1 _4992_ (.A1(_1346_),
    .A2(_0345_),
    .B1(_1470_),
    .B2(_0349_),
    .Y(_1471_));
 sky130_fd_sc_hd__a22o_1 _4993_ (.A1(_0352_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[45] ),
    .B1(_0355_),
    .B2(_0389_),
    .X(_1472_));
 sky130_fd_sc_hd__nor2_1 _4994_ (.A(_1471_),
    .B(_1472_),
    .Y(_1473_));
 sky130_fd_sc_hd__nand2_1 _4995_ (.A(_0371_),
    .B(_0323_),
    .Y(_1474_));
 sky130_fd_sc_hd__o21ai_1 _4996_ (.A1(_1095_),
    .A2(_0369_),
    .B1(_1474_),
    .Y(_1475_));
 sky130_fd_sc_hd__a221oi_1 _4997_ (.A1(_0356_),
    .A2(_0362_),
    .B1(_0339_),
    .B2(_0366_),
    .C1(_1475_),
    .Y(_1476_));
 sky130_fd_sc_hd__nand2_1 _4998_ (.A(_0388_),
    .B(_0703_),
    .Y(_1477_));
 sky130_fd_sc_hd__o21ai_1 _4999_ (.A1(_0700_),
    .A2(_0386_),
    .B1(_1477_),
    .Y(_1478_));
 sky130_fd_sc_hd__a221oi_1 _5000_ (.A1(_0433_),
    .A2(_0379_),
    .B1(_0404_),
    .B2(_0383_),
    .C1(_1478_),
    .Y(_1479_));
 sky130_fd_sc_hd__and4_1 _5001_ (.A(_1469_),
    .B(_1473_),
    .C(_1476_),
    .D(_1479_),
    .X(_1480_));
 sky130_fd_sc_hd__nand2_1 _5002_ (.A(_0399_),
    .B(_0451_),
    .Y(_1481_));
 sky130_fd_sc_hd__nand2_1 _5003_ (.A(_0403_),
    .B(_0411_),
    .Y(_1482_));
 sky130_fd_sc_hd__or2_1 _5004_ (.A(_0981_),
    .B(_0408_),
    .X(_1483_));
 sky130_fd_sc_hd__o2111a_1 _5005_ (.A1(_0708_),
    .A2(_0397_),
    .B1(_1481_),
    .C1(_1482_),
    .D1(_1483_),
    .X(_1484_));
 sky130_fd_sc_hd__nand2_1 _5006_ (.A(_0416_),
    .B(_0455_),
    .Y(_1485_));
 sky130_fd_sc_hd__nand2_1 _5007_ (.A(_0420_),
    .B(_3115_),
    .Y(_1486_));
 sky130_fd_sc_hd__or2_1 _5008_ (.A(_3108_),
    .B(_0426_),
    .X(_1487_));
 sky130_fd_sc_hd__o2111a_1 _5009_ (.A1(_0767_),
    .A2(_0414_),
    .B1(_1485_),
    .C1(_1486_),
    .D1(_1487_),
    .X(_1488_));
 sky130_fd_sc_hd__nand2_1 _5010_ (.A(_0442_),
    .B(_0417_),
    .Y(_1489_));
 sky130_fd_sc_hd__o21ai_1 _5011_ (.A1(_0406_),
    .A2(_0440_),
    .B1(_1489_),
    .Y(_1490_));
 sky130_fd_sc_hd__a221oi_1 _5012_ (.A1(_0423_),
    .A2(_0432_),
    .B1(_0421_),
    .B2(_0436_),
    .C1(_1490_),
    .Y(_1491_));
 sky130_fd_sc_hd__nand2_1 _5013_ (.A(_0460_),
    .B(_3136_),
    .Y(_1492_));
 sky130_fd_sc_hd__o21ai_1 _5014_ (.A1(_0620_),
    .A2(_0458_),
    .B1(_1492_),
    .Y(_1493_));
 sky130_fd_sc_hd__a221oi_1 _5015_ (.A1(_3102_),
    .A2(_0450_),
    .B1(_3129_),
    .B2(_0454_),
    .C1(_1493_),
    .Y(_1494_));
 sky130_fd_sc_hd__and4_1 _5016_ (.A(_1484_),
    .B(_1488_),
    .C(_1491_),
    .D(_1494_),
    .X(_1495_));
 sky130_fd_sc_hd__and2_1 _5017_ (.A(_1480_),
    .B(_1495_),
    .X(_1496_));
 sky130_fd_sc_hd__inv_2 _5018_ (.A(\egd_top.BitStream_buffer.BS_buffer[31] ),
    .Y(_1497_));
 sky130_fd_sc_hd__nand2_1 _5019_ (.A(_0474_),
    .B(_0359_),
    .Y(_1498_));
 sky130_fd_sc_hd__a22o_1 _5020_ (.A1(_0478_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[33] ),
    .B1(_0481_),
    .B2(_0689_),
    .X(_1499_));
 sky130_fd_sc_hd__inv_2 _5021_ (.A(_1499_),
    .Y(_1500_));
 sky130_fd_sc_hd__o211a_1 _5022_ (.A1(_1497_),
    .A2(_0472_),
    .B1(_1498_),
    .C1(_1500_),
    .X(_1501_));
 sky130_fd_sc_hd__nand2_1 _5023_ (.A(_0498_),
    .B(_0479_),
    .Y(_1502_));
 sky130_fd_sc_hd__o21ai_1 _5024_ (.A1(_0723_),
    .A2(_0496_),
    .B1(_1502_),
    .Y(_1503_));
 sky130_fd_sc_hd__a221oi_1 _5025_ (.A1(_0503_),
    .A2(_0488_),
    .B1(_0467_),
    .B2(_0492_),
    .C1(_1503_),
    .Y(_1504_));
 sky130_fd_sc_hd__nand2_1 _5026_ (.A(_0508_),
    .B(_0531_),
    .Y(_1505_));
 sky130_fd_sc_hd__nand2_1 _5027_ (.A(_0512_),
    .B(_0482_),
    .Y(_1506_));
 sky130_fd_sc_hd__or2_1 _5028_ (.A(_1123_),
    .B(_0518_),
    .X(_1507_));
 sky130_fd_sc_hd__o2111a_1 _5029_ (.A1(_1373_),
    .A2(_0506_),
    .B1(_1505_),
    .C1(_1506_),
    .D1(_1507_),
    .X(_1508_));
 sky130_fd_sc_hd__nand2_1 _5030_ (.A(_0530_),
    .B(_0691_),
    .Y(_1509_));
 sky130_fd_sc_hd__nand2_1 _5031_ (.A(_0534_),
    .B(_0372_),
    .Y(_1510_));
 sky130_fd_sc_hd__nand2_1 _5032_ (.A(_1509_),
    .B(_1510_),
    .Y(_1511_));
 sky130_fd_sc_hd__a221oi_1 _5033_ (.A1(_0346_),
    .A2(_0524_),
    .B1(_0353_),
    .B2(_0528_),
    .C1(_1511_),
    .Y(_1512_));
 sky130_fd_sc_hd__and4_1 _5034_ (.A(_1501_),
    .B(_1504_),
    .C(_1508_),
    .D(_1512_),
    .X(_1513_));
 sky130_fd_sc_hd__nand2_1 _5035_ (.A(_0547_),
    .B(\egd_top.BitStream_buffer.BS_buffer[13] ),
    .Y(_1514_));
 sky130_fd_sc_hd__nand2_1 _5036_ (.A(_0551_),
    .B(\egd_top.BitStream_buffer.BS_buffer[11] ),
    .Y(_1515_));
 sky130_fd_sc_hd__or2_1 _5037_ (.A(_0756_),
    .B(_0556_),
    .X(_1516_));
 sky130_fd_sc_hd__o2111a_1 _5038_ (.A1(_0593_),
    .A2(_0545_),
    .B1(_1514_),
    .C1(_1515_),
    .D1(_1516_),
    .X(_1517_));
 sky130_fd_sc_hd__nand2_1 _5039_ (.A(_0563_),
    .B(_0489_),
    .Y(_1518_));
 sky130_fd_sc_hd__nand2_1 _5040_ (.A(_0566_),
    .B(\egd_top.BitStream_buffer.BS_buffer[15] ),
    .Y(_1519_));
 sky130_fd_sc_hd__or2_1 _5041_ (.A(_1022_),
    .B(_0570_),
    .X(_1520_));
 sky130_fd_sc_hd__o2111a_1 _5042_ (.A1(_0494_),
    .A2(_0561_),
    .B1(_1518_),
    .C1(_1519_),
    .D1(_1520_),
    .X(_1521_));
 sky130_fd_sc_hd__or2_1 _5043_ (.A(_0750_),
    .B(_0584_),
    .X(_1522_));
 sky130_fd_sc_hd__o221a_1 _5044_ (.A1(_0568_),
    .A2(_0576_),
    .B1(_0745_),
    .B2(_0580_),
    .C1(_1522_),
    .X(_1523_));
 sky130_fd_sc_hd__o22ai_1 _5045_ (.A1(_0728_),
    .A2(_0595_),
    .B1(_0867_),
    .B2(_0598_),
    .Y(_1524_));
 sky130_fd_sc_hd__a221oi_1 _5046_ (.A1(_0515_),
    .A2(_0589_),
    .B1(_0509_),
    .B2(_0592_),
    .C1(_1524_),
    .Y(_1525_));
 sky130_fd_sc_hd__and4_1 _5047_ (.A(_1517_),
    .B(_1521_),
    .C(_1523_),
    .D(_1525_),
    .X(_1526_));
 sky130_fd_sc_hd__and3_1 _5048_ (.A(_1496_),
    .B(_1513_),
    .C(_1526_),
    .X(_1527_));
 sky130_fd_sc_hd__nand2_1 _5049_ (.A(_0606_),
    .B(\egd_top.BitStream_buffer.BS_buffer[7] ),
    .Y(_1528_));
 sky130_fd_sc_hd__nand3_1 _5050_ (.A(_1465_),
    .B(_1527_),
    .C(_1528_),
    .Y(_1529_));
 sky130_fd_sc_hd__inv_2 _5051_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[8] ),
    .Y(_1530_));
 sky130_fd_sc_hd__a21oi_1 _5052_ (.A1(_1530_),
    .A2(_0898_),
    .B1(_2938_),
    .Y(_1531_));
 sky130_fd_sc_hd__o21a_1 _5053_ (.A1(_3056_),
    .A2(_1529_),
    .B1(_1531_),
    .X(_0290_));
 sky130_fd_sc_hd__inv_2 _5054_ (.A(\egd_top.BitStream_buffer.BS_buffer[81] ),
    .Y(_1532_));
 sky130_fd_sc_hd__o22ai_1 _5055_ (.A1(_1408_),
    .A2(_3084_),
    .B1(_1532_),
    .B2(_3092_),
    .Y(_1533_));
 sky130_fd_sc_hd__a221oi_1 _5056_ (.A1(_3259_),
    .A2(_3068_),
    .B1(_3251_),
    .B2(_3075_),
    .C1(_1533_),
    .Y(_1534_));
 sky130_fd_sc_hd__nand2_1 _5057_ (.A(_3114_),
    .B(_3085_),
    .Y(_1535_));
 sky130_fd_sc_hd__o21ai_1 _5058_ (.A1(_3077_),
    .A2(_3111_),
    .B1(_1535_),
    .Y(_1536_));
 sky130_fd_sc_hd__a221oi_1 _5059_ (.A1(_3057_),
    .A2(_3101_),
    .B1(_3069_),
    .B2(_3106_),
    .C1(_1536_),
    .Y(_1537_));
 sky130_fd_sc_hd__nand2_1 _5060_ (.A(_3128_),
    .B(_3161_),
    .Y(_1538_));
 sky130_fd_sc_hd__nand2_1 _5061_ (.A(_3133_),
    .B(_3144_),
    .Y(_1539_));
 sky130_fd_sc_hd__or2_1 _5062_ (.A(_1031_),
    .B(_3141_),
    .X(_1540_));
 sky130_fd_sc_hd__o2111a_1 _5063_ (.A1(_1284_),
    .A2(_3124_),
    .B1(_1538_),
    .C1(_1539_),
    .D1(_1540_),
    .X(_1541_));
 sky130_fd_sc_hd__nand2_1 _5064_ (.A(_3155_),
    .B(_3265_),
    .Y(_1542_));
 sky130_fd_sc_hd__nand2_1 _5065_ (.A(_3160_),
    .B(_0646_),
    .Y(_1543_));
 sky130_fd_sc_hd__nand2_1 _5066_ (.A(_1542_),
    .B(_1543_),
    .Y(_1544_));
 sky130_fd_sc_hd__a221oi_1 _5067_ (.A1(_3272_),
    .A2(_3148_),
    .B1(_3275_),
    .B2(_3152_),
    .C1(_1544_),
    .Y(_1545_));
 sky130_fd_sc_hd__and4_1 _5068_ (.A(_1534_),
    .B(_1537_),
    .C(_1541_),
    .D(_1545_),
    .X(_1546_));
 sky130_fd_sc_hd__o22ai_1 _5069_ (.A1(_3216_),
    .A2(_3176_),
    .B1(_3219_),
    .B2(_3179_),
    .Y(_1547_));
 sky130_fd_sc_hd__a221oi_1 _5070_ (.A1(_3050_),
    .A2(_3170_),
    .B1(_3053_),
    .B2(_3173_),
    .C1(_1547_),
    .Y(_1548_));
 sky130_fd_sc_hd__nand2_1 _5071_ (.A(_3192_),
    .B(_0573_),
    .Y(_1549_));
 sky130_fd_sc_hd__o21ai_1 _5072_ (.A1(_0582_),
    .A2(_3190_),
    .B1(_1549_),
    .Y(_1550_));
 sky130_fd_sc_hd__a221oi_1 _5073_ (.A1(_0607_),
    .A2(_3184_),
    .B1(_0577_),
    .B2(_3187_),
    .C1(_1550_),
    .Y(_1551_));
 sky130_fd_sc_hd__nand2_1 _5074_ (.A(_3206_),
    .B(_3034_),
    .Y(_1552_));
 sky130_fd_sc_hd__o21ai_1 _5075_ (.A1(_0916_),
    .A2(_3204_),
    .B1(_1552_),
    .Y(_1553_));
 sky130_fd_sc_hd__a221oi_1 _5076_ (.A1(_3037_),
    .A2(_3198_),
    .B1(_3040_),
    .B2(_3201_),
    .C1(_1553_),
    .Y(_1554_));
 sky130_fd_sc_hd__o22ai_1 _5077_ (.A1(_0753_),
    .A2(_3218_),
    .B1(_0541_),
    .B2(_3221_),
    .Y(_1555_));
 sky130_fd_sc_hd__a221oi_1 _5078_ (.A1(_0548_),
    .A2(_3212_),
    .B1(\egd_top.BitStream_buffer.BS_buffer[7] ),
    .B2(_3215_),
    .C1(_1555_),
    .Y(_1556_));
 sky130_fd_sc_hd__and4_1 _5079_ (.A(_1548_),
    .B(_1551_),
    .C(_1554_),
    .D(_1556_),
    .X(_1557_));
 sky130_fd_sc_hd__o22ai_1 _5080_ (.A1(_0940_),
    .A2(_3238_),
    .B1(_1069_),
    .B2(_3241_),
    .Y(_1558_));
 sky130_fd_sc_hd__a221oi_1 _5081_ (.A1(_3331_),
    .A2(_3231_),
    .B1(_3327_),
    .B2(_3235_),
    .C1(_1558_),
    .Y(_1559_));
 sky130_fd_sc_hd__nand2_1 _5082_ (.A(_3246_),
    .B(_0804_),
    .Y(_1560_));
 sky130_fd_sc_hd__nand2_1 _5083_ (.A(_3250_),
    .B(_3232_),
    .Y(_1561_));
 sky130_fd_sc_hd__nand2_1 _5084_ (.A(_3254_),
    .B(_0653_),
    .Y(_1562_));
 sky130_fd_sc_hd__nand2_1 _5085_ (.A(_3258_),
    .B(_3225_),
    .Y(_1563_));
 sky130_fd_sc_hd__and4_1 _5086_ (.A(_1560_),
    .B(_1561_),
    .C(_1562_),
    .D(_1563_),
    .X(_1564_));
 sky130_fd_sc_hd__o22ai_1 _5087_ (.A1(_3287_),
    .A2(_3264_),
    .B1(_3291_),
    .B2(_3268_),
    .Y(_1565_));
 sky130_fd_sc_hd__a22o_1 _5088_ (.A1(_3271_),
    .A2(_3278_),
    .B1(_3274_),
    .B2(_3282_),
    .X(_1566_));
 sky130_fd_sc_hd__nor2_1 _5089_ (.A(_1565_),
    .B(_1566_),
    .Y(_1567_));
 sky130_fd_sc_hd__o22ai_1 _5090_ (.A1(_1444_),
    .A2(_3289_),
    .B1(_3348_),
    .B2(_3293_),
    .Y(_1568_));
 sky130_fd_sc_hd__a221oi_1 _5091_ (.A1(_3345_),
    .A2(_3281_),
    .B1(_3335_),
    .B2(_3285_),
    .C1(_1568_),
    .Y(_1569_));
 sky130_fd_sc_hd__and4_1 _5092_ (.A(_1559_),
    .B(_1564_),
    .C(_1567_),
    .D(_1569_),
    .X(_1570_));
 sky130_fd_sc_hd__nand2_1 _5093_ (.A(_3309_),
    .B(_3010_),
    .Y(_1571_));
 sky130_fd_sc_hd__nand2_1 _5094_ (.A(_3313_),
    .B(_2998_),
    .Y(_1572_));
 sky130_fd_sc_hd__nand2_1 _5095_ (.A(_1571_),
    .B(_1572_),
    .Y(_1573_));
 sky130_fd_sc_hd__a221oi_1 _5096_ (.A1(_3013_),
    .A2(_3303_),
    .B1(_3016_),
    .B2(_3307_),
    .C1(_1573_),
    .Y(_1574_));
 sky130_fd_sc_hd__nand2_1 _5097_ (.A(_3326_),
    .B(_3304_),
    .Y(_1575_));
 sky130_fd_sc_hd__nand2_1 _5098_ (.A(_3330_),
    .B(_3297_),
    .Y(_1576_));
 sky130_fd_sc_hd__nand2_1 _5099_ (.A(_1575_),
    .B(_1576_),
    .Y(_1577_));
 sky130_fd_sc_hd__a221oi_1 _5100_ (.A1(_3314_),
    .A2(_3321_),
    .B1(_3310_),
    .B2(_3324_),
    .C1(_1577_),
    .Y(_1578_));
 sky130_fd_sc_hd__nand2_1 _5101_ (.A(_3340_),
    .B(\egd_top.BitStream_buffer.BS_buffer[108] ),
    .Y(_1579_));
 sky130_fd_sc_hd__nand2_1 _5102_ (.A(_3344_),
    .B(_0674_),
    .Y(_1580_));
 sky130_fd_sc_hd__or2_1 _5103_ (.A(_1332_),
    .B(_3350_),
    .X(_1581_));
 sky130_fd_sc_hd__o2111a_1 _5104_ (.A1(_3361_),
    .A2(_3338_),
    .B1(_1579_),
    .C1(_1580_),
    .D1(_1581_),
    .X(_1582_));
 sky130_fd_sc_hd__nand2_1 _5105_ (.A(_3365_),
    .B(_3025_),
    .Y(_1583_));
 sky130_fd_sc_hd__o21ai_1 _5106_ (.A1(_0780_),
    .A2(_3363_),
    .B1(_1583_),
    .Y(_1584_));
 sky130_fd_sc_hd__a221oi_1 _5107_ (.A1(_3019_),
    .A2(_3356_),
    .B1(_3022_),
    .B2(_3360_),
    .C1(_1584_),
    .Y(_1585_));
 sky130_fd_sc_hd__and4_1 _5108_ (.A(_1574_),
    .B(_1578_),
    .C(_1582_),
    .D(_1585_),
    .X(_1586_));
 sky130_fd_sc_hd__and4_1 _5109_ (.A(_1546_),
    .B(_1557_),
    .C(_1570_),
    .D(_1586_),
    .X(_1587_));
 sky130_fd_sc_hd__nand2_1 _5110_ (.A(_0334_),
    .B(_0443_),
    .Y(_1588_));
 sky130_fd_sc_hd__nand2_1 _5111_ (.A(_0338_),
    .B(_0437_),
    .Y(_1589_));
 sky130_fd_sc_hd__nand2_1 _5112_ (.A(_1588_),
    .B(_1589_),
    .Y(_1590_));
 sky130_fd_sc_hd__a221oi_1 _5113_ (.A1(_0429_),
    .A2(_0328_),
    .B1(_0433_),
    .B2(_0332_),
    .C1(_1590_),
    .Y(_1591_));
 sky130_fd_sc_hd__inv_2 _5114_ (.A(\egd_top.BitStream_buffer.BS_buffer[45] ),
    .Y(_1592_));
 sky130_fd_sc_hd__o22ai_1 _5115_ (.A1(_1470_),
    .A2(_0345_),
    .B1(_1592_),
    .B2(_0349_),
    .Y(_1593_));
 sky130_fd_sc_hd__a22o_1 _5116_ (.A1(_0352_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[46] ),
    .B1(_0355_),
    .B2(_0695_),
    .X(_1594_));
 sky130_fd_sc_hd__nor2_1 _5117_ (.A(_1593_),
    .B(_1594_),
    .Y(_1595_));
 sky130_fd_sc_hd__nand2_1 _5118_ (.A(_0371_),
    .B(_0329_),
    .Y(_1596_));
 sky130_fd_sc_hd__o21ai_1 _5119_ (.A1(_1222_),
    .A2(_0369_),
    .B1(_1596_),
    .Y(_1597_));
 sky130_fd_sc_hd__a221oi_1 _5120_ (.A1(_0339_),
    .A2(_0362_),
    .B1(_0335_),
    .B2(_0366_),
    .C1(_1597_),
    .Y(_1598_));
 sky130_fd_sc_hd__nand2_1 _5121_ (.A(_0388_),
    .B(_0400_),
    .Y(_1599_));
 sky130_fd_sc_hd__o21ai_1 _5122_ (.A1(_0406_),
    .A2(_0386_),
    .B1(_1599_),
    .Y(_1600_));
 sky130_fd_sc_hd__a221oi_1 _5123_ (.A1(_0404_),
    .A2(_0379_),
    .B1(_0703_),
    .B2(_0383_),
    .C1(_1600_),
    .Y(_1601_));
 sky130_fd_sc_hd__and4_1 _5124_ (.A(_1591_),
    .B(_1595_),
    .C(_1598_),
    .D(_1601_),
    .X(_1602_));
 sky130_fd_sc_hd__nand2_1 _5125_ (.A(_0399_),
    .B(_0461_),
    .Y(_1603_));
 sky130_fd_sc_hd__nand2_1 _5126_ (.A(_0403_),
    .B(_0447_),
    .Y(_1604_));
 sky130_fd_sc_hd__or2_1 _5127_ (.A(_0456_),
    .B(_0408_),
    .X(_1605_));
 sky130_fd_sc_hd__o2111a_1 _5128_ (.A1(_0848_),
    .A2(_0397_),
    .B1(_1603_),
    .C1(_1604_),
    .D1(_1605_),
    .X(_1606_));
 sky130_fd_sc_hd__nand2_1 _5129_ (.A(_0416_),
    .B(_3107_),
    .Y(_1607_));
 sky130_fd_sc_hd__nand2_1 _5130_ (.A(_0420_),
    .B(_3095_),
    .Y(_1608_));
 sky130_fd_sc_hd__or2_1 _5131_ (.A(_0614_),
    .B(_0426_),
    .X(_1609_));
 sky130_fd_sc_hd__o2111a_1 _5132_ (.A1(_0903_),
    .A2(_0414_),
    .B1(_1607_),
    .C1(_1608_),
    .D1(_1609_),
    .X(_1610_));
 sky130_fd_sc_hd__nand2_1 _5133_ (.A(_0442_),
    .B(_0423_),
    .Y(_1611_));
 sky130_fd_sc_hd__o21ai_1 _5134_ (.A1(_0705_),
    .A2(_0440_),
    .B1(_1611_),
    .Y(_1612_));
 sky130_fd_sc_hd__a221oi_1 _5135_ (.A1(_0421_),
    .A2(_0432_),
    .B1(_0411_),
    .B2(_0436_),
    .C1(_1612_),
    .Y(_1613_));
 sky130_fd_sc_hd__nand2_1 _5136_ (.A(_0460_),
    .B(_3134_),
    .Y(_1614_));
 sky130_fd_sc_hd__o21ai_1 _5137_ (.A1(_3120_),
    .A2(_0458_),
    .B1(_1614_),
    .Y(_1615_));
 sky130_fd_sc_hd__a221oi_1 _5138_ (.A1(_3129_),
    .A2(_0450_),
    .B1(_3136_),
    .B2(_0454_),
    .C1(_1615_),
    .Y(_1616_));
 sky130_fd_sc_hd__and4_1 _5139_ (.A(_1606_),
    .B(_1610_),
    .C(_1613_),
    .D(_1616_),
    .X(_1617_));
 sky130_fd_sc_hd__and2_1 _5140_ (.A(_1602_),
    .B(_1617_),
    .X(_1618_));
 sky130_fd_sc_hd__inv_2 _5141_ (.A(\egd_top.BitStream_buffer.BS_buffer[32] ),
    .Y(_1619_));
 sky130_fd_sc_hd__nand2_1 _5142_ (.A(_0474_),
    .B(_0363_),
    .Y(_1620_));
 sky130_fd_sc_hd__a22o_1 _5143_ (.A1(_0478_),
    .A2(_0689_),
    .B1(_0481_),
    .B2(_0372_),
    .X(_1621_));
 sky130_fd_sc_hd__inv_2 _5144_ (.A(_1621_),
    .Y(_1622_));
 sky130_fd_sc_hd__o211a_1 _5145_ (.A1(_1619_),
    .A2(_0472_),
    .B1(_1620_),
    .C1(_1622_),
    .X(_1623_));
 sky130_fd_sc_hd__nand2_1 _5146_ (.A(_0498_),
    .B(_0482_),
    .Y(_1624_));
 sky130_fd_sc_hd__o21ai_1 _5147_ (.A1(_0862_),
    .A2(_0496_),
    .B1(_1624_),
    .Y(_1625_));
 sky130_fd_sc_hd__a221oi_1 _5148_ (.A1(_0467_),
    .A2(_0488_),
    .B1(_0475_),
    .B2(_0492_),
    .C1(_1625_),
    .Y(_1626_));
 sky130_fd_sc_hd__nand2_1 _5149_ (.A(_0508_),
    .B(_0521_),
    .Y(_1627_));
 sky130_fd_sc_hd__nand2_1 _5150_ (.A(_0512_),
    .B(_0535_),
    .Y(_1628_));
 sky130_fd_sc_hd__or2_1 _5151_ (.A(_1249_),
    .B(_0518_),
    .X(_1629_));
 sky130_fd_sc_hd__o2111a_1 _5152_ (.A1(_1497_),
    .A2(_0506_),
    .B1(_1627_),
    .C1(_1628_),
    .D1(_1629_),
    .X(_1630_));
 sky130_fd_sc_hd__nand2_1 _5153_ (.A(_0530_),
    .B(_0346_),
    .Y(_1631_));
 sky130_fd_sc_hd__nand2_1 _5154_ (.A(_0534_),
    .B(_0691_),
    .Y(_1632_));
 sky130_fd_sc_hd__nand2_1 _5155_ (.A(_1631_),
    .B(_1632_),
    .Y(_1633_));
 sky130_fd_sc_hd__a221oi_1 _5156_ (.A1(_0353_),
    .A2(_0524_),
    .B1(_0356_),
    .B2(_0528_),
    .C1(_1633_),
    .Y(_1634_));
 sky130_fd_sc_hd__and4_1 _5157_ (.A(_1623_),
    .B(_1626_),
    .C(_1630_),
    .D(_1634_),
    .X(_1635_));
 sky130_fd_sc_hd__nand2_1 _5158_ (.A(_0547_),
    .B(\egd_top.BitStream_buffer.BS_buffer[14] ),
    .Y(_1636_));
 sky130_fd_sc_hd__nand2_1 _5159_ (.A(_0551_),
    .B(\egd_top.BitStream_buffer.BS_buffer[12] ),
    .Y(_1637_));
 sky130_fd_sc_hd__or2_1 _5160_ (.A(_0890_),
    .B(_0556_),
    .X(_1638_));
 sky130_fd_sc_hd__o2111a_1 _5161_ (.A1(_0596_),
    .A2(_0545_),
    .B1(_1636_),
    .C1(_1637_),
    .D1(_1638_),
    .X(_1639_));
 sky130_fd_sc_hd__nand2_1 _5162_ (.A(_0563_),
    .B(_0493_),
    .Y(_1640_));
 sky130_fd_sc_hd__nand2_1 _5163_ (.A(_0566_),
    .B(\egd_top.BitStream_buffer.BS_buffer[16] ),
    .Y(_1641_));
 sky130_fd_sc_hd__or2_1 _5164_ (.A(_1150_),
    .B(_0570_),
    .X(_1642_));
 sky130_fd_sc_hd__o2111a_1 _5165_ (.A1(_0728_),
    .A2(_0561_),
    .B1(_1640_),
    .C1(_1641_),
    .D1(_1642_),
    .X(_1643_));
 sky130_fd_sc_hd__or2_1 _5166_ (.A(_0559_),
    .B(_0584_),
    .X(_1644_));
 sky130_fd_sc_hd__o221a_1 _5167_ (.A1(_0750_),
    .A2(_0576_),
    .B1(_0568_),
    .B2(_0580_),
    .C1(_1644_),
    .X(_1645_));
 sky130_fd_sc_hd__o22ai_1 _5168_ (.A1(_0867_),
    .A2(_0595_),
    .B1(_0516_),
    .B2(_0598_),
    .Y(_1646_));
 sky130_fd_sc_hd__a221oi_1 _5169_ (.A1(_0509_),
    .A2(_0589_),
    .B1(_0503_),
    .B2(_0592_),
    .C1(_1646_),
    .Y(_1647_));
 sky130_fd_sc_hd__and4_1 _5170_ (.A(_1639_),
    .B(_1643_),
    .C(_1645_),
    .D(_1647_),
    .X(_1648_));
 sky130_fd_sc_hd__and3_1 _5171_ (.A(_1618_),
    .B(_1635_),
    .C(_1648_),
    .X(_1649_));
 sky130_fd_sc_hd__nand2_1 _5172_ (.A(_0606_),
    .B(\egd_top.BitStream_buffer.BS_buffer[8] ),
    .Y(_1650_));
 sky130_fd_sc_hd__nand3_1 _5173_ (.A(_1587_),
    .B(_1649_),
    .C(_1650_),
    .Y(_1651_));
 sky130_fd_sc_hd__inv_2 _5174_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[7] ),
    .Y(_1652_));
 sky130_fd_sc_hd__a21oi_1 _5175_ (.A1(_1652_),
    .A2(_0898_),
    .B1(_2938_),
    .Y(_1653_));
 sky130_fd_sc_hd__o21a_1 _5176_ (.A1(_3056_),
    .A2(_1651_),
    .B1(_1653_),
    .X(_0289_));
 sky130_fd_sc_hd__inv_2 _5177_ (.A(\egd_top.BitStream_buffer.BS_buffer[82] ),
    .Y(_1654_));
 sky130_fd_sc_hd__o22ai_1 _5178_ (.A1(_1532_),
    .A2(_3084_),
    .B1(_1654_),
    .B2(_3092_),
    .Y(_1655_));
 sky130_fd_sc_hd__a221oi_1 _5179_ (.A1(_3251_),
    .A2(_3068_),
    .B1(_0646_),
    .B2(_3075_),
    .C1(_1655_),
    .Y(_1656_));
 sky130_fd_sc_hd__nand2_1 _5180_ (.A(_3114_),
    .B(_3057_),
    .Y(_1657_));
 sky130_fd_sc_hd__o21ai_1 _5181_ (.A1(_3086_),
    .A2(_3111_),
    .B1(_1657_),
    .Y(_1658_));
 sky130_fd_sc_hd__a221oi_1 _5182_ (.A1(_3069_),
    .A2(_3101_),
    .B1(_3161_),
    .B2(_3106_),
    .C1(_1658_),
    .Y(_1659_));
 sky130_fd_sc_hd__nand2_1 _5183_ (.A(_3128_),
    .B(_3156_),
    .Y(_1660_));
 sky130_fd_sc_hd__nand2_1 _5184_ (.A(_3133_),
    .B(_3149_),
    .Y(_1661_));
 sky130_fd_sc_hd__or2_1 _5185_ (.A(_1159_),
    .B(_3141_),
    .X(_1662_));
 sky130_fd_sc_hd__o2111a_1 _5186_ (.A1(_1408_),
    .A2(_3124_),
    .B1(_1660_),
    .C1(_1661_),
    .D1(_1662_),
    .X(_1663_));
 sky130_fd_sc_hd__nand2_1 _5187_ (.A(_3155_),
    .B(_3272_),
    .Y(_1664_));
 sky130_fd_sc_hd__nand2_1 _5188_ (.A(_3160_),
    .B(_3265_),
    .Y(_1665_));
 sky130_fd_sc_hd__nand2_1 _5189_ (.A(_1664_),
    .B(_1665_),
    .Y(_1666_));
 sky130_fd_sc_hd__a221oi_2 _5190_ (.A1(_3275_),
    .A2(_3148_),
    .B1(_0653_),
    .B2(_3152_),
    .C1(_1666_),
    .Y(_1667_));
 sky130_fd_sc_hd__and4_1 _5191_ (.A(_1656_),
    .B(_1659_),
    .C(_1663_),
    .D(_1667_),
    .X(_1668_));
 sky130_fd_sc_hd__o22ai_1 _5192_ (.A1(_3219_),
    .A2(_3176_),
    .B1(_0638_),
    .B2(_3179_),
    .Y(_1669_));
 sky130_fd_sc_hd__a221oi_1 _5193_ (.A1(_3053_),
    .A2(_3170_),
    .B1(_0607_),
    .B2(_3173_),
    .C1(_1669_),
    .Y(_1670_));
 sky130_fd_sc_hd__nand2_1 _5194_ (.A(_3192_),
    .B(_0581_),
    .Y(_1671_));
 sky130_fd_sc_hd__o21ai_1 _5195_ (.A1(_0753_),
    .A2(_3190_),
    .B1(_1671_),
    .Y(_1672_));
 sky130_fd_sc_hd__a221oi_1 _5196_ (.A1(_0577_),
    .A2(_3184_),
    .B1(_0573_),
    .B2(_3187_),
    .C1(_1672_),
    .Y(_1673_));
 sky130_fd_sc_hd__nand2_1 _5197_ (.A(_3206_),
    .B(_3037_),
    .Y(_1674_));
 sky130_fd_sc_hd__o21ai_1 _5198_ (.A1(_1047_),
    .A2(_3204_),
    .B1(_1674_),
    .Y(_1675_));
 sky130_fd_sc_hd__a221oi_1 _5199_ (.A1(_3040_),
    .A2(_3198_),
    .B1(_3044_),
    .B2(_3201_),
    .C1(_1675_),
    .Y(_1676_));
 sky130_fd_sc_hd__o22ai_1 _5200_ (.A1(_0541_),
    .A2(_3218_),
    .B1(_0742_),
    .B2(_3221_),
    .Y(_1677_));
 sky130_fd_sc_hd__a221oi_1 _5201_ (.A1(\egd_top.BitStream_buffer.BS_buffer[7] ),
    .A2(_3212_),
    .B1(\egd_top.BitStream_buffer.BS_buffer[8] ),
    .B2(_3215_),
    .C1(_1677_),
    .Y(_1678_));
 sky130_fd_sc_hd__and4_1 _5202_ (.A(_1670_),
    .B(_1673_),
    .C(_1676_),
    .D(_1678_),
    .X(_1679_));
 sky130_fd_sc_hd__o22ai_1 _5203_ (.A1(_1069_),
    .A2(_3238_),
    .B1(_1196_),
    .B2(_3241_),
    .Y(_1680_));
 sky130_fd_sc_hd__a221oi_1 _5204_ (.A1(_3327_),
    .A2(_3231_),
    .B1(_3341_),
    .B2(_3235_),
    .C1(_1680_),
    .Y(_1681_));
 sky130_fd_sc_hd__nand2_1 _5205_ (.A(_3246_),
    .B(_3225_),
    .Y(_1682_));
 sky130_fd_sc_hd__nand2_1 _5206_ (.A(_3250_),
    .B(_3286_),
    .Y(_1683_));
 sky130_fd_sc_hd__nand2_1 _5207_ (.A(_3254_),
    .B(_0804_),
    .Y(_1684_));
 sky130_fd_sc_hd__nand2_1 _5208_ (.A(_3258_),
    .B(_3232_),
    .Y(_1685_));
 sky130_fd_sc_hd__and4_1 _5209_ (.A(_1682_),
    .B(_1683_),
    .C(_1684_),
    .D(_1685_),
    .X(_1686_));
 sky130_fd_sc_hd__o22ai_1 _5210_ (.A1(_3291_),
    .A2(_3264_),
    .B1(_0656_),
    .B2(_3268_),
    .Y(_1687_));
 sky130_fd_sc_hd__a22o_1 _5211_ (.A1(_3271_),
    .A2(_3282_),
    .B1(_3274_),
    .B2(_3318_),
    .X(_1688_));
 sky130_fd_sc_hd__nor2_1 _5212_ (.A(_1687_),
    .B(_1688_),
    .Y(_1689_));
 sky130_fd_sc_hd__o22ai_1 _5213_ (.A1(_3348_),
    .A2(_3289_),
    .B1(_0671_),
    .B2(_3293_),
    .Y(_1690_));
 sky130_fd_sc_hd__a221oi_2 _5214_ (.A1(_3335_),
    .A2(_3281_),
    .B1(_3314_),
    .B2(_3285_),
    .C1(_1690_),
    .Y(_1691_));
 sky130_fd_sc_hd__and4_1 _5215_ (.A(_1681_),
    .B(_1686_),
    .C(_1689_),
    .D(_1691_),
    .X(_1692_));
 sky130_fd_sc_hd__nand2_1 _5216_ (.A(_3309_),
    .B(_3013_),
    .Y(_1693_));
 sky130_fd_sc_hd__nand2_1 _5217_ (.A(_3313_),
    .B(_3010_),
    .Y(_1694_));
 sky130_fd_sc_hd__nand2_1 _5218_ (.A(_1693_),
    .B(_1694_),
    .Y(_1695_));
 sky130_fd_sc_hd__a221oi_1 _5219_ (.A1(_3016_),
    .A2(_3303_),
    .B1(_3019_),
    .B2(_3307_),
    .C1(_1695_),
    .Y(_1696_));
 sky130_fd_sc_hd__nand2_1 _5220_ (.A(_3326_),
    .B(_3353_),
    .Y(_1697_));
 sky130_fd_sc_hd__nand2_1 _5221_ (.A(_3330_),
    .B(_3304_),
    .Y(_1698_));
 sky130_fd_sc_hd__nand2_1 _5222_ (.A(_1697_),
    .B(_1698_),
    .Y(_1699_));
 sky130_fd_sc_hd__a221oi_1 _5223_ (.A1(_3310_),
    .A2(_3321_),
    .B1(_3297_),
    .B2(_3324_),
    .C1(_1699_),
    .Y(_1700_));
 sky130_fd_sc_hd__nand2_1 _5224_ (.A(_3340_),
    .B(\egd_top.BitStream_buffer.BS_buffer[109] ),
    .Y(_1701_));
 sky130_fd_sc_hd__nand2_1 _5225_ (.A(_3344_),
    .B(_0675_),
    .Y(_1702_));
 sky130_fd_sc_hd__or2_1 _5226_ (.A(_1456_),
    .B(_3350_),
    .X(_1703_));
 sky130_fd_sc_hd__o2111a_1 _5227_ (.A1(_3202_),
    .A2(_3338_),
    .B1(_1701_),
    .C1(_1702_),
    .D1(_1703_),
    .X(_1704_));
 sky130_fd_sc_hd__nand2_1 _5228_ (.A(_3365_),
    .B(_3028_),
    .Y(_1705_));
 sky130_fd_sc_hd__o21ai_1 _5229_ (.A1(_0916_),
    .A2(_3363_),
    .B1(_1705_),
    .Y(_1706_));
 sky130_fd_sc_hd__a221oi_1 _5230_ (.A1(_3022_),
    .A2(_3356_),
    .B1(_3025_),
    .B2(_3360_),
    .C1(_1706_),
    .Y(_1707_));
 sky130_fd_sc_hd__and4_1 _5231_ (.A(_1696_),
    .B(_1700_),
    .C(_1704_),
    .D(_1707_),
    .X(_1708_));
 sky130_fd_sc_hd__and4_1 _5232_ (.A(_1668_),
    .B(_1679_),
    .C(_1692_),
    .D(_1708_),
    .X(_1709_));
 sky130_fd_sc_hd__nand2_1 _5233_ (.A(_0334_),
    .B(_0429_),
    .Y(_1710_));
 sky130_fd_sc_hd__nand2_1 _5234_ (.A(_0338_),
    .B(_0443_),
    .Y(_1711_));
 sky130_fd_sc_hd__nand2_1 _5235_ (.A(_1710_),
    .B(_1711_),
    .Y(_1712_));
 sky130_fd_sc_hd__a221oi_1 _5236_ (.A1(_0433_),
    .A2(_0328_),
    .B1(_0404_),
    .B2(_0332_),
    .C1(_1712_),
    .Y(_1713_));
 sky130_fd_sc_hd__inv_2 _5237_ (.A(\egd_top.BitStream_buffer.BS_buffer[46] ),
    .Y(_1714_));
 sky130_fd_sc_hd__o22ai_1 _5238_ (.A1(_1592_),
    .A2(_0345_),
    .B1(_1714_),
    .B2(_0349_),
    .Y(_1715_));
 sky130_fd_sc_hd__a22o_1 _5239_ (.A1(_0352_),
    .A2(_0695_),
    .B1(_0355_),
    .B2(_0437_),
    .X(_1716_));
 sky130_fd_sc_hd__nor2_1 _5240_ (.A(_1715_),
    .B(_1716_),
    .Y(_1717_));
 sky130_fd_sc_hd__nand2_1 _5241_ (.A(_0371_),
    .B(_0376_),
    .Y(_1718_));
 sky130_fd_sc_hd__o21ai_1 _5242_ (.A1(_1346_),
    .A2(_0369_),
    .B1(_1718_),
    .Y(_1719_));
 sky130_fd_sc_hd__a221oi_1 _5243_ (.A1(_0335_),
    .A2(_0362_),
    .B1(_0323_),
    .B2(_0366_),
    .C1(_1719_),
    .Y(_1720_));
 sky130_fd_sc_hd__nand2_1 _5244_ (.A(_0388_),
    .B(_0701_),
    .Y(_1721_));
 sky130_fd_sc_hd__o21ai_1 _5245_ (.A1(_0705_),
    .A2(_0386_),
    .B1(_1721_),
    .Y(_1722_));
 sky130_fd_sc_hd__a221oi_1 _5246_ (.A1(_0703_),
    .A2(_0379_),
    .B1(_0400_),
    .B2(_0383_),
    .C1(_1722_),
    .Y(_1723_));
 sky130_fd_sc_hd__and4_1 _5247_ (.A(_1713_),
    .B(_1717_),
    .C(_1720_),
    .D(_1723_),
    .X(_1724_));
 sky130_fd_sc_hd__nand2_1 _5248_ (.A(_0399_),
    .B(_0455_),
    .Y(_1725_));
 sky130_fd_sc_hd__nand2_1 _5249_ (.A(_0403_),
    .B(_0451_),
    .Y(_1726_));
 sky130_fd_sc_hd__or2_1 _5250_ (.A(_3108_),
    .B(_0408_),
    .X(_1727_));
 sky130_fd_sc_hd__o2111a_1 _5251_ (.A1(_0981_),
    .A2(_0397_),
    .B1(_1725_),
    .C1(_1726_),
    .D1(_1727_),
    .X(_1728_));
 sky130_fd_sc_hd__nand2_1 _5252_ (.A(_0416_),
    .B(_3115_),
    .Y(_1729_));
 sky130_fd_sc_hd__nand2_1 _5253_ (.A(_0420_),
    .B(_3102_),
    .Y(_1730_));
 sky130_fd_sc_hd__or2_1 _5254_ (.A(_0767_),
    .B(_0426_),
    .X(_1731_));
 sky130_fd_sc_hd__o2111a_1 _5255_ (.A1(_1034_),
    .A2(_0414_),
    .B1(_1729_),
    .C1(_1730_),
    .D1(_1731_),
    .X(_1732_));
 sky130_fd_sc_hd__nand2_1 _5256_ (.A(_0442_),
    .B(_0421_),
    .Y(_1733_));
 sky130_fd_sc_hd__o21ai_1 _5257_ (.A1(_0424_),
    .A2(_0440_),
    .B1(_1733_),
    .Y(_1734_));
 sky130_fd_sc_hd__a221oi_1 _5258_ (.A1(_0411_),
    .A2(_0432_),
    .B1(_0447_),
    .B2(_0436_),
    .C1(_1734_),
    .Y(_1735_));
 sky130_fd_sc_hd__nand2_1 _5259_ (.A(_0460_),
    .B(_3119_),
    .Y(_1736_));
 sky130_fd_sc_hd__o21ai_1 _5260_ (.A1(_3077_),
    .A2(_0458_),
    .B1(_1736_),
    .Y(_1737_));
 sky130_fd_sc_hd__a221oi_1 _5261_ (.A1(_3136_),
    .A2(_0450_),
    .B1(_3134_),
    .B2(_0454_),
    .C1(_1737_),
    .Y(_1738_));
 sky130_fd_sc_hd__and4_1 _5262_ (.A(_1728_),
    .B(_1732_),
    .C(_1735_),
    .D(_1738_),
    .X(_1739_));
 sky130_fd_sc_hd__and2_1 _5263_ (.A(_1724_),
    .B(_1739_),
    .X(_1740_));
 sky130_fd_sc_hd__inv_2 _5264_ (.A(\egd_top.BitStream_buffer.BS_buffer[33] ),
    .Y(_1741_));
 sky130_fd_sc_hd__nand2_1 _5265_ (.A(_0474_),
    .B(_0689_),
    .Y(_1742_));
 sky130_fd_sc_hd__a22o_1 _5266_ (.A1(_0478_),
    .A2(_0372_),
    .B1(_0481_),
    .B2(_0691_),
    .X(_1743_));
 sky130_fd_sc_hd__inv_2 _5267_ (.A(_1743_),
    .Y(_1744_));
 sky130_fd_sc_hd__o211a_1 _5268_ (.A1(_1741_),
    .A2(_0472_),
    .B1(_1742_),
    .C1(_1744_),
    .X(_1745_));
 sky130_fd_sc_hd__nand2_1 _5269_ (.A(_0498_),
    .B(_0535_),
    .Y(_1746_));
 sky130_fd_sc_hd__o21ai_1 _5270_ (.A1(_0995_),
    .A2(_0496_),
    .B1(_1746_),
    .Y(_1747_));
 sky130_fd_sc_hd__a221oi_1 _5271_ (.A1(_0475_),
    .A2(_0488_),
    .B1(_0479_),
    .B2(_0492_),
    .C1(_1747_),
    .Y(_1748_));
 sky130_fd_sc_hd__nand2_1 _5272_ (.A(_0508_),
    .B(_0525_),
    .Y(_1749_));
 sky130_fd_sc_hd__nand2_1 _5273_ (.A(_0512_),
    .B(_0531_),
    .Y(_1750_));
 sky130_fd_sc_hd__or2_1 _5274_ (.A(_1373_),
    .B(_0518_),
    .X(_1751_));
 sky130_fd_sc_hd__o2111a_1 _5275_ (.A1(_1619_),
    .A2(_0506_),
    .B1(_1749_),
    .C1(_1750_),
    .D1(_1751_),
    .X(_1752_));
 sky130_fd_sc_hd__nand2_1 _5276_ (.A(_0530_),
    .B(_0353_),
    .Y(_1753_));
 sky130_fd_sc_hd__nand2_1 _5277_ (.A(_0534_),
    .B(_0346_),
    .Y(_1754_));
 sky130_fd_sc_hd__nand2_1 _5278_ (.A(_1753_),
    .B(_1754_),
    .Y(_1755_));
 sky130_fd_sc_hd__a221oi_1 _5279_ (.A1(_0356_),
    .A2(_0524_),
    .B1(_0339_),
    .B2(_0528_),
    .C1(_1755_),
    .Y(_1756_));
 sky130_fd_sc_hd__and4_1 _5280_ (.A(_1745_),
    .B(_1748_),
    .C(_1752_),
    .D(_1756_),
    .X(_1757_));
 sky130_fd_sc_hd__nand2_1 _5281_ (.A(_0547_),
    .B(\egd_top.BitStream_buffer.BS_buffer[15] ),
    .Y(_1758_));
 sky130_fd_sc_hd__nand2_1 _5282_ (.A(_0551_),
    .B(\egd_top.BitStream_buffer.BS_buffer[13] ),
    .Y(_1759_));
 sky130_fd_sc_hd__or2_1 _5283_ (.A(_1022_),
    .B(_0556_),
    .X(_1760_));
 sky130_fd_sc_hd__o2111a_1 _5284_ (.A1(_0756_),
    .A2(_0545_),
    .B1(_1758_),
    .C1(_1759_),
    .D1(_1760_),
    .X(_1761_));
 sky130_fd_sc_hd__nand2_1 _5285_ (.A(_0563_),
    .B(_0499_),
    .Y(_1762_));
 sky130_fd_sc_hd__nand2_1 _5286_ (.A(_0566_),
    .B(_0489_),
    .Y(_1763_));
 sky130_fd_sc_hd__or2_1 _5287_ (.A(_0494_),
    .B(_0570_),
    .X(_1764_));
 sky130_fd_sc_hd__o2111a_1 _5288_ (.A1(_0867_),
    .A2(_0561_),
    .B1(_1762_),
    .C1(_1763_),
    .D1(_1764_),
    .X(_1765_));
 sky130_fd_sc_hd__or2_1 _5289_ (.A(_0593_),
    .B(_0584_),
    .X(_1766_));
 sky130_fd_sc_hd__o221a_1 _5290_ (.A1(_0559_),
    .A2(_0576_),
    .B1(_0750_),
    .B2(_0580_),
    .C1(_1766_),
    .X(_1767_));
 sky130_fd_sc_hd__o22ai_1 _5291_ (.A1(_0516_),
    .A2(_0595_),
    .B1(_0734_),
    .B2(_0598_),
    .Y(_1768_));
 sky130_fd_sc_hd__a221oi_1 _5292_ (.A1(_0503_),
    .A2(_0589_),
    .B1(_0467_),
    .B2(_0592_),
    .C1(_1768_),
    .Y(_1769_));
 sky130_fd_sc_hd__and4_1 _5293_ (.A(_1761_),
    .B(_1765_),
    .C(_1767_),
    .D(_1769_),
    .X(_1770_));
 sky130_fd_sc_hd__and3_1 _5294_ (.A(_1740_),
    .B(_1757_),
    .C(_1770_),
    .X(_1771_));
 sky130_fd_sc_hd__nand2_1 _5295_ (.A(_0606_),
    .B(\egd_top.BitStream_buffer.BS_buffer[9] ),
    .Y(_1772_));
 sky130_fd_sc_hd__nand3_1 _5296_ (.A(_1709_),
    .B(_1771_),
    .C(_1772_),
    .Y(_1773_));
 sky130_fd_sc_hd__inv_2 _5297_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[6] ),
    .Y(_1774_));
 sky130_fd_sc_hd__a21oi_1 _5298_ (.A1(_1774_),
    .A2(_0898_),
    .B1(_2938_),
    .Y(_1775_));
 sky130_fd_sc_hd__o21a_1 _5299_ (.A1(_3056_),
    .A2(_1773_),
    .B1(_1775_),
    .X(_0288_));
 sky130_fd_sc_hd__inv_2 _5300_ (.A(\egd_top.BitStream_buffer.BS_buffer[83] ),
    .Y(_1776_));
 sky130_fd_sc_hd__o22ai_1 _5301_ (.A1(_1654_),
    .A2(_3084_),
    .B1(_1776_),
    .B2(_3092_),
    .Y(_1777_));
 sky130_fd_sc_hd__a221oi_1 _5302_ (.A1(_0646_),
    .A2(_3068_),
    .B1(_3265_),
    .B2(_3075_),
    .C1(_1777_),
    .Y(_1778_));
 sky130_fd_sc_hd__nand2_1 _5303_ (.A(_3114_),
    .B(_3069_),
    .Y(_1779_));
 sky130_fd_sc_hd__o21ai_1 _5304_ (.A1(_0611_),
    .A2(_3111_),
    .B1(_1779_),
    .Y(_1780_));
 sky130_fd_sc_hd__a221oi_2 _5305_ (.A1(_3161_),
    .A2(_3101_),
    .B1(_3156_),
    .B2(_3106_),
    .C1(_1780_),
    .Y(_1781_));
 sky130_fd_sc_hd__nand2_1 _5306_ (.A(_3128_),
    .B(_3144_),
    .Y(_1782_));
 sky130_fd_sc_hd__nand2_1 _5307_ (.A(_3133_),
    .B(_3255_),
    .Y(_1783_));
 sky130_fd_sc_hd__or2_1 _5308_ (.A(_1284_),
    .B(_3141_),
    .X(_1784_));
 sky130_fd_sc_hd__o2111a_1 _5309_ (.A1(_1532_),
    .A2(_3124_),
    .B1(_1782_),
    .C1(_1783_),
    .D1(_1784_),
    .X(_1785_));
 sky130_fd_sc_hd__nand2_1 _5310_ (.A(_3155_),
    .B(_3275_),
    .Y(_1786_));
 sky130_fd_sc_hd__nand2_1 _5311_ (.A(_3160_),
    .B(_3272_),
    .Y(_1787_));
 sky130_fd_sc_hd__nand2_1 _5312_ (.A(_1786_),
    .B(_1787_),
    .Y(_1788_));
 sky130_fd_sc_hd__a221oi_1 _5313_ (.A1(_0653_),
    .A2(_3148_),
    .B1(_0804_),
    .B2(_3152_),
    .C1(_1788_),
    .Y(_1789_));
 sky130_fd_sc_hd__and4_1 _5314_ (.A(_1778_),
    .B(_1781_),
    .C(_1785_),
    .D(_1789_),
    .X(_1790_));
 sky130_fd_sc_hd__o22ai_1 _5315_ (.A1(_0638_),
    .A2(_3176_),
    .B1(_0790_),
    .B2(_3179_),
    .Y(_1791_));
 sky130_fd_sc_hd__a221oi_1 _5316_ (.A1(_0607_),
    .A2(_3170_),
    .B1(_0577_),
    .B2(_3173_),
    .C1(_1791_),
    .Y(_1792_));
 sky130_fd_sc_hd__nand2_1 _5317_ (.A(_3192_),
    .B(_0552_),
    .Y(_1793_));
 sky130_fd_sc_hd__o21ai_1 _5318_ (.A1(_0541_),
    .A2(_3190_),
    .B1(_1793_),
    .Y(_1794_));
 sky130_fd_sc_hd__a221oi_1 _5319_ (.A1(_0573_),
    .A2(_3184_),
    .B1(_0581_),
    .B2(_3187_),
    .C1(_1794_),
    .Y(_1795_));
 sky130_fd_sc_hd__nand2_1 _5320_ (.A(_3206_),
    .B(_3040_),
    .Y(_1796_));
 sky130_fd_sc_hd__o21ai_1 _5321_ (.A1(_1174_),
    .A2(_3204_),
    .B1(_1796_),
    .Y(_1797_));
 sky130_fd_sc_hd__a221oi_1 _5322_ (.A1(_3044_),
    .A2(_3198_),
    .B1(_3047_),
    .B2(_3201_),
    .C1(_1797_),
    .Y(_1798_));
 sky130_fd_sc_hd__o22ai_1 _5323_ (.A1(_0742_),
    .A2(_3218_),
    .B1(_0554_),
    .B2(_3221_),
    .Y(_1799_));
 sky130_fd_sc_hd__a221oi_1 _5324_ (.A1(\egd_top.BitStream_buffer.BS_buffer[8] ),
    .A2(_3212_),
    .B1(\egd_top.BitStream_buffer.BS_buffer[9] ),
    .B2(_3215_),
    .C1(_1799_),
    .Y(_1800_));
 sky130_fd_sc_hd__and4_1 _5325_ (.A(_1792_),
    .B(_1795_),
    .C(_1798_),
    .D(_1800_),
    .X(_1801_));
 sky130_fd_sc_hd__o22ai_1 _5326_ (.A1(_1196_),
    .A2(_3238_),
    .B1(_1320_),
    .B2(_3241_),
    .Y(_1802_));
 sky130_fd_sc_hd__a221oi_1 _5327_ (.A1(_3341_),
    .A2(_3231_),
    .B1(_3347_),
    .B2(_3235_),
    .C1(_1802_),
    .Y(_1803_));
 sky130_fd_sc_hd__nand2_1 _5328_ (.A(_3246_),
    .B(_3232_),
    .Y(_1804_));
 sky130_fd_sc_hd__nand2_1 _5329_ (.A(_3250_),
    .B(_3290_),
    .Y(_1805_));
 sky130_fd_sc_hd__nand2_1 _5330_ (.A(_3254_),
    .B(_3225_),
    .Y(_1806_));
 sky130_fd_sc_hd__nand2_1 _5331_ (.A(_3258_),
    .B(_3286_),
    .Y(_1807_));
 sky130_fd_sc_hd__and4_1 _5332_ (.A(_1804_),
    .B(_1805_),
    .C(_1806_),
    .D(_1807_),
    .X(_1808_));
 sky130_fd_sc_hd__o22ai_1 _5333_ (.A1(_0656_),
    .A2(_3264_),
    .B1(_0807_),
    .B2(_3268_),
    .Y(_1809_));
 sky130_fd_sc_hd__a22o_1 _5334_ (.A1(_3271_),
    .A2(_3318_),
    .B1(_3274_),
    .B2(_3322_),
    .X(_1810_));
 sky130_fd_sc_hd__nor2_1 _5335_ (.A(_1809_),
    .B(_1810_),
    .Y(_1811_));
 sky130_fd_sc_hd__o22ai_1 _5336_ (.A1(_0671_),
    .A2(_3289_),
    .B1(_3336_),
    .B2(_3293_),
    .Y(_1812_));
 sky130_fd_sc_hd__a221oi_1 _5337_ (.A1(_3314_),
    .A2(_3281_),
    .B1(_3310_),
    .B2(_3285_),
    .C1(_1812_),
    .Y(_1813_));
 sky130_fd_sc_hd__and4_1 _5338_ (.A(_1803_),
    .B(_1808_),
    .C(_1811_),
    .D(_1813_),
    .X(_1814_));
 sky130_fd_sc_hd__nand2_1 _5339_ (.A(_3309_),
    .B(_3016_),
    .Y(_1815_));
 sky130_fd_sc_hd__nand2_1 _5340_ (.A(_3313_),
    .B(_3013_),
    .Y(_1816_));
 sky130_fd_sc_hd__nand2_1 _5341_ (.A(_1815_),
    .B(_1816_),
    .Y(_1817_));
 sky130_fd_sc_hd__a221oi_1 _5342_ (.A1(_3019_),
    .A2(_3303_),
    .B1(_3022_),
    .B2(_3307_),
    .C1(_1817_),
    .Y(_1818_));
 sky130_fd_sc_hd__nand2_1 _5343_ (.A(_3326_),
    .B(_3357_),
    .Y(_1819_));
 sky130_fd_sc_hd__nand2_1 _5344_ (.A(_3330_),
    .B(_3353_),
    .Y(_1820_));
 sky130_fd_sc_hd__nand2_1 _5345_ (.A(_1819_),
    .B(_1820_),
    .Y(_1821_));
 sky130_fd_sc_hd__a221oi_1 _5346_ (.A1(_3297_),
    .A2(_3321_),
    .B1(_3304_),
    .B2(_3324_),
    .C1(_1821_),
    .Y(_1822_));
 sky130_fd_sc_hd__nand2_1 _5347_ (.A(_3340_),
    .B(\egd_top.BitStream_buffer.BS_buffer[110] ),
    .Y(_1823_));
 sky130_fd_sc_hd__nand2_1 _5348_ (.A(_3344_),
    .B(_2998_),
    .Y(_1824_));
 sky130_fd_sc_hd__or2_1 _5349_ (.A(_3361_),
    .B(_3350_),
    .X(_1825_));
 sky130_fd_sc_hd__o2111a_1 _5350_ (.A1(_0634_),
    .A2(_3338_),
    .B1(_1823_),
    .C1(_1824_),
    .D1(_1825_),
    .X(_1826_));
 sky130_fd_sc_hd__nand2_1 _5351_ (.A(_3365_),
    .B(_3031_),
    .Y(_1827_));
 sky130_fd_sc_hd__o21ai_1 _5352_ (.A1(_1047_),
    .A2(_3363_),
    .B1(_1827_),
    .Y(_1828_));
 sky130_fd_sc_hd__a221oi_1 _5353_ (.A1(_3025_),
    .A2(_3356_),
    .B1(_3028_),
    .B2(_3360_),
    .C1(_1828_),
    .Y(_1829_));
 sky130_fd_sc_hd__and4_1 _5354_ (.A(_1818_),
    .B(_1822_),
    .C(_1826_),
    .D(_1829_),
    .X(_1830_));
 sky130_fd_sc_hd__and4_1 _5355_ (.A(_1790_),
    .B(_1801_),
    .C(_1814_),
    .D(_1830_),
    .X(_1831_));
 sky130_fd_sc_hd__nand2_1 _5356_ (.A(_0334_),
    .B(_0433_),
    .Y(_1832_));
 sky130_fd_sc_hd__nand2_1 _5357_ (.A(_0338_),
    .B(_0429_),
    .Y(_1833_));
 sky130_fd_sc_hd__nand2_1 _5358_ (.A(_1832_),
    .B(_1833_),
    .Y(_1834_));
 sky130_fd_sc_hd__a221oi_1 _5359_ (.A1(_0404_),
    .A2(_0328_),
    .B1(_0703_),
    .B2(_0332_),
    .C1(_1834_),
    .Y(_1835_));
 sky130_fd_sc_hd__o22ai_1 _5360_ (.A1(_1714_),
    .A2(_0345_),
    .B1(_0384_),
    .B2(_0349_),
    .Y(_1836_));
 sky130_fd_sc_hd__a22o_1 _5361_ (.A1(_0352_),
    .A2(_0437_),
    .B1(_0355_),
    .B2(_0443_),
    .X(_1837_));
 sky130_fd_sc_hd__nor2_1 _5362_ (.A(_1836_),
    .B(_1837_),
    .Y(_1838_));
 sky130_fd_sc_hd__nand2_1 _5363_ (.A(_0371_),
    .B(_0380_),
    .Y(_1839_));
 sky130_fd_sc_hd__o21ai_1 _5364_ (.A1(_1470_),
    .A2(_0369_),
    .B1(_1839_),
    .Y(_1840_));
 sky130_fd_sc_hd__a221oi_1 _5365_ (.A1(_0323_),
    .A2(_0362_),
    .B1(_0329_),
    .B2(_0366_),
    .C1(_1840_),
    .Y(_1841_));
 sky130_fd_sc_hd__nand2_1 _5366_ (.A(_0388_),
    .B(_0417_),
    .Y(_1842_));
 sky130_fd_sc_hd__o21ai_1 _5367_ (.A1(_0424_),
    .A2(_0386_),
    .B1(_1842_),
    .Y(_1843_));
 sky130_fd_sc_hd__a221oi_1 _5368_ (.A1(_0400_),
    .A2(_0379_),
    .B1(_0701_),
    .B2(_0383_),
    .C1(_1843_),
    .Y(_1844_));
 sky130_fd_sc_hd__and4_1 _5369_ (.A(_1835_),
    .B(_1838_),
    .C(_1841_),
    .D(_1844_),
    .X(_1845_));
 sky130_fd_sc_hd__nand2_1 _5370_ (.A(_0399_),
    .B(_3107_),
    .Y(_1846_));
 sky130_fd_sc_hd__nand2_1 _5371_ (.A(_0403_),
    .B(_0461_),
    .Y(_1847_));
 sky130_fd_sc_hd__or2_1 _5372_ (.A(_0614_),
    .B(_0408_),
    .X(_1848_));
 sky130_fd_sc_hd__o2111a_1 _5373_ (.A1(_0456_),
    .A2(_0397_),
    .B1(_1846_),
    .C1(_1847_),
    .D1(_1848_),
    .X(_1849_));
 sky130_fd_sc_hd__nand2_1 _5374_ (.A(_0416_),
    .B(_3095_),
    .Y(_1850_));
 sky130_fd_sc_hd__nand2_1 _5375_ (.A(_0420_),
    .B(_3129_),
    .Y(_1851_));
 sky130_fd_sc_hd__or2_1 _5376_ (.A(_0903_),
    .B(_0426_),
    .X(_1852_));
 sky130_fd_sc_hd__o2111a_1 _5377_ (.A1(_3137_),
    .A2(_0414_),
    .B1(_1850_),
    .C1(_1851_),
    .D1(_1852_),
    .X(_1853_));
 sky130_fd_sc_hd__nand2_1 _5378_ (.A(_0442_),
    .B(_0411_),
    .Y(_1854_));
 sky130_fd_sc_hd__o21ai_1 _5379_ (.A1(_0711_),
    .A2(_0440_),
    .B1(_1854_),
    .Y(_1855_));
 sky130_fd_sc_hd__a221oi_1 _5380_ (.A1(_0447_),
    .A2(_0432_),
    .B1(_0451_),
    .B2(_0436_),
    .C1(_1855_),
    .Y(_1856_));
 sky130_fd_sc_hd__nand2_1 _5381_ (.A(_0460_),
    .B(_3076_),
    .Y(_1857_));
 sky130_fd_sc_hd__o21ai_1 _5382_ (.A1(_3086_),
    .A2(_0458_),
    .B1(_1857_),
    .Y(_1858_));
 sky130_fd_sc_hd__a221oi_1 _5383_ (.A1(_3134_),
    .A2(_0450_),
    .B1(_3119_),
    .B2(_0454_),
    .C1(_1858_),
    .Y(_1859_));
 sky130_fd_sc_hd__and4_1 _5384_ (.A(_1849_),
    .B(_1853_),
    .C(_1856_),
    .D(_1859_),
    .X(_1860_));
 sky130_fd_sc_hd__and2_1 _5385_ (.A(_1845_),
    .B(_1860_),
    .X(_1861_));
 sky130_fd_sc_hd__nand2_1 _5386_ (.A(_0474_),
    .B(_0372_),
    .Y(_1862_));
 sky130_fd_sc_hd__a22o_1 _5387_ (.A1(_0478_),
    .A2(_0691_),
    .B1(_0481_),
    .B2(_0346_),
    .X(_1863_));
 sky130_fd_sc_hd__inv_2 _5388_ (.A(_1863_),
    .Y(_1864_));
 sky130_fd_sc_hd__o211a_1 _5389_ (.A1(_0367_),
    .A2(_0472_),
    .B1(_1862_),
    .C1(_1864_),
    .X(_1865_));
 sky130_fd_sc_hd__nand2_1 _5390_ (.A(_0498_),
    .B(_0531_),
    .Y(_1866_));
 sky130_fd_sc_hd__o21ai_1 _5391_ (.A1(_1123_),
    .A2(_0496_),
    .B1(_1866_),
    .Y(_1867_));
 sky130_fd_sc_hd__a221oi_1 _5392_ (.A1(_0479_),
    .A2(_0488_),
    .B1(_0482_),
    .B2(_0492_),
    .C1(_1867_),
    .Y(_1868_));
 sky130_fd_sc_hd__nand2_1 _5393_ (.A(_0508_),
    .B(_0359_),
    .Y(_1869_));
 sky130_fd_sc_hd__nand2_1 _5394_ (.A(_0512_),
    .B(_0521_),
    .Y(_1870_));
 sky130_fd_sc_hd__or2_1 _5395_ (.A(_1497_),
    .B(_0518_),
    .X(_1871_));
 sky130_fd_sc_hd__o2111a_1 _5396_ (.A1(_1741_),
    .A2(_0506_),
    .B1(_1869_),
    .C1(_1870_),
    .D1(_1871_),
    .X(_1872_));
 sky130_fd_sc_hd__nand2_1 _5397_ (.A(_0530_),
    .B(_0356_),
    .Y(_1873_));
 sky130_fd_sc_hd__nand2_1 _5398_ (.A(_0534_),
    .B(_0353_),
    .Y(_1874_));
 sky130_fd_sc_hd__nand2_1 _5399_ (.A(_1873_),
    .B(_1874_),
    .Y(_1875_));
 sky130_fd_sc_hd__a221oi_1 _5400_ (.A1(_0339_),
    .A2(_0524_),
    .B1(_0335_),
    .B2(_0528_),
    .C1(_1875_),
    .Y(_1876_));
 sky130_fd_sc_hd__and4_1 _5401_ (.A(_1865_),
    .B(_1868_),
    .C(_1872_),
    .D(_1876_),
    .X(_1877_));
 sky130_fd_sc_hd__nand2_1 _5402_ (.A(_0547_),
    .B(\egd_top.BitStream_buffer.BS_buffer[16] ),
    .Y(_1878_));
 sky130_fd_sc_hd__nand2_1 _5403_ (.A(_0551_),
    .B(\egd_top.BitStream_buffer.BS_buffer[14] ),
    .Y(_1879_));
 sky130_fd_sc_hd__or2_1 _5404_ (.A(_1150_),
    .B(_0556_),
    .X(_1880_));
 sky130_fd_sc_hd__o2111a_1 _5405_ (.A1(_0890_),
    .A2(_0545_),
    .B1(_1878_),
    .C1(_1879_),
    .D1(_1880_),
    .X(_1881_));
 sky130_fd_sc_hd__nand2_1 _5406_ (.A(_0563_),
    .B(_0513_),
    .Y(_1882_));
 sky130_fd_sc_hd__nand2_1 _5407_ (.A(_0566_),
    .B(_0493_),
    .Y(_1883_));
 sky130_fd_sc_hd__or2_1 _5408_ (.A(_0728_),
    .B(_0570_),
    .X(_1884_));
 sky130_fd_sc_hd__o2111a_1 _5409_ (.A1(_0516_),
    .A2(_0561_),
    .B1(_1882_),
    .C1(_1883_),
    .D1(_1884_),
    .X(_1885_));
 sky130_fd_sc_hd__or2_1 _5410_ (.A(_0596_),
    .B(_0584_),
    .X(_1886_));
 sky130_fd_sc_hd__o221a_1 _5411_ (.A1(_0593_),
    .A2(_0576_),
    .B1(_0559_),
    .B2(_0580_),
    .C1(_1886_),
    .X(_1887_));
 sky130_fd_sc_hd__o22ai_1 _5412_ (.A1(_0734_),
    .A2(_0595_),
    .B1(_0504_),
    .B2(_0598_),
    .Y(_1888_));
 sky130_fd_sc_hd__a221oi_1 _5413_ (.A1(_0467_),
    .A2(_0589_),
    .B1(_0475_),
    .B2(_0592_),
    .C1(_1888_),
    .Y(_1889_));
 sky130_fd_sc_hd__and4_1 _5414_ (.A(_1881_),
    .B(_1885_),
    .C(_1887_),
    .D(_1889_),
    .X(_1890_));
 sky130_fd_sc_hd__and3_1 _5415_ (.A(_1861_),
    .B(_1877_),
    .C(_1890_),
    .X(_1891_));
 sky130_fd_sc_hd__nand2_1 _5416_ (.A(_0606_),
    .B(\egd_top.BitStream_buffer.BS_buffer[10] ),
    .Y(_1892_));
 sky130_fd_sc_hd__nand3_1 _5417_ (.A(_1831_),
    .B(_1891_),
    .C(_1892_),
    .Y(_1893_));
 sky130_fd_sc_hd__inv_2 _5418_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[5] ),
    .Y(_1894_));
 sky130_fd_sc_hd__a21oi_1 _5419_ (.A1(_1894_),
    .A2(_0898_),
    .B1(_2938_),
    .Y(_1895_));
 sky130_fd_sc_hd__o21a_1 _5420_ (.A1(_3056_),
    .A2(_1893_),
    .B1(_1895_),
    .X(_0287_));
 sky130_fd_sc_hd__o22ai_1 _5421_ (.A1(_1776_),
    .A2(_3084_),
    .B1(_3262_),
    .B2(_3092_),
    .Y(_1896_));
 sky130_fd_sc_hd__a221oi_1 _5422_ (.A1(_3265_),
    .A2(_3068_),
    .B1(_3272_),
    .B2(_3075_),
    .C1(_1896_),
    .Y(_1897_));
 sky130_fd_sc_hd__nand2_1 _5423_ (.A(_3114_),
    .B(_3161_),
    .Y(_1898_));
 sky130_fd_sc_hd__o21ai_1 _5424_ (.A1(_0764_),
    .A2(_3111_),
    .B1(_1898_),
    .Y(_1899_));
 sky130_fd_sc_hd__a221oi_1 _5425_ (.A1(_3156_),
    .A2(_3101_),
    .B1(_3144_),
    .B2(_3106_),
    .C1(_1899_),
    .Y(_1900_));
 sky130_fd_sc_hd__nand2_1 _5426_ (.A(_3128_),
    .B(_3149_),
    .Y(_1901_));
 sky130_fd_sc_hd__nand2_1 _5427_ (.A(_3133_),
    .B(_3247_),
    .Y(_1902_));
 sky130_fd_sc_hd__or2_1 _5428_ (.A(_1408_),
    .B(_3141_),
    .X(_1903_));
 sky130_fd_sc_hd__o2111a_1 _5429_ (.A1(_1654_),
    .A2(_3124_),
    .B1(_1901_),
    .C1(_1902_),
    .D1(_1903_),
    .X(_1904_));
 sky130_fd_sc_hd__nand2_1 _5430_ (.A(_3155_),
    .B(_0653_),
    .Y(_1905_));
 sky130_fd_sc_hd__nand2_1 _5431_ (.A(_3160_),
    .B(_3275_),
    .Y(_1906_));
 sky130_fd_sc_hd__nand2_1 _5432_ (.A(_1905_),
    .B(_1906_),
    .Y(_1907_));
 sky130_fd_sc_hd__a221oi_1 _5433_ (.A1(_0804_),
    .A2(_3148_),
    .B1(_3225_),
    .B2(_3152_),
    .C1(_1907_),
    .Y(_1908_));
 sky130_fd_sc_hd__and4_1 _5434_ (.A(_1897_),
    .B(_1900_),
    .C(_1904_),
    .D(_1908_),
    .X(_1909_));
 sky130_fd_sc_hd__o22ai_1 _5435_ (.A1(_0790_),
    .A2(_3176_),
    .B1(_0926_),
    .B2(_3179_),
    .Y(_1910_));
 sky130_fd_sc_hd__a221oi_1 _5436_ (.A1(_0577_),
    .A2(_3170_),
    .B1(_0573_),
    .B2(_3173_),
    .C1(_1910_),
    .Y(_1911_));
 sky130_fd_sc_hd__nand2_1 _5437_ (.A(_3192_),
    .B(_0540_),
    .Y(_1912_));
 sky130_fd_sc_hd__o21ai_1 _5438_ (.A1(_0742_),
    .A2(_3190_),
    .B1(_1912_),
    .Y(_1913_));
 sky130_fd_sc_hd__a221oi_1 _5439_ (.A1(_0581_),
    .A2(_3184_),
    .B1(_0552_),
    .B2(_3187_),
    .C1(_1913_),
    .Y(_1914_));
 sky130_fd_sc_hd__nand2_1 _5440_ (.A(_3206_),
    .B(_3044_),
    .Y(_1915_));
 sky130_fd_sc_hd__o21ai_1 _5441_ (.A1(_3188_),
    .A2(_3204_),
    .B1(_1915_),
    .Y(_1916_));
 sky130_fd_sc_hd__a221oi_1 _5442_ (.A1(_3047_),
    .A2(_3198_),
    .B1(_3050_),
    .B2(_3201_),
    .C1(_1916_),
    .Y(_1917_));
 sky130_fd_sc_hd__o22ai_1 _5443_ (.A1(_0554_),
    .A2(_3218_),
    .B1(_0745_),
    .B2(_3221_),
    .Y(_1918_));
 sky130_fd_sc_hd__a221oi_1 _5444_ (.A1(\egd_top.BitStream_buffer.BS_buffer[9] ),
    .A2(_3212_),
    .B1(\egd_top.BitStream_buffer.BS_buffer[10] ),
    .B2(_3215_),
    .C1(_1918_),
    .Y(_1919_));
 sky130_fd_sc_hd__and4_1 _5445_ (.A(_1911_),
    .B(_1914_),
    .C(_1917_),
    .D(_1919_),
    .X(_1920_));
 sky130_fd_sc_hd__o22ai_1 _5446_ (.A1(_1320_),
    .A2(_3238_),
    .B1(_1444_),
    .B2(_3241_),
    .Y(_1921_));
 sky130_fd_sc_hd__a221oi_1 _5447_ (.A1(_3347_),
    .A2(_3231_),
    .B1(_3345_),
    .B2(_3235_),
    .C1(_1921_),
    .Y(_1922_));
 sky130_fd_sc_hd__nand2_1 _5448_ (.A(_3246_),
    .B(_3286_),
    .Y(_1923_));
 sky130_fd_sc_hd__nand2_1 _5449_ (.A(_3250_),
    .B(_3278_),
    .Y(_1924_));
 sky130_fd_sc_hd__nand2_1 _5450_ (.A(_3254_),
    .B(_3232_),
    .Y(_1925_));
 sky130_fd_sc_hd__nand2_1 _5451_ (.A(_3258_),
    .B(_3290_),
    .Y(_1926_));
 sky130_fd_sc_hd__and4_1 _5452_ (.A(_1923_),
    .B(_1924_),
    .C(_1925_),
    .D(_1926_),
    .X(_1927_));
 sky130_fd_sc_hd__o22ai_1 _5453_ (.A1(_0807_),
    .A2(_3264_),
    .B1(_0940_),
    .B2(_3268_),
    .Y(_1928_));
 sky130_fd_sc_hd__a22o_1 _5454_ (.A1(_3271_),
    .A2(_3322_),
    .B1(_3274_),
    .B2(_3331_),
    .X(_1929_));
 sky130_fd_sc_hd__nor2_1 _5455_ (.A(_1928_),
    .B(_1929_),
    .Y(_1930_));
 sky130_fd_sc_hd__o22ai_1 _5456_ (.A1(_3336_),
    .A2(_3289_),
    .B1(_0668_),
    .B2(_3293_),
    .Y(_1931_));
 sky130_fd_sc_hd__a221oi_1 _5457_ (.A1(_3310_),
    .A2(_3281_),
    .B1(_3297_),
    .B2(_3285_),
    .C1(_1931_),
    .Y(_1932_));
 sky130_fd_sc_hd__and4_1 _5458_ (.A(_1922_),
    .B(_1927_),
    .C(_1930_),
    .D(_1932_),
    .X(_1933_));
 sky130_fd_sc_hd__nand2_1 _5459_ (.A(_3309_),
    .B(_3019_),
    .Y(_1934_));
 sky130_fd_sc_hd__nand2_1 _5460_ (.A(_3313_),
    .B(_3016_),
    .Y(_1935_));
 sky130_fd_sc_hd__nand2_1 _5461_ (.A(_1934_),
    .B(_1935_),
    .Y(_1936_));
 sky130_fd_sc_hd__a221oi_1 _5462_ (.A1(_3022_),
    .A2(_3303_),
    .B1(_3025_),
    .B2(_3307_),
    .C1(_1936_),
    .Y(_1937_));
 sky130_fd_sc_hd__nand2_1 _5463_ (.A(_3326_),
    .B(_0674_),
    .Y(_1938_));
 sky130_fd_sc_hd__nand2_1 _5464_ (.A(_3330_),
    .B(_3357_),
    .Y(_1939_));
 sky130_fd_sc_hd__nand2_1 _5465_ (.A(_1938_),
    .B(_1939_),
    .Y(_1940_));
 sky130_fd_sc_hd__a221oi_1 _5466_ (.A1(_3304_),
    .A2(_3321_),
    .B1(_3353_),
    .B2(_3324_),
    .C1(_1940_),
    .Y(_1941_));
 sky130_fd_sc_hd__nand2_1 _5467_ (.A(_3340_),
    .B(\egd_top.BitStream_buffer.BS_buffer[111] ),
    .Y(_1942_));
 sky130_fd_sc_hd__nand2_1 _5468_ (.A(_3344_),
    .B(_3010_),
    .Y(_1943_));
 sky130_fd_sc_hd__or2_1 _5469_ (.A(_3202_),
    .B(_3350_),
    .X(_1944_));
 sky130_fd_sc_hd__o2111a_1 _5470_ (.A1(_0786_),
    .A2(_3338_),
    .B1(_1942_),
    .C1(_1943_),
    .D1(_1944_),
    .X(_1945_));
 sky130_fd_sc_hd__nand2_1 _5471_ (.A(_3365_),
    .B(_3034_),
    .Y(_1946_));
 sky130_fd_sc_hd__o21ai_1 _5472_ (.A1(_1174_),
    .A2(_3363_),
    .B1(_1946_),
    .Y(_1947_));
 sky130_fd_sc_hd__a221oi_1 _5473_ (.A1(_3028_),
    .A2(_3356_),
    .B1(_3031_),
    .B2(_3360_),
    .C1(_1947_),
    .Y(_1948_));
 sky130_fd_sc_hd__and4_1 _5474_ (.A(_1937_),
    .B(_1941_),
    .C(_1945_),
    .D(_1948_),
    .X(_1949_));
 sky130_fd_sc_hd__and4_1 _5475_ (.A(_1909_),
    .B(_1920_),
    .C(_1933_),
    .D(_1949_),
    .X(_1950_));
 sky130_fd_sc_hd__nand2_1 _5476_ (.A(_0334_),
    .B(_0404_),
    .Y(_1951_));
 sky130_fd_sc_hd__nand2_1 _5477_ (.A(_0338_),
    .B(_0433_),
    .Y(_1952_));
 sky130_fd_sc_hd__nand2_1 _5478_ (.A(_1951_),
    .B(_1952_),
    .Y(_1953_));
 sky130_fd_sc_hd__a221oi_1 _5479_ (.A1(_0703_),
    .A2(_0328_),
    .B1(_0400_),
    .B2(_0332_),
    .C1(_1953_),
    .Y(_1954_));
 sky130_fd_sc_hd__o22ai_1 _5480_ (.A1(_0384_),
    .A2(_0345_),
    .B1(_0438_),
    .B2(_0349_),
    .Y(_1955_));
 sky130_fd_sc_hd__a22o_1 _5481_ (.A1(_0352_),
    .A2(_0443_),
    .B1(_0355_),
    .B2(_0429_),
    .X(_1956_));
 sky130_fd_sc_hd__nor2_1 _5482_ (.A(_1955_),
    .B(_1956_),
    .Y(_1957_));
 sky130_fd_sc_hd__nand2_1 _5483_ (.A(_0371_),
    .B(_0389_),
    .Y(_1958_));
 sky130_fd_sc_hd__o21ai_1 _5484_ (.A1(_1592_),
    .A2(_0369_),
    .B1(_1958_),
    .Y(_1959_));
 sky130_fd_sc_hd__a221oi_1 _5485_ (.A1(_0329_),
    .A2(_0362_),
    .B1(_0376_),
    .B2(_0366_),
    .C1(_1959_),
    .Y(_1960_));
 sky130_fd_sc_hd__nand2_1 _5486_ (.A(_0388_),
    .B(_0423_),
    .Y(_1961_));
 sky130_fd_sc_hd__o21ai_1 _5487_ (.A1(_0711_),
    .A2(_0386_),
    .B1(_1961_),
    .Y(_1962_));
 sky130_fd_sc_hd__a221oi_1 _5488_ (.A1(_0701_),
    .A2(_0379_),
    .B1(_0417_),
    .B2(_0383_),
    .C1(_1962_),
    .Y(_1963_));
 sky130_fd_sc_hd__and4_1 _5489_ (.A(_1954_),
    .B(_1957_),
    .C(_1960_),
    .D(_1963_),
    .X(_1964_));
 sky130_fd_sc_hd__nand2_1 _5490_ (.A(_0399_),
    .B(_3115_),
    .Y(_1965_));
 sky130_fd_sc_hd__nand2_1 _5491_ (.A(_0403_),
    .B(_0455_),
    .Y(_1966_));
 sky130_fd_sc_hd__or2_1 _5492_ (.A(_0767_),
    .B(_0408_),
    .X(_1967_));
 sky130_fd_sc_hd__o2111a_1 _5493_ (.A1(_3108_),
    .A2(_0397_),
    .B1(_1965_),
    .C1(_1966_),
    .D1(_1967_),
    .X(_1968_));
 sky130_fd_sc_hd__nand2_1 _5494_ (.A(_0416_),
    .B(_3102_),
    .Y(_1969_));
 sky130_fd_sc_hd__nand2_1 _5495_ (.A(_0420_),
    .B(_3136_),
    .Y(_1970_));
 sky130_fd_sc_hd__or2_1 _5496_ (.A(_1034_),
    .B(_0426_),
    .X(_1971_));
 sky130_fd_sc_hd__o2111a_1 _5497_ (.A1(_0620_),
    .A2(_0414_),
    .B1(_1969_),
    .C1(_1970_),
    .D1(_1971_),
    .X(_1972_));
 sky130_fd_sc_hd__nand2_1 _5498_ (.A(_0442_),
    .B(_0447_),
    .Y(_1973_));
 sky130_fd_sc_hd__o21ai_1 _5499_ (.A1(_0412_),
    .A2(_0440_),
    .B1(_1973_),
    .Y(_1974_));
 sky130_fd_sc_hd__a221oi_1 _5500_ (.A1(_0451_),
    .A2(_0432_),
    .B1(_0461_),
    .B2(_0436_),
    .C1(_1974_),
    .Y(_1975_));
 sky130_fd_sc_hd__nand2_1 _5501_ (.A(_0460_),
    .B(_3085_),
    .Y(_1976_));
 sky130_fd_sc_hd__o21ai_1 _5502_ (.A1(_0611_),
    .A2(_0458_),
    .B1(_1976_),
    .Y(_1977_));
 sky130_fd_sc_hd__a221oi_1 _5503_ (.A1(_3119_),
    .A2(_0450_),
    .B1(_3076_),
    .B2(_0454_),
    .C1(_1977_),
    .Y(_1978_));
 sky130_fd_sc_hd__and4_1 _5504_ (.A(_1968_),
    .B(_1972_),
    .C(_1975_),
    .D(_1978_),
    .X(_1979_));
 sky130_fd_sc_hd__and2_1 _5505_ (.A(_1964_),
    .B(_1979_),
    .X(_1980_));
 sky130_fd_sc_hd__nand2_1 _5506_ (.A(_0474_),
    .B(_0691_),
    .Y(_1981_));
 sky130_fd_sc_hd__a22o_1 _5507_ (.A1(_0478_),
    .A2(_0346_),
    .B1(_0481_),
    .B2(_0353_),
    .X(_1982_));
 sky130_fd_sc_hd__inv_2 _5508_ (.A(_1982_),
    .Y(_1983_));
 sky130_fd_sc_hd__o211a_1 _5509_ (.A1(_0690_),
    .A2(_0472_),
    .B1(_1981_),
    .C1(_1983_),
    .X(_1984_));
 sky130_fd_sc_hd__nand2_1 _5510_ (.A(_0498_),
    .B(_0521_),
    .Y(_1985_));
 sky130_fd_sc_hd__o21ai_1 _5511_ (.A1(_1249_),
    .A2(_0496_),
    .B1(_1985_),
    .Y(_1986_));
 sky130_fd_sc_hd__a221oi_1 _5512_ (.A1(_0482_),
    .A2(_0488_),
    .B1(_0535_),
    .B2(_0492_),
    .C1(_1986_),
    .Y(_1987_));
 sky130_fd_sc_hd__nand2_1 _5513_ (.A(_0508_),
    .B(_0363_),
    .Y(_1988_));
 sky130_fd_sc_hd__nand2_1 _5514_ (.A(_0512_),
    .B(_0525_),
    .Y(_1989_));
 sky130_fd_sc_hd__or2_1 _5515_ (.A(_1619_),
    .B(_0518_),
    .X(_1990_));
 sky130_fd_sc_hd__o2111a_1 _5516_ (.A1(_0367_),
    .A2(_0506_),
    .B1(_1988_),
    .C1(_1989_),
    .D1(_1990_),
    .X(_1991_));
 sky130_fd_sc_hd__nand2_1 _5517_ (.A(_0530_),
    .B(_0339_),
    .Y(_1992_));
 sky130_fd_sc_hd__nand2_1 _5518_ (.A(_0534_),
    .B(_0356_),
    .Y(_1993_));
 sky130_fd_sc_hd__nand2_1 _5519_ (.A(_1992_),
    .B(_1993_),
    .Y(_1994_));
 sky130_fd_sc_hd__a221oi_1 _5520_ (.A1(_0335_),
    .A2(_0524_),
    .B1(_0323_),
    .B2(_0528_),
    .C1(_1994_),
    .Y(_1995_));
 sky130_fd_sc_hd__and4_1 _5521_ (.A(_1984_),
    .B(_1987_),
    .C(_1991_),
    .D(_1995_),
    .X(_1996_));
 sky130_fd_sc_hd__nand2_1 _5522_ (.A(_0547_),
    .B(_0489_),
    .Y(_1997_));
 sky130_fd_sc_hd__nand2_1 _5523_ (.A(_0551_),
    .B(\egd_top.BitStream_buffer.BS_buffer[15] ),
    .Y(_1998_));
 sky130_fd_sc_hd__or2_1 _5524_ (.A(_0494_),
    .B(_0556_),
    .X(_1999_));
 sky130_fd_sc_hd__o2111a_1 _5525_ (.A1(_1022_),
    .A2(_0545_),
    .B1(_1997_),
    .C1(_1998_),
    .D1(_1999_),
    .X(_2000_));
 sky130_fd_sc_hd__nand2_1 _5526_ (.A(_0563_),
    .B(_0515_),
    .Y(_2001_));
 sky130_fd_sc_hd__nand2_1 _5527_ (.A(_0566_),
    .B(_0499_),
    .Y(_2002_));
 sky130_fd_sc_hd__or2_1 _5528_ (.A(_0867_),
    .B(_0570_),
    .X(_2003_));
 sky130_fd_sc_hd__o2111a_1 _5529_ (.A1(_0734_),
    .A2(_0561_),
    .B1(_2001_),
    .C1(_2002_),
    .D1(_2003_),
    .X(_2004_));
 sky130_fd_sc_hd__or2_1 _5530_ (.A(_0756_),
    .B(_0584_),
    .X(_2005_));
 sky130_fd_sc_hd__o221a_1 _5531_ (.A1(_0596_),
    .A2(_0576_),
    .B1(_0593_),
    .B2(_0580_),
    .C1(_2005_),
    .X(_2006_));
 sky130_fd_sc_hd__o22ai_1 _5532_ (.A1(_0504_),
    .A2(_0595_),
    .B1(_0468_),
    .B2(_0598_),
    .Y(_2007_));
 sky130_fd_sc_hd__a221oi_1 _5533_ (.A1(_0475_),
    .A2(_0589_),
    .B1(_0479_),
    .B2(_0592_),
    .C1(_2007_),
    .Y(_2008_));
 sky130_fd_sc_hd__and4_1 _5534_ (.A(_2000_),
    .B(_2004_),
    .C(_2006_),
    .D(_2008_),
    .X(_2009_));
 sky130_fd_sc_hd__and3_1 _5535_ (.A(_1980_),
    .B(_1996_),
    .C(_2009_),
    .X(_2010_));
 sky130_fd_sc_hd__nand2_1 _5536_ (.A(_0606_),
    .B(\egd_top.BitStream_buffer.BS_buffer[11] ),
    .Y(_2011_));
 sky130_fd_sc_hd__nand3_1 _5537_ (.A(_1950_),
    .B(_2010_),
    .C(_2011_),
    .Y(_2012_));
 sky130_fd_sc_hd__inv_2 _5538_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[4] ),
    .Y(_2013_));
 sky130_fd_sc_hd__a21oi_1 _5539_ (.A1(_2013_),
    .A2(_2996_),
    .B1(_2938_),
    .Y(_2014_));
 sky130_fd_sc_hd__o21a_1 _5540_ (.A1(_3056_),
    .A2(_2012_),
    .B1(_2014_),
    .X(_0286_));
 sky130_fd_sc_hd__o22ai_1 _5541_ (.A1(_3262_),
    .A2(_3083_),
    .B1(_3266_),
    .B2(_3091_),
    .Y(_2015_));
 sky130_fd_sc_hd__a221oi_1 _5542_ (.A1(_3272_),
    .A2(_3067_),
    .B1(_3275_),
    .B2(_3074_),
    .C1(_2015_),
    .Y(_2016_));
 sky130_fd_sc_hd__nand2_1 _5543_ (.A(_3113_),
    .B(_3156_),
    .Y(_2017_));
 sky130_fd_sc_hd__o21ai_1 _5544_ (.A1(_0900_),
    .A2(_3110_),
    .B1(_2017_),
    .Y(_2018_));
 sky130_fd_sc_hd__a221oi_1 _5545_ (.A1(_3144_),
    .A2(_3100_),
    .B1(_3149_),
    .B2(_3105_),
    .C1(_2018_),
    .Y(_2019_));
 sky130_fd_sc_hd__nand2_1 _5546_ (.A(_3127_),
    .B(_3255_),
    .Y(_2020_));
 sky130_fd_sc_hd__nand2_1 _5547_ (.A(_3132_),
    .B(_3259_),
    .Y(_2021_));
 sky130_fd_sc_hd__or2_1 _5548_ (.A(_1532_),
    .B(_3140_),
    .X(_2022_));
 sky130_fd_sc_hd__o2111a_1 _5549_ (.A1(_1776_),
    .A2(_3123_),
    .B1(_2020_),
    .C1(_2021_),
    .D1(_2022_),
    .X(_2023_));
 sky130_fd_sc_hd__nand2_1 _5550_ (.A(_3154_),
    .B(_0804_),
    .Y(_2024_));
 sky130_fd_sc_hd__nand2_1 _5551_ (.A(_3159_),
    .B(_0653_),
    .Y(_2025_));
 sky130_fd_sc_hd__nand2_1 _5552_ (.A(_2024_),
    .B(_2025_),
    .Y(_2026_));
 sky130_fd_sc_hd__a221oi_1 _5553_ (.A1(_3225_),
    .A2(_3147_),
    .B1(_3232_),
    .B2(_3151_),
    .C1(_2026_),
    .Y(_2027_));
 sky130_fd_sc_hd__and4_1 _5554_ (.A(_2016_),
    .B(_2019_),
    .C(_2023_),
    .D(_2027_),
    .X(_2028_));
 sky130_fd_sc_hd__o22ai_1 _5555_ (.A1(_0926_),
    .A2(_3175_),
    .B1(_0578_),
    .B2(_3178_),
    .Y(_2029_));
 sky130_fd_sc_hd__a221oi_1 _5556_ (.A1(_0573_),
    .A2(_3169_),
    .B1(_0581_),
    .B2(_3172_),
    .C1(_2029_),
    .Y(_2030_));
 sky130_fd_sc_hd__nand2_1 _5557_ (.A(_3191_),
    .B(_0548_),
    .Y(_2031_));
 sky130_fd_sc_hd__o21ai_1 _5558_ (.A1(_0554_),
    .A2(_3189_),
    .B1(_2031_),
    .Y(_2032_));
 sky130_fd_sc_hd__a221oi_1 _5559_ (.A1(_0552_),
    .A2(_3183_),
    .B1(_0540_),
    .B2(_3186_),
    .C1(_2032_),
    .Y(_2033_));
 sky130_fd_sc_hd__nand2_1 _5560_ (.A(_3205_),
    .B(_3047_),
    .Y(_2034_));
 sky130_fd_sc_hd__o21ai_1 _5561_ (.A1(_3216_),
    .A2(_3203_),
    .B1(_2034_),
    .Y(_2035_));
 sky130_fd_sc_hd__a221oi_1 _5562_ (.A1(_3050_),
    .A2(_3197_),
    .B1(_3053_),
    .B2(_3200_),
    .C1(_2035_),
    .Y(_2036_));
 sky130_fd_sc_hd__o22ai_1 _5563_ (.A1(_0745_),
    .A2(_3217_),
    .B1(_0568_),
    .B2(_3220_),
    .Y(_2037_));
 sky130_fd_sc_hd__a221oi_1 _5564_ (.A1(\egd_top.BitStream_buffer.BS_buffer[10] ),
    .A2(_3211_),
    .B1(\egd_top.BitStream_buffer.BS_buffer[11] ),
    .B2(_3214_),
    .C1(_2037_),
    .Y(_2038_));
 sky130_fd_sc_hd__and4_1 _5565_ (.A(_2030_),
    .B(_2033_),
    .C(_2036_),
    .D(_2038_),
    .X(_2039_));
 sky130_fd_sc_hd__o22ai_1 _5566_ (.A1(_1444_),
    .A2(_3237_),
    .B1(_3348_),
    .B2(_3240_),
    .Y(_2040_));
 sky130_fd_sc_hd__a221oi_1 _5567_ (.A1(_3345_),
    .A2(_3230_),
    .B1(_3335_),
    .B2(_3234_),
    .C1(_2040_),
    .Y(_2041_));
 sky130_fd_sc_hd__nand2_1 _5568_ (.A(_3245_),
    .B(_3290_),
    .Y(_2042_));
 sky130_fd_sc_hd__nand2_1 _5569_ (.A(_3249_),
    .B(_3282_),
    .Y(_2043_));
 sky130_fd_sc_hd__nand2_1 _5570_ (.A(_3253_),
    .B(_3286_),
    .Y(_2044_));
 sky130_fd_sc_hd__nand2_1 _5571_ (.A(_3257_),
    .B(_3278_),
    .Y(_2045_));
 sky130_fd_sc_hd__and4_1 _5572_ (.A(_2042_),
    .B(_2043_),
    .C(_2044_),
    .D(_2045_),
    .X(_2046_));
 sky130_fd_sc_hd__o22ai_1 _5573_ (.A1(_0940_),
    .A2(_3263_),
    .B1(_1069_),
    .B2(_3267_),
    .Y(_2047_));
 sky130_fd_sc_hd__a22o_1 _5574_ (.A1(_3270_),
    .A2(_3331_),
    .B1(_3273_),
    .B2(_3327_),
    .X(_2048_));
 sky130_fd_sc_hd__nor2_1 _5575_ (.A(_2047_),
    .B(_2048_),
    .Y(_2049_));
 sky130_fd_sc_hd__o22ai_1 _5576_ (.A1(_0668_),
    .A2(_3288_),
    .B1(_0819_),
    .B2(_3292_),
    .Y(_2050_));
 sky130_fd_sc_hd__a221oi_1 _5577_ (.A1(_3297_),
    .A2(_3280_),
    .B1(_3304_),
    .B2(_3284_),
    .C1(_2050_),
    .Y(_2051_));
 sky130_fd_sc_hd__and4_1 _5578_ (.A(_2041_),
    .B(_2046_),
    .C(_2049_),
    .D(_2051_),
    .X(_2052_));
 sky130_fd_sc_hd__nand2_1 _5579_ (.A(_3308_),
    .B(_3022_),
    .Y(_2053_));
 sky130_fd_sc_hd__nand2_1 _5580_ (.A(_3312_),
    .B(_3019_),
    .Y(_2054_));
 sky130_fd_sc_hd__nand2_1 _5581_ (.A(_2053_),
    .B(_2054_),
    .Y(_2055_));
 sky130_fd_sc_hd__a221oi_1 _5582_ (.A1(_3025_),
    .A2(_3302_),
    .B1(_3028_),
    .B2(_3306_),
    .C1(_2055_),
    .Y(_2056_));
 sky130_fd_sc_hd__nand2_1 _5583_ (.A(_3325_),
    .B(_0675_),
    .Y(_2057_));
 sky130_fd_sc_hd__nand2_1 _5584_ (.A(_3329_),
    .B(_0674_),
    .Y(_2058_));
 sky130_fd_sc_hd__nand2_1 _5585_ (.A(_2057_),
    .B(_2058_),
    .Y(_2059_));
 sky130_fd_sc_hd__a221oi_1 _5586_ (.A1(_3353_),
    .A2(_3320_),
    .B1(_3357_),
    .B2(_3323_),
    .C1(_2059_),
    .Y(_2060_));
 sky130_fd_sc_hd__nand2_1 _5587_ (.A(_3339_),
    .B(_2998_),
    .Y(_2061_));
 sky130_fd_sc_hd__nand2_1 _5588_ (.A(_3343_),
    .B(_3013_),
    .Y(_2062_));
 sky130_fd_sc_hd__or2_1 _5589_ (.A(_0634_),
    .B(_3349_),
    .X(_2063_));
 sky130_fd_sc_hd__o2111a_1 _5590_ (.A1(_0922_),
    .A2(_3337_),
    .B1(_2061_),
    .C1(_2062_),
    .D1(_2063_),
    .X(_2064_));
 sky130_fd_sc_hd__nand2_1 _5591_ (.A(_3364_),
    .B(_3037_),
    .Y(_2065_));
 sky130_fd_sc_hd__o21ai_1 _5592_ (.A1(_3188_),
    .A2(_3362_),
    .B1(_2065_),
    .Y(_2066_));
 sky130_fd_sc_hd__a221oi_1 _5593_ (.A1(_3031_),
    .A2(_3355_),
    .B1(_3034_),
    .B2(_3359_),
    .C1(_2066_),
    .Y(_2067_));
 sky130_fd_sc_hd__and4_1 _5594_ (.A(_2056_),
    .B(_2060_),
    .C(_2064_),
    .D(_2067_),
    .X(_2068_));
 sky130_fd_sc_hd__and4_1 _5595_ (.A(_2028_),
    .B(_2039_),
    .C(_2052_),
    .D(_2068_),
    .X(_2069_));
 sky130_fd_sc_hd__nand2_1 _5596_ (.A(_0333_),
    .B(_0703_),
    .Y(_2070_));
 sky130_fd_sc_hd__nand2_1 _5597_ (.A(_0337_),
    .B(_0404_),
    .Y(_2071_));
 sky130_fd_sc_hd__nand2_1 _5598_ (.A(_2070_),
    .B(_2071_),
    .Y(_2072_));
 sky130_fd_sc_hd__a221oi_1 _5599_ (.A1(_0400_),
    .A2(_0327_),
    .B1(_0701_),
    .B2(_0331_),
    .C1(_2072_),
    .Y(_2073_));
 sky130_fd_sc_hd__o22ai_1 _5600_ (.A1(_0438_),
    .A2(_0344_),
    .B1(_0714_),
    .B2(_0348_),
    .Y(_2074_));
 sky130_fd_sc_hd__a22o_1 _5601_ (.A1(_0351_),
    .A2(_0429_),
    .B1(_0354_),
    .B2(_0433_),
    .X(_2075_));
 sky130_fd_sc_hd__nor2_1 _5602_ (.A(_2074_),
    .B(_2075_),
    .Y(_2076_));
 sky130_fd_sc_hd__nand2_1 _5603_ (.A(_0370_),
    .B(_0695_),
    .Y(_2077_));
 sky130_fd_sc_hd__o21ai_1 _5604_ (.A1(_1714_),
    .A2(_0368_),
    .B1(_2077_),
    .Y(_2078_));
 sky130_fd_sc_hd__a221oi_1 _5605_ (.A1(_0376_),
    .A2(_0361_),
    .B1(_0380_),
    .B2(_0365_),
    .C1(_2078_),
    .Y(_2079_));
 sky130_fd_sc_hd__nand2_1 _5606_ (.A(_0387_),
    .B(_0421_),
    .Y(_2080_));
 sky130_fd_sc_hd__o21ai_1 _5607_ (.A1(_0412_),
    .A2(_0385_),
    .B1(_2080_),
    .Y(_2081_));
 sky130_fd_sc_hd__a221oi_1 _5608_ (.A1(_0417_),
    .A2(_0378_),
    .B1(_0423_),
    .B2(_0382_),
    .C1(_2081_),
    .Y(_2082_));
 sky130_fd_sc_hd__and4_1 _5609_ (.A(_2073_),
    .B(_2076_),
    .C(_2079_),
    .D(_2082_),
    .X(_2083_));
 sky130_fd_sc_hd__nand2_1 _5610_ (.A(_0398_),
    .B(_3095_),
    .Y(_2084_));
 sky130_fd_sc_hd__nand2_1 _5611_ (.A(_0402_),
    .B(_3107_),
    .Y(_2085_));
 sky130_fd_sc_hd__or2_1 _5612_ (.A(_0903_),
    .B(_0407_),
    .X(_2086_));
 sky130_fd_sc_hd__o2111a_1 _5613_ (.A1(_0614_),
    .A2(_0396_),
    .B1(_2084_),
    .C1(_2085_),
    .D1(_2086_),
    .X(_2087_));
 sky130_fd_sc_hd__nand2_1 _5614_ (.A(_0415_),
    .B(_3129_),
    .Y(_2088_));
 sky130_fd_sc_hd__nand2_1 _5615_ (.A(_0419_),
    .B(_3134_),
    .Y(_2089_));
 sky130_fd_sc_hd__or2_1 _5616_ (.A(_3137_),
    .B(_0425_),
    .X(_2090_));
 sky130_fd_sc_hd__o2111a_1 _5617_ (.A1(_3120_),
    .A2(_0413_),
    .B1(_2088_),
    .C1(_2089_),
    .D1(_2090_),
    .X(_2091_));
 sky130_fd_sc_hd__nand2_1 _5618_ (.A(_0441_),
    .B(_0451_),
    .Y(_2092_));
 sky130_fd_sc_hd__o21ai_1 _5619_ (.A1(_0708_),
    .A2(_0439_),
    .B1(_2092_),
    .Y(_2093_));
 sky130_fd_sc_hd__a221oi_1 _5620_ (.A1(_0461_),
    .A2(_0431_),
    .B1(_0455_),
    .B2(_0435_),
    .C1(_2093_),
    .Y(_2094_));
 sky130_fd_sc_hd__nand2_1 _5621_ (.A(_0459_),
    .B(_3057_),
    .Y(_2095_));
 sky130_fd_sc_hd__o21ai_1 _5622_ (.A1(_0764_),
    .A2(_0457_),
    .B1(_2095_),
    .Y(_2096_));
 sky130_fd_sc_hd__a221oi_1 _5623_ (.A1(_3076_),
    .A2(_0449_),
    .B1(_3085_),
    .B2(_0453_),
    .C1(_2096_),
    .Y(_2097_));
 sky130_fd_sc_hd__and4_1 _5624_ (.A(_2087_),
    .B(_2091_),
    .C(_2094_),
    .D(_2097_),
    .X(_2098_));
 sky130_fd_sc_hd__and2_1 _5625_ (.A(_2083_),
    .B(_2098_),
    .X(_2099_));
 sky130_fd_sc_hd__nand2_1 _5626_ (.A(_0473_),
    .B(_0346_),
    .Y(_2100_));
 sky130_fd_sc_hd__a22o_1 _5627_ (.A1(_0477_),
    .A2(_0353_),
    .B1(_0480_),
    .B2(_0356_),
    .X(_2101_));
 sky130_fd_sc_hd__inv_2 _5628_ (.A(_2101_),
    .Y(_2102_));
 sky130_fd_sc_hd__o211a_1 _5629_ (.A1(_0343_),
    .A2(_0471_),
    .B1(_2100_),
    .C1(_2102_),
    .X(_2103_));
 sky130_fd_sc_hd__nand2_1 _5630_ (.A(_0497_),
    .B(_0525_),
    .Y(_2104_));
 sky130_fd_sc_hd__o21ai_1 _5631_ (.A1(_1373_),
    .A2(_0495_),
    .B1(_2104_),
    .Y(_2105_));
 sky130_fd_sc_hd__a221oi_1 _5632_ (.A1(_0535_),
    .A2(_0487_),
    .B1(_0531_),
    .B2(_0491_),
    .C1(_2105_),
    .Y(_2106_));
 sky130_fd_sc_hd__nand2_1 _5633_ (.A(_0507_),
    .B(_0689_),
    .Y(_2107_));
 sky130_fd_sc_hd__nand2_1 _5634_ (.A(_0511_),
    .B(_0359_),
    .Y(_2108_));
 sky130_fd_sc_hd__or2_1 _5635_ (.A(_1741_),
    .B(_0517_),
    .X(_2109_));
 sky130_fd_sc_hd__o2111a_1 _5636_ (.A1(_0690_),
    .A2(_0505_),
    .B1(_2107_),
    .C1(_2108_),
    .D1(_2109_),
    .X(_2110_));
 sky130_fd_sc_hd__nand2_1 _5637_ (.A(_0529_),
    .B(_0335_),
    .Y(_2111_));
 sky130_fd_sc_hd__nand2_1 _5638_ (.A(_0533_),
    .B(_0339_),
    .Y(_2112_));
 sky130_fd_sc_hd__nand2_1 _5639_ (.A(_2111_),
    .B(_2112_),
    .Y(_2113_));
 sky130_fd_sc_hd__a221oi_1 _5640_ (.A1(_0323_),
    .A2(_0523_),
    .B1(_0329_),
    .B2(_0527_),
    .C1(_2113_),
    .Y(_2114_));
 sky130_fd_sc_hd__and4_1 _5641_ (.A(_2103_),
    .B(_2106_),
    .C(_2110_),
    .D(_2114_),
    .X(_2115_));
 sky130_fd_sc_hd__nand2_1 _5642_ (.A(_0546_),
    .B(_0493_),
    .Y(_2116_));
 sky130_fd_sc_hd__nand2_1 _5643_ (.A(_0550_),
    .B(\egd_top.BitStream_buffer.BS_buffer[16] ),
    .Y(_2117_));
 sky130_fd_sc_hd__or2_1 _5644_ (.A(_0728_),
    .B(_0555_),
    .X(_2118_));
 sky130_fd_sc_hd__o2111a_1 _5645_ (.A1(_1150_),
    .A2(_0544_),
    .B1(_2116_),
    .C1(_2117_),
    .D1(_2118_),
    .X(_2119_));
 sky130_fd_sc_hd__nand2_1 _5646_ (.A(_0562_),
    .B(_0509_),
    .Y(_2120_));
 sky130_fd_sc_hd__nand2_1 _5647_ (.A(_0565_),
    .B(_0513_),
    .Y(_2121_));
 sky130_fd_sc_hd__or2_1 _5648_ (.A(_0516_),
    .B(_0569_),
    .X(_2122_));
 sky130_fd_sc_hd__o2111a_1 _5649_ (.A1(_0504_),
    .A2(_0560_),
    .B1(_2120_),
    .C1(_2121_),
    .D1(_2122_),
    .X(_2123_));
 sky130_fd_sc_hd__or2_1 _5650_ (.A(_0890_),
    .B(_0583_),
    .X(_2124_));
 sky130_fd_sc_hd__o221a_1 _5651_ (.A1(_0756_),
    .A2(_0575_),
    .B1(_0596_),
    .B2(_0579_),
    .C1(_2124_),
    .X(_2125_));
 sky130_fd_sc_hd__o22ai_1 _5652_ (.A1(_0468_),
    .A2(_0594_),
    .B1(_0723_),
    .B2(_0597_),
    .Y(_2126_));
 sky130_fd_sc_hd__a221oi_1 _5653_ (.A1(_0479_),
    .A2(_0588_),
    .B1(_0482_),
    .B2(_0591_),
    .C1(_2126_),
    .Y(_2127_));
 sky130_fd_sc_hd__and4_1 _5654_ (.A(_2119_),
    .B(_2123_),
    .C(_2125_),
    .D(_2127_),
    .X(_2128_));
 sky130_fd_sc_hd__and3_1 _5655_ (.A(_2099_),
    .B(_2115_),
    .C(_2128_),
    .X(_2129_));
 sky130_fd_sc_hd__nand2_1 _5656_ (.A(_0605_),
    .B(\egd_top.BitStream_buffer.BS_buffer[12] ),
    .Y(_2130_));
 sky130_fd_sc_hd__nand3_2 _5657_ (.A(_2069_),
    .B(_2129_),
    .C(_2130_),
    .Y(_2131_));
 sky130_fd_sc_hd__inv_2 _5658_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[3] ),
    .Y(_2132_));
 sky130_fd_sc_hd__a21oi_1 _5659_ (.A1(_2132_),
    .A2(_2996_),
    .B1(_2937_),
    .Y(_2133_));
 sky130_fd_sc_hd__o21a_1 _5660_ (.A1(_0898_),
    .A2(_2131_),
    .B1(_2133_),
    .X(_0285_));
 sky130_fd_sc_hd__o22ai_1 _5661_ (.A1(_3266_),
    .A2(_3083_),
    .B1(_0651_),
    .B2(_3091_),
    .Y(_2134_));
 sky130_fd_sc_hd__a221oi_1 _5662_ (.A1(_3275_),
    .A2(_3067_),
    .B1(_0653_),
    .B2(_3074_),
    .C1(_2134_),
    .Y(_2135_));
 sky130_fd_sc_hd__nand2_1 _5663_ (.A(_3113_),
    .B(_3144_),
    .Y(_2136_));
 sky130_fd_sc_hd__o21ai_1 _5664_ (.A1(_1031_),
    .A2(_3110_),
    .B1(_2136_),
    .Y(_2137_));
 sky130_fd_sc_hd__a221oi_1 _5665_ (.A1(_3149_),
    .A2(_3100_),
    .B1(_3255_),
    .B2(_3105_),
    .C1(_2137_),
    .Y(_2138_));
 sky130_fd_sc_hd__nand2_1 _5666_ (.A(_3127_),
    .B(_3247_),
    .Y(_2139_));
 sky130_fd_sc_hd__nand2_1 _5667_ (.A(_3132_),
    .B(_3251_),
    .Y(_2140_));
 sky130_fd_sc_hd__or2_1 _5668_ (.A(_1654_),
    .B(_3140_),
    .X(_2141_));
 sky130_fd_sc_hd__o2111a_1 _5669_ (.A1(_3262_),
    .A2(_3123_),
    .B1(_2139_),
    .C1(_2140_),
    .D1(_2141_),
    .X(_2142_));
 sky130_fd_sc_hd__nand2_1 _5670_ (.A(_3154_),
    .B(_3225_),
    .Y(_2143_));
 sky130_fd_sc_hd__nand2_1 _5671_ (.A(_3159_),
    .B(_0804_),
    .Y(_2144_));
 sky130_fd_sc_hd__nand2_1 _5672_ (.A(_2143_),
    .B(_2144_),
    .Y(_2145_));
 sky130_fd_sc_hd__a221oi_2 _5673_ (.A1(_3232_),
    .A2(_3147_),
    .B1(_3286_),
    .B2(_3151_),
    .C1(_2145_),
    .Y(_2146_));
 sky130_fd_sc_hd__and4_1 _5674_ (.A(_2135_),
    .B(_2138_),
    .C(_2142_),
    .D(_2146_),
    .X(_2147_));
 sky130_fd_sc_hd__o22ai_1 _5675_ (.A1(_0578_),
    .A2(_3175_),
    .B1(_0574_),
    .B2(_3178_),
    .Y(_2148_));
 sky130_fd_sc_hd__a221oi_1 _5676_ (.A1(_0581_),
    .A2(_3169_),
    .B1(_0552_),
    .B2(_3172_),
    .C1(_2148_),
    .Y(_2149_));
 sky130_fd_sc_hd__nand2_1 _5677_ (.A(_3191_),
    .B(\egd_top.BitStream_buffer.BS_buffer[7] ),
    .Y(_2150_));
 sky130_fd_sc_hd__o21ai_1 _5678_ (.A1(_0745_),
    .A2(_3189_),
    .B1(_2150_),
    .Y(_2151_));
 sky130_fd_sc_hd__a221oi_1 _5679_ (.A1(_0540_),
    .A2(_3183_),
    .B1(_0548_),
    .B2(_3186_),
    .C1(_2151_),
    .Y(_2152_));
 sky130_fd_sc_hd__nand2_1 _5680_ (.A(_3205_),
    .B(_3050_),
    .Y(_2153_));
 sky130_fd_sc_hd__o21ai_1 _5681_ (.A1(_3219_),
    .A2(_3203_),
    .B1(_2153_),
    .Y(_2154_));
 sky130_fd_sc_hd__a221oi_1 _5682_ (.A1(_3053_),
    .A2(_3197_),
    .B1(_0607_),
    .B2(_3200_),
    .C1(_2154_),
    .Y(_2155_));
 sky130_fd_sc_hd__o22ai_1 _5683_ (.A1(_0568_),
    .A2(_3217_),
    .B1(_0750_),
    .B2(_3220_),
    .Y(_2156_));
 sky130_fd_sc_hd__a221oi_1 _5684_ (.A1(\egd_top.BitStream_buffer.BS_buffer[11] ),
    .A2(_3211_),
    .B1(\egd_top.BitStream_buffer.BS_buffer[12] ),
    .B2(_3214_),
    .C1(_2156_),
    .Y(_2157_));
 sky130_fd_sc_hd__and4_1 _5685_ (.A(_2149_),
    .B(_2152_),
    .C(_2155_),
    .D(_2157_),
    .X(_2158_));
 sky130_fd_sc_hd__o22ai_1 _5686_ (.A1(_3348_),
    .A2(_3237_),
    .B1(_0671_),
    .B2(_3240_),
    .Y(_2159_));
 sky130_fd_sc_hd__a221oi_1 _5687_ (.A1(_3335_),
    .A2(_3230_),
    .B1(_3314_),
    .B2(_3234_),
    .C1(_2159_),
    .Y(_2160_));
 sky130_fd_sc_hd__nand2_1 _5688_ (.A(_3245_),
    .B(_3278_),
    .Y(_2161_));
 sky130_fd_sc_hd__nand2_1 _5689_ (.A(_3249_),
    .B(_3318_),
    .Y(_2162_));
 sky130_fd_sc_hd__nand2_1 _5690_ (.A(_3253_),
    .B(_3290_),
    .Y(_2163_));
 sky130_fd_sc_hd__nand2_1 _5691_ (.A(_3257_),
    .B(_3282_),
    .Y(_2164_));
 sky130_fd_sc_hd__and4_1 _5692_ (.A(_2161_),
    .B(_2162_),
    .C(_2163_),
    .D(_2164_),
    .X(_2165_));
 sky130_fd_sc_hd__o22ai_1 _5693_ (.A1(_1069_),
    .A2(_3263_),
    .B1(_1196_),
    .B2(_3267_),
    .Y(_2166_));
 sky130_fd_sc_hd__a22o_1 _5694_ (.A1(_3270_),
    .A2(_3327_),
    .B1(_3273_),
    .B2(_3341_),
    .X(_2167_));
 sky130_fd_sc_hd__nor2_1 _5695_ (.A(_2166_),
    .B(_2167_),
    .Y(_2168_));
 sky130_fd_sc_hd__o22ai_1 _5696_ (.A1(_0819_),
    .A2(_3288_),
    .B1(_0952_),
    .B2(_3292_),
    .Y(_2169_));
 sky130_fd_sc_hd__a221oi_1 _5697_ (.A1(_3304_),
    .A2(_3280_),
    .B1(_3353_),
    .B2(_3284_),
    .C1(_2169_),
    .Y(_2170_));
 sky130_fd_sc_hd__and4_1 _5698_ (.A(_2160_),
    .B(_2165_),
    .C(_2168_),
    .D(_2170_),
    .X(_2171_));
 sky130_fd_sc_hd__nand2_1 _5699_ (.A(_3308_),
    .B(_3025_),
    .Y(_2172_));
 sky130_fd_sc_hd__nand2_1 _5700_ (.A(_3312_),
    .B(_3022_),
    .Y(_2173_));
 sky130_fd_sc_hd__nand2_1 _5701_ (.A(_2172_),
    .B(_2173_),
    .Y(_2174_));
 sky130_fd_sc_hd__a221oi_1 _5702_ (.A1(_3028_),
    .A2(_3302_),
    .B1(_3031_),
    .B2(_3306_),
    .C1(_2174_),
    .Y(_2175_));
 sky130_fd_sc_hd__nand2_1 _5703_ (.A(_3325_),
    .B(_2998_),
    .Y(_2176_));
 sky130_fd_sc_hd__nand2_1 _5704_ (.A(_3329_),
    .B(_0675_),
    .Y(_2177_));
 sky130_fd_sc_hd__nand2_1 _5705_ (.A(_2176_),
    .B(_2177_),
    .Y(_2178_));
 sky130_fd_sc_hd__a221oi_1 _5706_ (.A1(_3357_),
    .A2(_3320_),
    .B1(_0674_),
    .B2(_3323_),
    .C1(_2178_),
    .Y(_2179_));
 sky130_fd_sc_hd__nand2_1 _5707_ (.A(_3339_),
    .B(_3010_),
    .Y(_2180_));
 sky130_fd_sc_hd__nand2_1 _5708_ (.A(_3343_),
    .B(_3016_),
    .Y(_2181_));
 sky130_fd_sc_hd__or2_1 _5709_ (.A(_0786_),
    .B(_3349_),
    .X(_2182_));
 sky130_fd_sc_hd__o2111a_1 _5710_ (.A1(_3174_),
    .A2(_3337_),
    .B1(_2180_),
    .C1(_2181_),
    .D1(_2182_),
    .X(_2183_));
 sky130_fd_sc_hd__nand2_1 _5711_ (.A(_3364_),
    .B(_3040_),
    .Y(_2184_));
 sky130_fd_sc_hd__o21ai_1 _5712_ (.A1(_3216_),
    .A2(_3362_),
    .B1(_2184_),
    .Y(_2185_));
 sky130_fd_sc_hd__a221oi_1 _5713_ (.A1(_3034_),
    .A2(_3355_),
    .B1(_3037_),
    .B2(_3359_),
    .C1(_2185_),
    .Y(_2186_));
 sky130_fd_sc_hd__and4_1 _5714_ (.A(_2175_),
    .B(_2179_),
    .C(_2183_),
    .D(_2186_),
    .X(_2187_));
 sky130_fd_sc_hd__and4_1 _5715_ (.A(_2147_),
    .B(_2158_),
    .C(_2171_),
    .D(_2187_),
    .X(_2188_));
 sky130_fd_sc_hd__nand2_1 _5716_ (.A(_0333_),
    .B(_0400_),
    .Y(_2189_));
 sky130_fd_sc_hd__nand2_1 _5717_ (.A(_0337_),
    .B(_0703_),
    .Y(_2190_));
 sky130_fd_sc_hd__nand2_1 _5718_ (.A(_2189_),
    .B(_2190_),
    .Y(_2191_));
 sky130_fd_sc_hd__a221oi_1 _5719_ (.A1(_0701_),
    .A2(_0327_),
    .B1(_0417_),
    .B2(_0331_),
    .C1(_2191_),
    .Y(_2192_));
 sky130_fd_sc_hd__o22ai_1 _5720_ (.A1(_0714_),
    .A2(_0344_),
    .B1(_0853_),
    .B2(_0348_),
    .Y(_2193_));
 sky130_fd_sc_hd__a22o_1 _5721_ (.A1(_0351_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[51] ),
    .B1(_0354_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[52] ),
    .X(_2194_));
 sky130_fd_sc_hd__nor2_1 _5722_ (.A(_2193_),
    .B(_2194_),
    .Y(_2195_));
 sky130_fd_sc_hd__nand2_1 _5723_ (.A(_0370_),
    .B(_0437_),
    .Y(_2196_));
 sky130_fd_sc_hd__o21ai_1 _5724_ (.A1(_0384_),
    .A2(_0368_),
    .B1(_2196_),
    .Y(_2197_));
 sky130_fd_sc_hd__a221oi_1 _5725_ (.A1(_0380_),
    .A2(_0361_),
    .B1(_0389_),
    .B2(_0365_),
    .C1(_2197_),
    .Y(_2198_));
 sky130_fd_sc_hd__nand2_1 _5726_ (.A(_0387_),
    .B(_0411_),
    .Y(_2199_));
 sky130_fd_sc_hd__o21ai_1 _5727_ (.A1(_0708_),
    .A2(_0385_),
    .B1(_2199_),
    .Y(_2200_));
 sky130_fd_sc_hd__a221oi_1 _5728_ (.A1(_0423_),
    .A2(_0378_),
    .B1(_0421_),
    .B2(_0382_),
    .C1(_2200_),
    .Y(_2201_));
 sky130_fd_sc_hd__and4_1 _5729_ (.A(_2192_),
    .B(_2195_),
    .C(_2198_),
    .D(_2201_),
    .X(_2202_));
 sky130_fd_sc_hd__nand2_1 _5730_ (.A(_0398_),
    .B(_3102_),
    .Y(_2203_));
 sky130_fd_sc_hd__nand2_1 _5731_ (.A(_0402_),
    .B(_3115_),
    .Y(_2204_));
 sky130_fd_sc_hd__or2_1 _5732_ (.A(_1034_),
    .B(_0407_),
    .X(_2205_));
 sky130_fd_sc_hd__o2111a_1 _5733_ (.A1(_0767_),
    .A2(_0396_),
    .B1(_2203_),
    .C1(_2204_),
    .D1(_2205_),
    .X(_2206_));
 sky130_fd_sc_hd__nand2_1 _5734_ (.A(_0415_),
    .B(_3136_),
    .Y(_2207_));
 sky130_fd_sc_hd__nand2_1 _5735_ (.A(_0419_),
    .B(_3119_),
    .Y(_2208_));
 sky130_fd_sc_hd__or2_1 _5736_ (.A(_0620_),
    .B(_0425_),
    .X(_2209_));
 sky130_fd_sc_hd__o2111a_1 _5737_ (.A1(_3077_),
    .A2(_0413_),
    .B1(_2207_),
    .C1(_2208_),
    .D1(_2209_),
    .X(_2210_));
 sky130_fd_sc_hd__nand2_1 _5738_ (.A(_0441_),
    .B(_0461_),
    .Y(_2211_));
 sky130_fd_sc_hd__o21ai_1 _5739_ (.A1(_0848_),
    .A2(_0439_),
    .B1(_2211_),
    .Y(_2212_));
 sky130_fd_sc_hd__a221oi_1 _5740_ (.A1(_0455_),
    .A2(_0431_),
    .B1(_3107_),
    .B2(_0435_),
    .C1(_2212_),
    .Y(_2213_));
 sky130_fd_sc_hd__nand2_1 _5741_ (.A(_0459_),
    .B(_3069_),
    .Y(_2214_));
 sky130_fd_sc_hd__o21ai_1 _5742_ (.A1(_0900_),
    .A2(_0457_),
    .B1(_2214_),
    .Y(_2215_));
 sky130_fd_sc_hd__a221oi_1 _5743_ (.A1(_3085_),
    .A2(_0449_),
    .B1(_3057_),
    .B2(_0453_),
    .C1(_2215_),
    .Y(_2216_));
 sky130_fd_sc_hd__and4_1 _5744_ (.A(_2206_),
    .B(_2210_),
    .C(_2213_),
    .D(_2216_),
    .X(_2217_));
 sky130_fd_sc_hd__and2_1 _5745_ (.A(_2202_),
    .B(_2217_),
    .X(_2218_));
 sky130_fd_sc_hd__nand2_1 _5746_ (.A(_0473_),
    .B(_0353_),
    .Y(_2219_));
 sky130_fd_sc_hd__a22o_1 _5747_ (.A1(_0477_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[39] ),
    .B1(_0480_),
    .B2(_0339_),
    .X(_2220_));
 sky130_fd_sc_hd__inv_2 _5748_ (.A(_2220_),
    .Y(_2221_));
 sky130_fd_sc_hd__o211a_1 _5749_ (.A1(_0347_),
    .A2(_0471_),
    .B1(_2219_),
    .C1(_2221_),
    .X(_2222_));
 sky130_fd_sc_hd__nand2_1 _5750_ (.A(_0497_),
    .B(_0359_),
    .Y(_2223_));
 sky130_fd_sc_hd__o21ai_1 _5751_ (.A1(_1497_),
    .A2(_0495_),
    .B1(_2223_),
    .Y(_2224_));
 sky130_fd_sc_hd__a221oi_1 _5752_ (.A1(_0531_),
    .A2(_0487_),
    .B1(_0521_),
    .B2(_0491_),
    .C1(_2224_),
    .Y(_2225_));
 sky130_fd_sc_hd__nand2_1 _5753_ (.A(_0507_),
    .B(_0372_),
    .Y(_2226_));
 sky130_fd_sc_hd__nand2_1 _5754_ (.A(_0511_),
    .B(_0363_),
    .Y(_2227_));
 sky130_fd_sc_hd__or2_1 _5755_ (.A(_0367_),
    .B(_0517_),
    .X(_2228_));
 sky130_fd_sc_hd__o2111a_1 _5756_ (.A1(_0343_),
    .A2(_0505_),
    .B1(_2226_),
    .C1(_2227_),
    .D1(_2228_),
    .X(_2229_));
 sky130_fd_sc_hd__nand2_1 _5757_ (.A(_0529_),
    .B(_0323_),
    .Y(_2230_));
 sky130_fd_sc_hd__nand2_1 _5758_ (.A(_0533_),
    .B(_0335_),
    .Y(_2231_));
 sky130_fd_sc_hd__nand2_1 _5759_ (.A(_2230_),
    .B(_2231_),
    .Y(_2232_));
 sky130_fd_sc_hd__a221oi_1 _5760_ (.A1(_0329_),
    .A2(_0523_),
    .B1(_0376_),
    .B2(_0527_),
    .C1(_2232_),
    .Y(_2233_));
 sky130_fd_sc_hd__and4_1 _5761_ (.A(_2222_),
    .B(_2225_),
    .C(_2229_),
    .D(_2233_),
    .X(_2234_));
 sky130_fd_sc_hd__nand2_1 _5762_ (.A(_0546_),
    .B(_0499_),
    .Y(_2235_));
 sky130_fd_sc_hd__nand2_1 _5763_ (.A(_0550_),
    .B(_0489_),
    .Y(_2236_));
 sky130_fd_sc_hd__or2_1 _5764_ (.A(_0867_),
    .B(_0555_),
    .X(_2237_));
 sky130_fd_sc_hd__o2111a_1 _5765_ (.A1(_0494_),
    .A2(_0544_),
    .B1(_2235_),
    .C1(_2236_),
    .D1(_2237_),
    .X(_2238_));
 sky130_fd_sc_hd__nand2_1 _5766_ (.A(_0562_),
    .B(_0503_),
    .Y(_2239_));
 sky130_fd_sc_hd__nand2_1 _5767_ (.A(_0565_),
    .B(_0515_),
    .Y(_2240_));
 sky130_fd_sc_hd__or2_1 _5768_ (.A(_0734_),
    .B(_0569_),
    .X(_2241_));
 sky130_fd_sc_hd__o2111a_1 _5769_ (.A1(_0468_),
    .A2(_0560_),
    .B1(_2239_),
    .C1(_2240_),
    .D1(_2241_),
    .X(_2242_));
 sky130_fd_sc_hd__or2_1 _5770_ (.A(_1022_),
    .B(_0583_),
    .X(_2243_));
 sky130_fd_sc_hd__o221a_1 _5771_ (.A1(_0890_),
    .A2(_0575_),
    .B1(_0756_),
    .B2(_0579_),
    .C1(_2243_),
    .X(_2244_));
 sky130_fd_sc_hd__o22ai_1 _5772_ (.A1(_0723_),
    .A2(_0594_),
    .B1(_0862_),
    .B2(_0597_),
    .Y(_2245_));
 sky130_fd_sc_hd__a221oi_1 _5773_ (.A1(_0482_),
    .A2(_0588_),
    .B1(_0535_),
    .B2(_0591_),
    .C1(_2245_),
    .Y(_2246_));
 sky130_fd_sc_hd__and4_1 _5774_ (.A(_2238_),
    .B(_2242_),
    .C(_2244_),
    .D(_2246_),
    .X(_2247_));
 sky130_fd_sc_hd__and3_1 _5775_ (.A(_2218_),
    .B(_2234_),
    .C(_2247_),
    .X(_2248_));
 sky130_fd_sc_hd__nand2_1 _5776_ (.A(_0605_),
    .B(\egd_top.BitStream_buffer.BS_buffer[13] ),
    .Y(_2249_));
 sky130_fd_sc_hd__nand3_2 _5777_ (.A(_2188_),
    .B(_2248_),
    .C(_2249_),
    .Y(_2250_));
 sky130_fd_sc_hd__inv_2 _5778_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[2] ),
    .Y(_2251_));
 sky130_fd_sc_hd__a21oi_1 _5779_ (.A1(_2251_),
    .A2(_2996_),
    .B1(_2937_),
    .Y(_2252_));
 sky130_fd_sc_hd__o21a_1 _5780_ (.A1(_0898_),
    .A2(_2250_),
    .B1(_2252_),
    .X(_0284_));
 sky130_fd_sc_hd__o22ai_1 _5781_ (.A1(_0651_),
    .A2(_3083_),
    .B1(_0802_),
    .B2(_3091_),
    .Y(_2253_));
 sky130_fd_sc_hd__a221oi_1 _5782_ (.A1(_0653_),
    .A2(_3067_),
    .B1(_0804_),
    .B2(_3074_),
    .C1(_2253_),
    .Y(_2254_));
 sky130_fd_sc_hd__nand2_1 _5783_ (.A(_3113_),
    .B(_3149_),
    .Y(_2255_));
 sky130_fd_sc_hd__o21ai_1 _5784_ (.A1(_1159_),
    .A2(_3110_),
    .B1(_2255_),
    .Y(_2256_));
 sky130_fd_sc_hd__a221oi_1 _5785_ (.A1(_3255_),
    .A2(_3100_),
    .B1(_3247_),
    .B2(_3105_),
    .C1(_2256_),
    .Y(_2257_));
 sky130_fd_sc_hd__nand2_1 _5786_ (.A(_3127_),
    .B(_3259_),
    .Y(_2258_));
 sky130_fd_sc_hd__nand2_1 _5787_ (.A(_3132_),
    .B(_0646_),
    .Y(_2259_));
 sky130_fd_sc_hd__or2_1 _5788_ (.A(_1776_),
    .B(_3140_),
    .X(_2260_));
 sky130_fd_sc_hd__o2111a_1 _5789_ (.A1(_3266_),
    .A2(_3123_),
    .B1(_2258_),
    .C1(_2259_),
    .D1(_2260_),
    .X(_2261_));
 sky130_fd_sc_hd__nand2_1 _5790_ (.A(_3154_),
    .B(_3232_),
    .Y(_2262_));
 sky130_fd_sc_hd__nand2_1 _5791_ (.A(_3159_),
    .B(_3225_),
    .Y(_2263_));
 sky130_fd_sc_hd__nand2_1 _5792_ (.A(_2262_),
    .B(_2263_),
    .Y(_2264_));
 sky130_fd_sc_hd__a221oi_1 _5793_ (.A1(_3286_),
    .A2(_3147_),
    .B1(_3290_),
    .B2(_3151_),
    .C1(_2264_),
    .Y(_2265_));
 sky130_fd_sc_hd__and4_1 _5794_ (.A(_2254_),
    .B(_2257_),
    .C(_2261_),
    .D(_2265_),
    .X(_2266_));
 sky130_fd_sc_hd__o22ai_1 _5795_ (.A1(_0574_),
    .A2(_3175_),
    .B1(_0582_),
    .B2(_3178_),
    .Y(_2267_));
 sky130_fd_sc_hd__a221oi_1 _5796_ (.A1(_0552_),
    .A2(_3169_),
    .B1(_0540_),
    .B2(_3172_),
    .C1(_2267_),
    .Y(_2268_));
 sky130_fd_sc_hd__nand2_1 _5797_ (.A(_3191_),
    .B(\egd_top.BitStream_buffer.BS_buffer[8] ),
    .Y(_2269_));
 sky130_fd_sc_hd__o21ai_1 _5798_ (.A1(_0568_),
    .A2(_3189_),
    .B1(_2269_),
    .Y(_2270_));
 sky130_fd_sc_hd__a221oi_1 _5799_ (.A1(_0548_),
    .A2(_3183_),
    .B1(\egd_top.BitStream_buffer.BS_buffer[7] ),
    .B2(_3186_),
    .C1(_2270_),
    .Y(_2271_));
 sky130_fd_sc_hd__nand2_1 _5800_ (.A(_3205_),
    .B(_3053_),
    .Y(_2272_));
 sky130_fd_sc_hd__o21ai_1 _5801_ (.A1(_0638_),
    .A2(_3203_),
    .B1(_2272_),
    .Y(_2273_));
 sky130_fd_sc_hd__a221oi_1 _5802_ (.A1(_0607_),
    .A2(_3197_),
    .B1(_0577_),
    .B2(_3200_),
    .C1(_2273_),
    .Y(_2274_));
 sky130_fd_sc_hd__o22ai_1 _5803_ (.A1(_0750_),
    .A2(_3217_),
    .B1(_0559_),
    .B2(_3220_),
    .Y(_2275_));
 sky130_fd_sc_hd__a221oi_1 _5804_ (.A1(\egd_top.BitStream_buffer.BS_buffer[12] ),
    .A2(_3211_),
    .B1(\egd_top.BitStream_buffer.BS_buffer[13] ),
    .B2(_3214_),
    .C1(_2275_),
    .Y(_2276_));
 sky130_fd_sc_hd__and4_1 _5805_ (.A(_2268_),
    .B(_2271_),
    .C(_2274_),
    .D(_2276_),
    .X(_2277_));
 sky130_fd_sc_hd__o22ai_1 _5806_ (.A1(_0671_),
    .A2(_3237_),
    .B1(_3336_),
    .B2(_3240_),
    .Y(_2278_));
 sky130_fd_sc_hd__a221oi_1 _5807_ (.A1(_3314_),
    .A2(_3230_),
    .B1(_3310_),
    .B2(_3234_),
    .C1(_2278_),
    .Y(_2279_));
 sky130_fd_sc_hd__nand2_1 _5808_ (.A(_3245_),
    .B(_3282_),
    .Y(_2280_));
 sky130_fd_sc_hd__nand2_1 _5809_ (.A(_3249_),
    .B(_3322_),
    .Y(_2281_));
 sky130_fd_sc_hd__nand2_1 _5810_ (.A(_3253_),
    .B(_3278_),
    .Y(_2282_));
 sky130_fd_sc_hd__nand2_1 _5811_ (.A(_3257_),
    .B(_3318_),
    .Y(_2283_));
 sky130_fd_sc_hd__and4_1 _5812_ (.A(_2280_),
    .B(_2281_),
    .C(_2282_),
    .D(_2283_),
    .X(_2284_));
 sky130_fd_sc_hd__o22ai_1 _5813_ (.A1(_1196_),
    .A2(_3263_),
    .B1(_1320_),
    .B2(_3267_),
    .Y(_2285_));
 sky130_fd_sc_hd__a22o_1 _5814_ (.A1(_3270_),
    .A2(_3341_),
    .B1(_3273_),
    .B2(_3347_),
    .X(_2286_));
 sky130_fd_sc_hd__nor2_1 _5815_ (.A(_2285_),
    .B(_2286_),
    .Y(_2287_));
 sky130_fd_sc_hd__o22ai_1 _5816_ (.A1(_0952_),
    .A2(_3288_),
    .B1(_1081_),
    .B2(_3292_),
    .Y(_2288_));
 sky130_fd_sc_hd__a221oi_1 _5817_ (.A1(_3353_),
    .A2(_3280_),
    .B1(_3357_),
    .B2(_3284_),
    .C1(_2288_),
    .Y(_2289_));
 sky130_fd_sc_hd__and4_1 _5818_ (.A(_2279_),
    .B(_2284_),
    .C(_2287_),
    .D(_2289_),
    .X(_2290_));
 sky130_fd_sc_hd__nand2_1 _5819_ (.A(_3308_),
    .B(_3028_),
    .Y(_2291_));
 sky130_fd_sc_hd__nand2_1 _5820_ (.A(_3312_),
    .B(_3025_),
    .Y(_2292_));
 sky130_fd_sc_hd__nand2_1 _5821_ (.A(_2291_),
    .B(_2292_),
    .Y(_2293_));
 sky130_fd_sc_hd__a221oi_1 _5822_ (.A1(_3031_),
    .A2(_3302_),
    .B1(_3034_),
    .B2(_3306_),
    .C1(_2293_),
    .Y(_2294_));
 sky130_fd_sc_hd__nand2_1 _5823_ (.A(_3325_),
    .B(_3010_),
    .Y(_2295_));
 sky130_fd_sc_hd__nand2_1 _5824_ (.A(_3329_),
    .B(_2998_),
    .Y(_2296_));
 sky130_fd_sc_hd__nand2_1 _5825_ (.A(_2295_),
    .B(_2296_),
    .Y(_2297_));
 sky130_fd_sc_hd__a221oi_1 _5826_ (.A1(_0674_),
    .A2(_3320_),
    .B1(_0675_),
    .B2(_3323_),
    .C1(_2297_),
    .Y(_2298_));
 sky130_fd_sc_hd__nand2_1 _5827_ (.A(_3339_),
    .B(_3013_),
    .Y(_2299_));
 sky130_fd_sc_hd__nand2_1 _5828_ (.A(_3343_),
    .B(_3019_),
    .Y(_2300_));
 sky130_fd_sc_hd__or2_1 _5829_ (.A(_0922_),
    .B(_3349_),
    .X(_2301_));
 sky130_fd_sc_hd__o2111a_1 _5830_ (.A1(_3177_),
    .A2(_3337_),
    .B1(_2299_),
    .C1(_2300_),
    .D1(_2301_),
    .X(_2302_));
 sky130_fd_sc_hd__nand2_1 _5831_ (.A(_3364_),
    .B(_3044_),
    .Y(_2303_));
 sky130_fd_sc_hd__o21ai_1 _5832_ (.A1(_3219_),
    .A2(_3362_),
    .B1(_2303_),
    .Y(_2304_));
 sky130_fd_sc_hd__a221oi_1 _5833_ (.A1(_3037_),
    .A2(_3355_),
    .B1(_3040_),
    .B2(_3359_),
    .C1(_2304_),
    .Y(_2305_));
 sky130_fd_sc_hd__and4_1 _5834_ (.A(_2294_),
    .B(_2298_),
    .C(_2302_),
    .D(_2305_),
    .X(_2306_));
 sky130_fd_sc_hd__and4_1 _5835_ (.A(_2266_),
    .B(_2277_),
    .C(_2290_),
    .D(_2306_),
    .X(_2307_));
 sky130_fd_sc_hd__nand2_1 _5836_ (.A(_0333_),
    .B(_0701_),
    .Y(_2308_));
 sky130_fd_sc_hd__nand2_1 _5837_ (.A(_0337_),
    .B(_0400_),
    .Y(_2309_));
 sky130_fd_sc_hd__nand2_1 _5838_ (.A(_2308_),
    .B(_2309_),
    .Y(_2310_));
 sky130_fd_sc_hd__a221oi_1 _5839_ (.A1(_0417_),
    .A2(_0327_),
    .B1(_0423_),
    .B2(_0331_),
    .C1(_2310_),
    .Y(_2311_));
 sky130_fd_sc_hd__o22ai_1 _5840_ (.A1(_0853_),
    .A2(_0344_),
    .B1(_0986_),
    .B2(_0348_),
    .Y(_2312_));
 sky130_fd_sc_hd__a22o_1 _5841_ (.A1(_0351_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[52] ),
    .B1(_0354_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[53] ),
    .X(_2313_));
 sky130_fd_sc_hd__nor2_1 _5842_ (.A(_2312_),
    .B(_2313_),
    .Y(_2314_));
 sky130_fd_sc_hd__nand2_1 _5843_ (.A(_0370_),
    .B(_0443_),
    .Y(_2315_));
 sky130_fd_sc_hd__o21ai_1 _5844_ (.A1(_0438_),
    .A2(_0368_),
    .B1(_2315_),
    .Y(_2316_));
 sky130_fd_sc_hd__a221oi_1 _5845_ (.A1(_0389_),
    .A2(_0361_),
    .B1(_0695_),
    .B2(_0365_),
    .C1(_2316_),
    .Y(_2317_));
 sky130_fd_sc_hd__nand2_1 _5846_ (.A(_0387_),
    .B(_0447_),
    .Y(_2318_));
 sky130_fd_sc_hd__o21ai_1 _5847_ (.A1(_0848_),
    .A2(_0385_),
    .B1(_2318_),
    .Y(_2319_));
 sky130_fd_sc_hd__a221oi_1 _5848_ (.A1(_0421_),
    .A2(_0378_),
    .B1(_0411_),
    .B2(_0382_),
    .C1(_2319_),
    .Y(_2320_));
 sky130_fd_sc_hd__and4_1 _5849_ (.A(_2311_),
    .B(_2314_),
    .C(_2317_),
    .D(_2320_),
    .X(_2321_));
 sky130_fd_sc_hd__nand2_1 _5850_ (.A(_0398_),
    .B(_3129_),
    .Y(_2322_));
 sky130_fd_sc_hd__nand2_1 _5851_ (.A(_0402_),
    .B(_3095_),
    .Y(_2323_));
 sky130_fd_sc_hd__or2_1 _5852_ (.A(_3137_),
    .B(_0407_),
    .X(_2324_));
 sky130_fd_sc_hd__o2111a_1 _5853_ (.A1(_0903_),
    .A2(_0396_),
    .B1(_2322_),
    .C1(_2323_),
    .D1(_2324_),
    .X(_2325_));
 sky130_fd_sc_hd__nand2_1 _5854_ (.A(_0415_),
    .B(_3134_),
    .Y(_2326_));
 sky130_fd_sc_hd__nand2_1 _5855_ (.A(_0419_),
    .B(_3076_),
    .Y(_2327_));
 sky130_fd_sc_hd__or2_1 _5856_ (.A(_3120_),
    .B(_0425_),
    .X(_2328_));
 sky130_fd_sc_hd__o2111a_1 _5857_ (.A1(_3086_),
    .A2(_0413_),
    .B1(_2326_),
    .C1(_2327_),
    .D1(_2328_),
    .X(_2329_));
 sky130_fd_sc_hd__nand2_1 _5858_ (.A(_0441_),
    .B(_0455_),
    .Y(_2330_));
 sky130_fd_sc_hd__o21ai_1 _5859_ (.A1(_0981_),
    .A2(_0439_),
    .B1(_2330_),
    .Y(_2331_));
 sky130_fd_sc_hd__a221oi_1 _5860_ (.A1(_3107_),
    .A2(_0431_),
    .B1(_3115_),
    .B2(_0435_),
    .C1(_2331_),
    .Y(_2332_));
 sky130_fd_sc_hd__nand2_1 _5861_ (.A(_0459_),
    .B(_3161_),
    .Y(_2333_));
 sky130_fd_sc_hd__o21ai_1 _5862_ (.A1(_1031_),
    .A2(_0457_),
    .B1(_2333_),
    .Y(_2334_));
 sky130_fd_sc_hd__a221oi_1 _5863_ (.A1(_3057_),
    .A2(_0449_),
    .B1(_3069_),
    .B2(_0453_),
    .C1(_2334_),
    .Y(_2335_));
 sky130_fd_sc_hd__and4_1 _5864_ (.A(_2325_),
    .B(_2329_),
    .C(_2332_),
    .D(_2335_),
    .X(_2336_));
 sky130_fd_sc_hd__and2_1 _5865_ (.A(_2321_),
    .B(_2336_),
    .X(_2337_));
 sky130_fd_sc_hd__nand2_1 _5866_ (.A(_0473_),
    .B(_0356_),
    .Y(_2338_));
 sky130_fd_sc_hd__a22o_1 _5867_ (.A1(_0477_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[40] ),
    .B1(_0480_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[41] ),
    .X(_2339_));
 sky130_fd_sc_hd__inv_2 _5868_ (.A(_2339_),
    .Y(_2340_));
 sky130_fd_sc_hd__o211a_1 _5869_ (.A1(_0685_),
    .A2(_0471_),
    .B1(_2338_),
    .C1(_2340_),
    .X(_2341_));
 sky130_fd_sc_hd__nand2_1 _5870_ (.A(_0497_),
    .B(_0363_),
    .Y(_2342_));
 sky130_fd_sc_hd__o21ai_1 _5871_ (.A1(_1619_),
    .A2(_0495_),
    .B1(_2342_),
    .Y(_2343_));
 sky130_fd_sc_hd__a221oi_1 _5872_ (.A1(_0521_),
    .A2(_0487_),
    .B1(_0525_),
    .B2(_0491_),
    .C1(_2343_),
    .Y(_2344_));
 sky130_fd_sc_hd__nand2_1 _5873_ (.A(_0507_),
    .B(_0691_),
    .Y(_2345_));
 sky130_fd_sc_hd__nand2_1 _5874_ (.A(_0511_),
    .B(_0689_),
    .Y(_2346_));
 sky130_fd_sc_hd__or2_1 _5875_ (.A(_0690_),
    .B(_0517_),
    .X(_2347_));
 sky130_fd_sc_hd__o2111a_1 _5876_ (.A1(_0347_),
    .A2(_0505_),
    .B1(_2345_),
    .C1(_2346_),
    .D1(_2347_),
    .X(_2348_));
 sky130_fd_sc_hd__nand2_1 _5877_ (.A(_0529_),
    .B(_0329_),
    .Y(_2349_));
 sky130_fd_sc_hd__nand2_1 _5878_ (.A(_0533_),
    .B(_0323_),
    .Y(_2350_));
 sky130_fd_sc_hd__nand2_1 _5879_ (.A(_2349_),
    .B(_2350_),
    .Y(_2351_));
 sky130_fd_sc_hd__a221oi_1 _5880_ (.A1(_0376_),
    .A2(_0523_),
    .B1(_0380_),
    .B2(_0527_),
    .C1(_2351_),
    .Y(_2352_));
 sky130_fd_sc_hd__and4_1 _5881_ (.A(_2341_),
    .B(_2344_),
    .C(_2348_),
    .D(_2352_),
    .X(_2353_));
 sky130_fd_sc_hd__nand2_1 _5882_ (.A(_0546_),
    .B(_0513_),
    .Y(_2354_));
 sky130_fd_sc_hd__nand2_1 _5883_ (.A(_0550_),
    .B(_0493_),
    .Y(_2355_));
 sky130_fd_sc_hd__or2_1 _5884_ (.A(_0516_),
    .B(_0555_),
    .X(_2356_));
 sky130_fd_sc_hd__o2111a_1 _5885_ (.A1(_0728_),
    .A2(_0544_),
    .B1(_2354_),
    .C1(_2355_),
    .D1(_2356_),
    .X(_2357_));
 sky130_fd_sc_hd__nand2_1 _5886_ (.A(_0562_),
    .B(_0467_),
    .Y(_2358_));
 sky130_fd_sc_hd__nand2_1 _5887_ (.A(_0565_),
    .B(_0509_),
    .Y(_2359_));
 sky130_fd_sc_hd__or2_1 _5888_ (.A(_0504_),
    .B(_0569_),
    .X(_2360_));
 sky130_fd_sc_hd__o2111a_1 _5889_ (.A1(_0723_),
    .A2(_0560_),
    .B1(_2358_),
    .C1(_2359_),
    .D1(_2360_),
    .X(_2361_));
 sky130_fd_sc_hd__or2_1 _5890_ (.A(_1150_),
    .B(_0583_),
    .X(_2362_));
 sky130_fd_sc_hd__o221a_1 _5891_ (.A1(_1022_),
    .A2(_0575_),
    .B1(_0890_),
    .B2(_0579_),
    .C1(_2362_),
    .X(_2363_));
 sky130_fd_sc_hd__o22ai_1 _5892_ (.A1(_0862_),
    .A2(_0594_),
    .B1(_0995_),
    .B2(_0597_),
    .Y(_2364_));
 sky130_fd_sc_hd__a221oi_1 _5893_ (.A1(_0535_),
    .A2(_0588_),
    .B1(_0531_),
    .B2(_0591_),
    .C1(_2364_),
    .Y(_2365_));
 sky130_fd_sc_hd__and4_1 _5894_ (.A(_2357_),
    .B(_2361_),
    .C(_2363_),
    .D(_2365_),
    .X(_2366_));
 sky130_fd_sc_hd__and3_1 _5895_ (.A(_2337_),
    .B(_2353_),
    .C(_2366_),
    .X(_2367_));
 sky130_fd_sc_hd__nand2_1 _5896_ (.A(_0605_),
    .B(\egd_top.BitStream_buffer.BS_buffer[14] ),
    .Y(_2368_));
 sky130_fd_sc_hd__nand3_2 _5897_ (.A(_2307_),
    .B(_2367_),
    .C(_2368_),
    .Y(_2369_));
 sky130_fd_sc_hd__inv_2 _5898_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[1] ),
    .Y(_2370_));
 sky130_fd_sc_hd__a21oi_1 _5899_ (.A1(_2370_),
    .A2(_2996_),
    .B1(_2937_),
    .Y(_2371_));
 sky130_fd_sc_hd__o21a_1 _5900_ (.A1(_0898_),
    .A2(_2369_),
    .B1(_2371_),
    .X(_0283_));
 sky130_fd_sc_hd__clkbuf_4 _5901_ (.A(net19),
    .X(_2372_));
 sky130_fd_sc_hd__nand2_1 _5902_ (.A(_3004_),
    .B(_2978_),
    .Y(_2373_));
 sky130_fd_sc_hd__and3_1 _5903_ (.A(_3007_),
    .B(_2372_),
    .C(_2373_),
    .X(_2374_));
 sky130_fd_sc_hd__clkbuf_1 _5904_ (.A(_2374_),
    .X(_0282_));
 sky130_fd_sc_hd__nand2_1 _5905_ (.A(_3003_),
    .B(_2971_),
    .Y(_2375_));
 sky130_fd_sc_hd__and3_1 _5906_ (.A(_3004_),
    .B(_2372_),
    .C(_2375_),
    .X(_2376_));
 sky130_fd_sc_hd__clkbuf_1 _5907_ (.A(_2376_),
    .X(_0281_));
 sky130_fd_sc_hd__or2_1 _5908_ (.A(\egd_top.BitStream_buffer.buffer_index[4] ),
    .B(_3002_),
    .X(_2377_));
 sky130_fd_sc_hd__and3_1 _5909_ (.A(_2377_),
    .B(_2372_),
    .C(_3003_),
    .X(_2378_));
 sky130_fd_sc_hd__clkbuf_1 _5910_ (.A(_2378_),
    .X(_0280_));
 sky130_fd_sc_hd__nand2_2 _5911_ (.A(_3002_),
    .B(_2979_),
    .Y(_2379_));
 sky130_fd_sc_hd__buf_4 _5912_ (.A(_2379_),
    .X(_2380_));
 sky130_fd_sc_hd__mux2_1 _5913_ (.A0(net7),
    .A1(_0607_),
    .S(_2380_),
    .X(_2381_));
 sky130_fd_sc_hd__and2_1 _5914_ (.A(_2381_),
    .B(_3042_),
    .X(_2382_));
 sky130_fd_sc_hd__clkbuf_1 _5915_ (.A(_2382_),
    .X(_0279_));
 sky130_fd_sc_hd__mux2_1 _5916_ (.A0(net6),
    .A1(_0577_),
    .S(_2380_),
    .X(_2383_));
 sky130_fd_sc_hd__and2_1 _5917_ (.A(_2383_),
    .B(_3042_),
    .X(_2384_));
 sky130_fd_sc_hd__clkbuf_1 _5918_ (.A(_2384_),
    .X(_0278_));
 sky130_fd_sc_hd__mux2_1 _5919_ (.A0(net5),
    .A1(_0573_),
    .S(_2380_),
    .X(_2385_));
 sky130_fd_sc_hd__and2_1 _5920_ (.A(_2385_),
    .B(_3042_),
    .X(_2386_));
 sky130_fd_sc_hd__clkbuf_1 _5921_ (.A(_2386_),
    .X(_0277_));
 sky130_fd_sc_hd__mux2_1 _5922_ (.A0(net4),
    .A1(_0581_),
    .S(_2380_),
    .X(_2387_));
 sky130_fd_sc_hd__and2_1 _5923_ (.A(_2387_),
    .B(_3042_),
    .X(_2388_));
 sky130_fd_sc_hd__clkbuf_1 _5924_ (.A(_2388_),
    .X(_0276_));
 sky130_fd_sc_hd__mux2_1 _5925_ (.A0(net3),
    .A1(_0552_),
    .S(_2380_),
    .X(_2389_));
 sky130_fd_sc_hd__and2_1 _5926_ (.A(_2389_),
    .B(_3042_),
    .X(_2390_));
 sky130_fd_sc_hd__clkbuf_1 _5927_ (.A(_2390_),
    .X(_0275_));
 sky130_fd_sc_hd__mux2_1 _5928_ (.A0(net2),
    .A1(_0540_),
    .S(_2380_),
    .X(_2391_));
 sky130_fd_sc_hd__and2_1 _5929_ (.A(_2391_),
    .B(_3042_),
    .X(_2392_));
 sky130_fd_sc_hd__clkbuf_1 _5930_ (.A(_2392_),
    .X(_0274_));
 sky130_fd_sc_hd__mux2_1 _5931_ (.A0(net16),
    .A1(_0548_),
    .S(_2380_),
    .X(_2393_));
 sky130_fd_sc_hd__and2_1 _5932_ (.A(_2393_),
    .B(_3042_),
    .X(_2394_));
 sky130_fd_sc_hd__clkbuf_1 _5933_ (.A(_2394_),
    .X(_0273_));
 sky130_fd_sc_hd__mux2_1 _5934_ (.A0(net15),
    .A1(\egd_top.BitStream_buffer.BS_buffer[7] ),
    .S(_2380_),
    .X(_2395_));
 sky130_fd_sc_hd__buf_2 _5935_ (.A(_2932_),
    .X(_2396_));
 sky130_fd_sc_hd__and2_1 _5936_ (.A(_2395_),
    .B(_2396_),
    .X(_2397_));
 sky130_fd_sc_hd__clkbuf_1 _5937_ (.A(_2397_),
    .X(_0272_));
 sky130_fd_sc_hd__mux2_1 _5938_ (.A0(net14),
    .A1(\egd_top.BitStream_buffer.BS_buffer[8] ),
    .S(_2380_),
    .X(_2398_));
 sky130_fd_sc_hd__and2_1 _5939_ (.A(_2398_),
    .B(_2396_),
    .X(_2399_));
 sky130_fd_sc_hd__clkbuf_1 _5940_ (.A(_2399_),
    .X(_0271_));
 sky130_fd_sc_hd__mux2_1 _5941_ (.A0(net13),
    .A1(\egd_top.BitStream_buffer.BS_buffer[9] ),
    .S(_2380_),
    .X(_2400_));
 sky130_fd_sc_hd__and2_1 _5942_ (.A(_2400_),
    .B(_2396_),
    .X(_2401_));
 sky130_fd_sc_hd__clkbuf_1 _5943_ (.A(_2401_),
    .X(_0270_));
 sky130_fd_sc_hd__mux2_1 _5944_ (.A0(net12),
    .A1(\egd_top.BitStream_buffer.BS_buffer[10] ),
    .S(_2380_),
    .X(_2402_));
 sky130_fd_sc_hd__and2_1 _5945_ (.A(_2402_),
    .B(_2396_),
    .X(_2403_));
 sky130_fd_sc_hd__clkbuf_1 _5946_ (.A(_2403_),
    .X(_0269_));
 sky130_fd_sc_hd__mux2_1 _5947_ (.A0(net11),
    .A1(\egd_top.BitStream_buffer.BS_buffer[11] ),
    .S(_2380_),
    .X(_2404_));
 sky130_fd_sc_hd__and2_1 _5948_ (.A(_2404_),
    .B(_2396_),
    .X(_2405_));
 sky130_fd_sc_hd__clkbuf_1 _5949_ (.A(_2405_),
    .X(_0268_));
 sky130_fd_sc_hd__mux2_1 _5950_ (.A0(net10),
    .A1(\egd_top.BitStream_buffer.BS_buffer[12] ),
    .S(_2379_),
    .X(_2406_));
 sky130_fd_sc_hd__and2_1 _5951_ (.A(_2406_),
    .B(_2396_),
    .X(_2407_));
 sky130_fd_sc_hd__clkbuf_1 _5952_ (.A(_2407_),
    .X(_0267_));
 sky130_fd_sc_hd__mux2_1 _5953_ (.A0(net9),
    .A1(\egd_top.BitStream_buffer.BS_buffer[13] ),
    .S(_2379_),
    .X(_2408_));
 sky130_fd_sc_hd__and2_1 _5954_ (.A(_2408_),
    .B(_2396_),
    .X(_2409_));
 sky130_fd_sc_hd__clkbuf_1 _5955_ (.A(_2409_),
    .X(_0266_));
 sky130_fd_sc_hd__mux2_1 _5956_ (.A0(net8),
    .A1(\egd_top.BitStream_buffer.BS_buffer[14] ),
    .S(_2379_),
    .X(_2410_));
 sky130_fd_sc_hd__and2_1 _5957_ (.A(_2410_),
    .B(_2396_),
    .X(_2411_));
 sky130_fd_sc_hd__clkbuf_1 _5958_ (.A(_2411_),
    .X(_0265_));
 sky130_fd_sc_hd__mux2_1 _5959_ (.A0(net1),
    .A1(\egd_top.BitStream_buffer.BS_buffer[15] ),
    .S(_2379_),
    .X(_2412_));
 sky130_fd_sc_hd__and2_1 _5960_ (.A(_2412_),
    .B(_2396_),
    .X(_2413_));
 sky130_fd_sc_hd__clkbuf_1 _5961_ (.A(_2413_),
    .X(_0264_));
 sky130_fd_sc_hd__or4b_4 _5962_ (.A(\egd_top.BitStream_buffer.buffer_index[6] ),
    .B(\egd_top.BitStream_buffer.buffer_index[5] ),
    .C(_2972_),
    .D_N(_3002_),
    .X(_2414_));
 sky130_fd_sc_hd__buf_4 _5963_ (.A(_2414_),
    .X(_2415_));
 sky130_fd_sc_hd__mux2_1 _5964_ (.A0(net7),
    .A1(\egd_top.BitStream_buffer.BS_buffer[16] ),
    .S(_2415_),
    .X(_2416_));
 sky130_fd_sc_hd__and2_1 _5965_ (.A(_2416_),
    .B(_2396_),
    .X(_2417_));
 sky130_fd_sc_hd__clkbuf_1 _5966_ (.A(_2417_),
    .X(_0263_));
 sky130_fd_sc_hd__mux2_1 _5967_ (.A0(net6),
    .A1(_0489_),
    .S(_2415_),
    .X(_2418_));
 sky130_fd_sc_hd__and2_1 _5968_ (.A(_2418_),
    .B(_2396_),
    .X(_2419_));
 sky130_fd_sc_hd__clkbuf_1 _5969_ (.A(_2419_),
    .X(_0262_));
 sky130_fd_sc_hd__mux2_1 _5970_ (.A0(net5),
    .A1(_0493_),
    .S(_2415_),
    .X(_2420_));
 sky130_fd_sc_hd__and2_1 _5971_ (.A(_2420_),
    .B(_2396_),
    .X(_2421_));
 sky130_fd_sc_hd__clkbuf_1 _5972_ (.A(_2421_),
    .X(_0261_));
 sky130_fd_sc_hd__mux2_1 _5973_ (.A0(net4),
    .A1(_0499_),
    .S(_2415_),
    .X(_2422_));
 sky130_fd_sc_hd__buf_2 _5974_ (.A(_2932_),
    .X(_2423_));
 sky130_fd_sc_hd__and2_1 _5975_ (.A(_2422_),
    .B(_2423_),
    .X(_2424_));
 sky130_fd_sc_hd__clkbuf_1 _5976_ (.A(_2424_),
    .X(_0260_));
 sky130_fd_sc_hd__mux2_1 _5977_ (.A0(net3),
    .A1(_0513_),
    .S(_2415_),
    .X(_2425_));
 sky130_fd_sc_hd__and2_1 _5978_ (.A(_2425_),
    .B(_2423_),
    .X(_2426_));
 sky130_fd_sc_hd__clkbuf_1 _5979_ (.A(_2426_),
    .X(_0259_));
 sky130_fd_sc_hd__mux2_1 _5980_ (.A0(net2),
    .A1(_0515_),
    .S(_2415_),
    .X(_2427_));
 sky130_fd_sc_hd__and2_1 _5981_ (.A(_2427_),
    .B(_2423_),
    .X(_2428_));
 sky130_fd_sc_hd__clkbuf_1 _5982_ (.A(_2428_),
    .X(_0258_));
 sky130_fd_sc_hd__mux2_1 _5983_ (.A0(net16),
    .A1(_0509_),
    .S(_2415_),
    .X(_2429_));
 sky130_fd_sc_hd__and2_1 _5984_ (.A(_2429_),
    .B(_2423_),
    .X(_2430_));
 sky130_fd_sc_hd__clkbuf_1 _5985_ (.A(_2430_),
    .X(_0257_));
 sky130_fd_sc_hd__mux2_1 _5986_ (.A0(net15),
    .A1(_0503_),
    .S(_2415_),
    .X(_2431_));
 sky130_fd_sc_hd__and2_1 _5987_ (.A(_2431_),
    .B(_2423_),
    .X(_2432_));
 sky130_fd_sc_hd__clkbuf_1 _5988_ (.A(_2432_),
    .X(_0256_));
 sky130_fd_sc_hd__mux2_1 _5989_ (.A0(net14),
    .A1(_0467_),
    .S(_2415_),
    .X(_2433_));
 sky130_fd_sc_hd__and2_1 _5990_ (.A(_2433_),
    .B(_2423_),
    .X(_2434_));
 sky130_fd_sc_hd__clkbuf_1 _5991_ (.A(_2434_),
    .X(_0255_));
 sky130_fd_sc_hd__mux2_1 _5992_ (.A0(net13),
    .A1(_0475_),
    .S(_2415_),
    .X(_2435_));
 sky130_fd_sc_hd__and2_1 _5993_ (.A(_2435_),
    .B(_2423_),
    .X(_2436_));
 sky130_fd_sc_hd__clkbuf_1 _5994_ (.A(_2436_),
    .X(_0254_));
 sky130_fd_sc_hd__mux2_1 _5995_ (.A0(net12),
    .A1(_0479_),
    .S(_2415_),
    .X(_2437_));
 sky130_fd_sc_hd__and2_1 _5996_ (.A(_2437_),
    .B(_2423_),
    .X(_2438_));
 sky130_fd_sc_hd__clkbuf_1 _5997_ (.A(_2438_),
    .X(_0253_));
 sky130_fd_sc_hd__mux2_1 _5998_ (.A0(net11),
    .A1(_0482_),
    .S(_2415_),
    .X(_2439_));
 sky130_fd_sc_hd__and2_1 _5999_ (.A(_2439_),
    .B(_2423_),
    .X(_2440_));
 sky130_fd_sc_hd__clkbuf_1 _6000_ (.A(_2440_),
    .X(_0252_));
 sky130_fd_sc_hd__mux2_1 _6001_ (.A0(net10),
    .A1(_0535_),
    .S(_2414_),
    .X(_2441_));
 sky130_fd_sc_hd__and2_1 _6002_ (.A(_2441_),
    .B(_2423_),
    .X(_2442_));
 sky130_fd_sc_hd__clkbuf_1 _6003_ (.A(_2442_),
    .X(_0251_));
 sky130_fd_sc_hd__mux2_1 _6004_ (.A0(net9),
    .A1(_0531_),
    .S(_2414_),
    .X(_2443_));
 sky130_fd_sc_hd__and2_1 _6005_ (.A(_2443_),
    .B(_2423_),
    .X(_2444_));
 sky130_fd_sc_hd__clkbuf_1 _6006_ (.A(_2444_),
    .X(_0250_));
 sky130_fd_sc_hd__mux2_1 _6007_ (.A0(net8),
    .A1(_0521_),
    .S(_2414_),
    .X(_2445_));
 sky130_fd_sc_hd__and2_1 _6008_ (.A(_2445_),
    .B(_2423_),
    .X(_2446_));
 sky130_fd_sc_hd__clkbuf_1 _6009_ (.A(_2446_),
    .X(_0249_));
 sky130_fd_sc_hd__mux2_1 _6010_ (.A0(net1),
    .A1(_0525_),
    .S(_2414_),
    .X(_2447_));
 sky130_fd_sc_hd__buf_2 _6011_ (.A(_2932_),
    .X(_2448_));
 sky130_fd_sc_hd__and2_1 _6012_ (.A(_2447_),
    .B(_2448_),
    .X(_2449_));
 sky130_fd_sc_hd__clkbuf_1 _6013_ (.A(_2449_),
    .X(_0248_));
 sky130_fd_sc_hd__or4b_4 _6014_ (.A(net200),
    .B(_2971_),
    .C(net196),
    .D_N(_3002_),
    .X(_2450_));
 sky130_fd_sc_hd__buf_4 _6015_ (.A(_2450_),
    .X(_2451_));
 sky130_fd_sc_hd__mux2_1 _6016_ (.A0(net7),
    .A1(_0359_),
    .S(_2451_),
    .X(_2452_));
 sky130_fd_sc_hd__and2_1 _6017_ (.A(_2452_),
    .B(_2448_),
    .X(_2453_));
 sky130_fd_sc_hd__clkbuf_1 _6018_ (.A(_2453_),
    .X(_0247_));
 sky130_fd_sc_hd__mux2_1 _6019_ (.A0(net6),
    .A1(_0363_),
    .S(_2451_),
    .X(_2454_));
 sky130_fd_sc_hd__and2_1 _6020_ (.A(_2454_),
    .B(_2448_),
    .X(_2455_));
 sky130_fd_sc_hd__clkbuf_1 _6021_ (.A(_2455_),
    .X(_0246_));
 sky130_fd_sc_hd__mux2_1 _6022_ (.A0(net5),
    .A1(_0689_),
    .S(_2451_),
    .X(_2456_));
 sky130_fd_sc_hd__and2_1 _6023_ (.A(_2456_),
    .B(_2448_),
    .X(_2457_));
 sky130_fd_sc_hd__clkbuf_1 _6024_ (.A(_2457_),
    .X(_0245_));
 sky130_fd_sc_hd__mux2_1 _6025_ (.A0(net4),
    .A1(_0372_),
    .S(_2451_),
    .X(_2458_));
 sky130_fd_sc_hd__and2_1 _6026_ (.A(_2458_),
    .B(_2448_),
    .X(_2459_));
 sky130_fd_sc_hd__clkbuf_1 _6027_ (.A(_2459_),
    .X(_0244_));
 sky130_fd_sc_hd__mux2_1 _6028_ (.A0(net3),
    .A1(_0691_),
    .S(_2451_),
    .X(_2460_));
 sky130_fd_sc_hd__and2_1 _6029_ (.A(_2460_),
    .B(_2448_),
    .X(_2461_));
 sky130_fd_sc_hd__clkbuf_1 _6030_ (.A(_2461_),
    .X(_0243_));
 sky130_fd_sc_hd__mux2_1 _6031_ (.A0(net2),
    .A1(_0346_),
    .S(_2451_),
    .X(_2462_));
 sky130_fd_sc_hd__and2_1 _6032_ (.A(_2462_),
    .B(_2448_),
    .X(_2463_));
 sky130_fd_sc_hd__clkbuf_1 _6033_ (.A(_2463_),
    .X(_0242_));
 sky130_fd_sc_hd__mux2_1 _6034_ (.A0(net16),
    .A1(_0353_),
    .S(_2451_),
    .X(_2464_));
 sky130_fd_sc_hd__and2_1 _6035_ (.A(_2464_),
    .B(_2448_),
    .X(_2465_));
 sky130_fd_sc_hd__clkbuf_1 _6036_ (.A(_2465_),
    .X(_0241_));
 sky130_fd_sc_hd__mux2_1 _6037_ (.A0(net15),
    .A1(_0356_),
    .S(_2451_),
    .X(_2466_));
 sky130_fd_sc_hd__and2_1 _6038_ (.A(_2466_),
    .B(_2448_),
    .X(_2467_));
 sky130_fd_sc_hd__clkbuf_1 _6039_ (.A(_2467_),
    .X(_0240_));
 sky130_fd_sc_hd__mux2_1 _6040_ (.A0(net14),
    .A1(_0339_),
    .S(_2451_),
    .X(_2468_));
 sky130_fd_sc_hd__and2_1 _6041_ (.A(_2468_),
    .B(_2448_),
    .X(_2469_));
 sky130_fd_sc_hd__clkbuf_1 _6042_ (.A(_2469_),
    .X(_0239_));
 sky130_fd_sc_hd__mux2_1 _6043_ (.A0(net13),
    .A1(_0335_),
    .S(_2451_),
    .X(_2470_));
 sky130_fd_sc_hd__and2_1 _6044_ (.A(_2470_),
    .B(_2448_),
    .X(_2471_));
 sky130_fd_sc_hd__clkbuf_1 _6045_ (.A(_2471_),
    .X(_0238_));
 sky130_fd_sc_hd__mux2_1 _6046_ (.A0(net12),
    .A1(_0323_),
    .S(_2451_),
    .X(_2472_));
 sky130_fd_sc_hd__and2_1 _6047_ (.A(_2472_),
    .B(_2448_),
    .X(_2473_));
 sky130_fd_sc_hd__clkbuf_1 _6048_ (.A(_2473_),
    .X(_0237_));
 sky130_fd_sc_hd__mux2_1 _6049_ (.A0(net11),
    .A1(_0329_),
    .S(_2451_),
    .X(_2474_));
 sky130_fd_sc_hd__buf_2 _6050_ (.A(_2932_),
    .X(_2475_));
 sky130_fd_sc_hd__and2_1 _6051_ (.A(_2474_),
    .B(_2475_),
    .X(_2476_));
 sky130_fd_sc_hd__clkbuf_1 _6052_ (.A(_2476_),
    .X(_0236_));
 sky130_fd_sc_hd__mux2_1 _6053_ (.A0(net10),
    .A1(_0376_),
    .S(_2450_),
    .X(_2477_));
 sky130_fd_sc_hd__and2_1 _6054_ (.A(_2477_),
    .B(_2475_),
    .X(_2478_));
 sky130_fd_sc_hd__clkbuf_1 _6055_ (.A(_2478_),
    .X(_0235_));
 sky130_fd_sc_hd__mux2_1 _6056_ (.A0(net9),
    .A1(_0380_),
    .S(_2450_),
    .X(_2479_));
 sky130_fd_sc_hd__and2_1 _6057_ (.A(_2479_),
    .B(_2475_),
    .X(_2480_));
 sky130_fd_sc_hd__clkbuf_1 _6058_ (.A(_2480_),
    .X(_0234_));
 sky130_fd_sc_hd__mux2_1 _6059_ (.A0(net8),
    .A1(_0389_),
    .S(net203),
    .X(_2481_));
 sky130_fd_sc_hd__and2_1 _6060_ (.A(_2481_),
    .B(_2475_),
    .X(_2482_));
 sky130_fd_sc_hd__clkbuf_1 _6061_ (.A(_2482_),
    .X(_0233_));
 sky130_fd_sc_hd__mux2_1 _6062_ (.A0(net1),
    .A1(_0695_),
    .S(_2450_),
    .X(_2483_));
 sky130_fd_sc_hd__and2_1 _6063_ (.A(_2483_),
    .B(_2475_),
    .X(_2484_));
 sky130_fd_sc_hd__clkbuf_1 _6064_ (.A(_2484_),
    .X(_0232_));
 sky130_fd_sc_hd__or2_4 _6065_ (.A(net200),
    .B(_3004_),
    .X(_2485_));
 sky130_fd_sc_hd__buf_4 _6066_ (.A(_2485_),
    .X(_2486_));
 sky130_fd_sc_hd__mux2_1 _6067_ (.A0(net7),
    .A1(_0437_),
    .S(_2486_),
    .X(_2487_));
 sky130_fd_sc_hd__and2_1 _6068_ (.A(_2487_),
    .B(_2475_),
    .X(_2488_));
 sky130_fd_sc_hd__clkbuf_1 _6069_ (.A(_2488_),
    .X(_0231_));
 sky130_fd_sc_hd__mux2_1 _6070_ (.A0(net6),
    .A1(_0443_),
    .S(_2486_),
    .X(_2489_));
 sky130_fd_sc_hd__and2_1 _6071_ (.A(_2489_),
    .B(_2475_),
    .X(_2490_));
 sky130_fd_sc_hd__clkbuf_1 _6072_ (.A(_2490_),
    .X(_0230_));
 sky130_fd_sc_hd__mux2_1 _6073_ (.A0(net5),
    .A1(_0429_),
    .S(_2486_),
    .X(_2491_));
 sky130_fd_sc_hd__and2_1 _6074_ (.A(_2491_),
    .B(_2475_),
    .X(_2492_));
 sky130_fd_sc_hd__clkbuf_1 _6075_ (.A(_2492_),
    .X(_0229_));
 sky130_fd_sc_hd__mux2_1 _6076_ (.A0(net4),
    .A1(_0433_),
    .S(_2486_),
    .X(_2493_));
 sky130_fd_sc_hd__and2_1 _6077_ (.A(_2493_),
    .B(_2475_),
    .X(_2494_));
 sky130_fd_sc_hd__clkbuf_1 _6078_ (.A(_2494_),
    .X(_0228_));
 sky130_fd_sc_hd__mux2_1 _6079_ (.A0(net3),
    .A1(_0404_),
    .S(_2486_),
    .X(_2495_));
 sky130_fd_sc_hd__and2_1 _6080_ (.A(_2495_),
    .B(_2475_),
    .X(_2496_));
 sky130_fd_sc_hd__clkbuf_1 _6081_ (.A(_2496_),
    .X(_0227_));
 sky130_fd_sc_hd__mux2_1 _6082_ (.A0(net2),
    .A1(_0703_),
    .S(_2486_),
    .X(_2497_));
 sky130_fd_sc_hd__and2_1 _6083_ (.A(_2497_),
    .B(_2475_),
    .X(_2498_));
 sky130_fd_sc_hd__clkbuf_1 _6084_ (.A(_2498_),
    .X(_0226_));
 sky130_fd_sc_hd__mux2_1 _6085_ (.A0(net16),
    .A1(_0400_),
    .S(_2486_),
    .X(_2499_));
 sky130_fd_sc_hd__and2_1 _6086_ (.A(_2499_),
    .B(_2475_),
    .X(_2500_));
 sky130_fd_sc_hd__clkbuf_1 _6087_ (.A(_2500_),
    .X(_0225_));
 sky130_fd_sc_hd__mux2_1 _6088_ (.A0(net15),
    .A1(_0701_),
    .S(_2486_),
    .X(_2501_));
 sky130_fd_sc_hd__buf_2 _6089_ (.A(_2932_),
    .X(_2502_));
 sky130_fd_sc_hd__and2_1 _6090_ (.A(_2501_),
    .B(_2502_),
    .X(_2503_));
 sky130_fd_sc_hd__clkbuf_1 _6091_ (.A(_2503_),
    .X(_0224_));
 sky130_fd_sc_hd__mux2_1 _6092_ (.A0(net14),
    .A1(_0417_),
    .S(_2486_),
    .X(_2504_));
 sky130_fd_sc_hd__and2_1 _6093_ (.A(_2504_),
    .B(_2502_),
    .X(_2505_));
 sky130_fd_sc_hd__clkbuf_1 _6094_ (.A(_2505_),
    .X(_0223_));
 sky130_fd_sc_hd__mux2_1 _6095_ (.A0(net13),
    .A1(_0423_),
    .S(_2486_),
    .X(_2506_));
 sky130_fd_sc_hd__and2_1 _6096_ (.A(_2506_),
    .B(_2502_),
    .X(_2507_));
 sky130_fd_sc_hd__clkbuf_1 _6097_ (.A(_2507_),
    .X(_0222_));
 sky130_fd_sc_hd__mux2_1 _6098_ (.A0(net12),
    .A1(_0421_),
    .S(_2486_),
    .X(_2508_));
 sky130_fd_sc_hd__and2_1 _6099_ (.A(_2508_),
    .B(_2502_),
    .X(_2509_));
 sky130_fd_sc_hd__clkbuf_1 _6100_ (.A(_2509_),
    .X(_0221_));
 sky130_fd_sc_hd__mux2_1 _6101_ (.A0(net11),
    .A1(_0411_),
    .S(_2486_),
    .X(_2510_));
 sky130_fd_sc_hd__and2_1 _6102_ (.A(_2510_),
    .B(_2502_),
    .X(_2511_));
 sky130_fd_sc_hd__clkbuf_1 _6103_ (.A(_2511_),
    .X(_0220_));
 sky130_fd_sc_hd__mux2_1 _6104_ (.A0(net10),
    .A1(_0447_),
    .S(_2485_),
    .X(_2512_));
 sky130_fd_sc_hd__and2_1 _6105_ (.A(_2512_),
    .B(_2502_),
    .X(_2513_));
 sky130_fd_sc_hd__clkbuf_1 _6106_ (.A(_2513_),
    .X(_0219_));
 sky130_fd_sc_hd__mux2_1 _6107_ (.A0(net9),
    .A1(_0451_),
    .S(_2485_),
    .X(_2514_));
 sky130_fd_sc_hd__and2_1 _6108_ (.A(_2514_),
    .B(_2502_),
    .X(_2515_));
 sky130_fd_sc_hd__clkbuf_1 _6109_ (.A(_2515_),
    .X(_0218_));
 sky130_fd_sc_hd__mux2_1 _6110_ (.A0(net8),
    .A1(_0461_),
    .S(_2485_),
    .X(_2516_));
 sky130_fd_sc_hd__and2_1 _6111_ (.A(_2516_),
    .B(_2502_),
    .X(_2517_));
 sky130_fd_sc_hd__clkbuf_1 _6112_ (.A(_2517_),
    .X(_0217_));
 sky130_fd_sc_hd__mux2_1 _6113_ (.A0(net1),
    .A1(_0455_),
    .S(_2485_),
    .X(_2518_));
 sky130_fd_sc_hd__and2_1 _6114_ (.A(_2518_),
    .B(_2502_),
    .X(_2519_));
 sky130_fd_sc_hd__clkbuf_1 _6115_ (.A(_2519_),
    .X(_0216_));
 sky130_fd_sc_hd__nand2_2 _6116_ (.A(_3002_),
    .B(_2973_),
    .Y(_2520_));
 sky130_fd_sc_hd__buf_4 _6117_ (.A(_2520_),
    .X(_2521_));
 sky130_fd_sc_hd__mux2_1 _6118_ (.A0(net7),
    .A1(_3107_),
    .S(_2521_),
    .X(_2522_));
 sky130_fd_sc_hd__and2_1 _6119_ (.A(_2522_),
    .B(_2502_),
    .X(_2523_));
 sky130_fd_sc_hd__clkbuf_1 _6120_ (.A(_2523_),
    .X(_0215_));
 sky130_fd_sc_hd__mux2_1 _6121_ (.A0(net6),
    .A1(_3115_),
    .S(_2521_),
    .X(_2524_));
 sky130_fd_sc_hd__and2_1 _6122_ (.A(_2524_),
    .B(_2502_),
    .X(_2525_));
 sky130_fd_sc_hd__clkbuf_1 _6123_ (.A(_2525_),
    .X(_0214_));
 sky130_fd_sc_hd__mux2_1 _6124_ (.A0(net5),
    .A1(_3095_),
    .S(_2521_),
    .X(_2526_));
 sky130_fd_sc_hd__and2_1 _6125_ (.A(_2526_),
    .B(_2502_),
    .X(_2527_));
 sky130_fd_sc_hd__clkbuf_1 _6126_ (.A(_2527_),
    .X(_0213_));
 sky130_fd_sc_hd__mux2_1 _6127_ (.A0(net4),
    .A1(_3102_),
    .S(_2521_),
    .X(_2528_));
 sky130_fd_sc_hd__buf_2 _6128_ (.A(_2932_),
    .X(_2529_));
 sky130_fd_sc_hd__and2_1 _6129_ (.A(_2528_),
    .B(_2529_),
    .X(_2530_));
 sky130_fd_sc_hd__clkbuf_1 _6130_ (.A(_2530_),
    .X(_0212_));
 sky130_fd_sc_hd__mux2_1 _6131_ (.A0(net3),
    .A1(_3129_),
    .S(_2521_),
    .X(_2531_));
 sky130_fd_sc_hd__and2_1 _6132_ (.A(_2531_),
    .B(_2529_),
    .X(_2532_));
 sky130_fd_sc_hd__clkbuf_1 _6133_ (.A(_2532_),
    .X(_0211_));
 sky130_fd_sc_hd__mux2_1 _6134_ (.A0(net2),
    .A1(_3136_),
    .S(_2521_),
    .X(_2533_));
 sky130_fd_sc_hd__and2_1 _6135_ (.A(_2533_),
    .B(_2529_),
    .X(_2534_));
 sky130_fd_sc_hd__clkbuf_1 _6136_ (.A(_2534_),
    .X(_0210_));
 sky130_fd_sc_hd__mux2_1 _6137_ (.A0(net16),
    .A1(_3134_),
    .S(_2521_),
    .X(_2535_));
 sky130_fd_sc_hd__and2_1 _6138_ (.A(_2535_),
    .B(_2529_),
    .X(_2536_));
 sky130_fd_sc_hd__clkbuf_1 _6139_ (.A(_2536_),
    .X(_0209_));
 sky130_fd_sc_hd__mux2_1 _6140_ (.A0(net15),
    .A1(_3119_),
    .S(_2521_),
    .X(_2537_));
 sky130_fd_sc_hd__and2_1 _6141_ (.A(_2537_),
    .B(_2529_),
    .X(_2538_));
 sky130_fd_sc_hd__clkbuf_1 _6142_ (.A(_2538_),
    .X(_0208_));
 sky130_fd_sc_hd__mux2_1 _6143_ (.A0(net14),
    .A1(_3076_),
    .S(_2521_),
    .X(_2539_));
 sky130_fd_sc_hd__and2_1 _6144_ (.A(_2539_),
    .B(_2529_),
    .X(_2540_));
 sky130_fd_sc_hd__clkbuf_1 _6145_ (.A(_2540_),
    .X(_0207_));
 sky130_fd_sc_hd__mux2_1 _6146_ (.A0(net13),
    .A1(_3085_),
    .S(_2521_),
    .X(_2541_));
 sky130_fd_sc_hd__and2_1 _6147_ (.A(_2541_),
    .B(_2529_),
    .X(_2542_));
 sky130_fd_sc_hd__clkbuf_1 _6148_ (.A(_2542_),
    .X(_0206_));
 sky130_fd_sc_hd__mux2_1 _6149_ (.A0(net12),
    .A1(_3057_),
    .S(_2521_),
    .X(_2543_));
 sky130_fd_sc_hd__and2_1 _6150_ (.A(_2543_),
    .B(_2529_),
    .X(_2544_));
 sky130_fd_sc_hd__clkbuf_1 _6151_ (.A(_2544_),
    .X(_0205_));
 sky130_fd_sc_hd__mux2_1 _6152_ (.A0(net11),
    .A1(_3069_),
    .S(_2521_),
    .X(_2545_));
 sky130_fd_sc_hd__and2_1 _6153_ (.A(_2545_),
    .B(_2529_),
    .X(_2546_));
 sky130_fd_sc_hd__clkbuf_1 _6154_ (.A(_2546_),
    .X(_0204_));
 sky130_fd_sc_hd__mux2_1 _6155_ (.A0(net10),
    .A1(_3161_),
    .S(_2520_),
    .X(_2547_));
 sky130_fd_sc_hd__and2_1 _6156_ (.A(_2547_),
    .B(_2529_),
    .X(_2548_));
 sky130_fd_sc_hd__clkbuf_1 _6157_ (.A(_2548_),
    .X(_0203_));
 sky130_fd_sc_hd__mux2_1 _6158_ (.A0(net9),
    .A1(_3156_),
    .S(_2520_),
    .X(_2549_));
 sky130_fd_sc_hd__and2_1 _6159_ (.A(_2549_),
    .B(_2529_),
    .X(_2550_));
 sky130_fd_sc_hd__clkbuf_1 _6160_ (.A(_2550_),
    .X(_0202_));
 sky130_fd_sc_hd__mux2_1 _6161_ (.A0(net8),
    .A1(_3144_),
    .S(_2520_),
    .X(_2551_));
 sky130_fd_sc_hd__and2_1 _6162_ (.A(_2551_),
    .B(_2529_),
    .X(_2552_));
 sky130_fd_sc_hd__clkbuf_1 _6163_ (.A(_2552_),
    .X(_0201_));
 sky130_fd_sc_hd__mux2_1 _6164_ (.A0(net1),
    .A1(_3149_),
    .S(_2520_),
    .X(_2553_));
 sky130_fd_sc_hd__clkbuf_4 _6165_ (.A(_2932_),
    .X(_2554_));
 sky130_fd_sc_hd__and2_1 _6166_ (.A(_2553_),
    .B(_2554_),
    .X(_2555_));
 sky130_fd_sc_hd__clkbuf_1 _6167_ (.A(_2555_),
    .X(_0200_));
 sky130_fd_sc_hd__or4b_2 _6168_ (.A(_2978_),
    .B(_2971_),
    .C(net196),
    .D_N(_3002_),
    .X(_2556_));
 sky130_fd_sc_hd__buf_4 _6169_ (.A(_2556_),
    .X(_2557_));
 sky130_fd_sc_hd__mux2_1 _6170_ (.A0(net7),
    .A1(_3318_),
    .S(_2557_),
    .X(_2558_));
 sky130_fd_sc_hd__and2_1 _6171_ (.A(_2558_),
    .B(_2554_),
    .X(_2559_));
 sky130_fd_sc_hd__clkbuf_1 _6172_ (.A(_2559_),
    .X(_0199_));
 sky130_fd_sc_hd__mux2_1 _6173_ (.A0(net6),
    .A1(_3322_),
    .S(_2557_),
    .X(_2560_));
 sky130_fd_sc_hd__and2_1 _6174_ (.A(_2560_),
    .B(_2554_),
    .X(_2561_));
 sky130_fd_sc_hd__clkbuf_1 _6175_ (.A(_2561_),
    .X(_0198_));
 sky130_fd_sc_hd__mux2_1 _6176_ (.A0(net5),
    .A1(_3331_),
    .S(_2557_),
    .X(_2562_));
 sky130_fd_sc_hd__and2_1 _6177_ (.A(_2562_),
    .B(_2554_),
    .X(_2563_));
 sky130_fd_sc_hd__clkbuf_1 _6178_ (.A(_2563_),
    .X(_0197_));
 sky130_fd_sc_hd__mux2_1 _6179_ (.A0(net4),
    .A1(_3327_),
    .S(_2557_),
    .X(_2564_));
 sky130_fd_sc_hd__and2_1 _6180_ (.A(_2564_),
    .B(_2554_),
    .X(_2565_));
 sky130_fd_sc_hd__clkbuf_1 _6181_ (.A(_2565_),
    .X(_0196_));
 sky130_fd_sc_hd__mux2_1 _6182_ (.A0(net3),
    .A1(_3341_),
    .S(_2557_),
    .X(_2566_));
 sky130_fd_sc_hd__and2_1 _6183_ (.A(_2566_),
    .B(_2554_),
    .X(_2567_));
 sky130_fd_sc_hd__clkbuf_1 _6184_ (.A(_2567_),
    .X(_0195_));
 sky130_fd_sc_hd__mux2_1 _6185_ (.A0(net2),
    .A1(_3347_),
    .S(_2557_),
    .X(_2568_));
 sky130_fd_sc_hd__and2_1 _6186_ (.A(_2568_),
    .B(_2554_),
    .X(_2569_));
 sky130_fd_sc_hd__clkbuf_1 _6187_ (.A(_2569_),
    .X(_0194_));
 sky130_fd_sc_hd__mux2_1 _6188_ (.A0(net16),
    .A1(_3345_),
    .S(_2557_),
    .X(_2570_));
 sky130_fd_sc_hd__and2_1 _6189_ (.A(_2570_),
    .B(_2554_),
    .X(_2571_));
 sky130_fd_sc_hd__clkbuf_1 _6190_ (.A(_2571_),
    .X(_0193_));
 sky130_fd_sc_hd__mux2_1 _6191_ (.A0(net15),
    .A1(_3335_),
    .S(_2557_),
    .X(_2572_));
 sky130_fd_sc_hd__and2_1 _6192_ (.A(_2572_),
    .B(_2554_),
    .X(_2573_));
 sky130_fd_sc_hd__clkbuf_1 _6193_ (.A(_2573_),
    .X(_0192_));
 sky130_fd_sc_hd__mux2_1 _6194_ (.A0(net14),
    .A1(_3314_),
    .S(_2557_),
    .X(_2574_));
 sky130_fd_sc_hd__and2_1 _6195_ (.A(_2574_),
    .B(_2554_),
    .X(_2575_));
 sky130_fd_sc_hd__clkbuf_1 _6196_ (.A(_2575_),
    .X(_0191_));
 sky130_fd_sc_hd__mux2_1 _6197_ (.A0(net13),
    .A1(_3310_),
    .S(_2557_),
    .X(_2576_));
 sky130_fd_sc_hd__and2_1 _6198_ (.A(_2576_),
    .B(_2554_),
    .X(_2577_));
 sky130_fd_sc_hd__clkbuf_1 _6199_ (.A(_2577_),
    .X(_0190_));
 sky130_fd_sc_hd__mux2_1 _6200_ (.A0(net12),
    .A1(_3297_),
    .S(_2557_),
    .X(_2578_));
 sky130_fd_sc_hd__and2_1 _6201_ (.A(_2578_),
    .B(_2554_),
    .X(_2579_));
 sky130_fd_sc_hd__clkbuf_1 _6202_ (.A(_2579_),
    .X(_0189_));
 sky130_fd_sc_hd__mux2_1 _6203_ (.A0(net11),
    .A1(_3304_),
    .S(_2557_),
    .X(_2580_));
 sky130_fd_sc_hd__clkbuf_4 _6204_ (.A(_2932_),
    .X(_2581_));
 sky130_fd_sc_hd__and2_1 _6205_ (.A(_2580_),
    .B(_2581_),
    .X(_2582_));
 sky130_fd_sc_hd__clkbuf_1 _6206_ (.A(_2582_),
    .X(_0188_));
 sky130_fd_sc_hd__mux2_1 _6207_ (.A0(net10),
    .A1(_3353_),
    .S(net197),
    .X(_2583_));
 sky130_fd_sc_hd__and2_1 _6208_ (.A(_2583_),
    .B(_2581_),
    .X(_2584_));
 sky130_fd_sc_hd__clkbuf_1 _6209_ (.A(_2584_),
    .X(_0187_));
 sky130_fd_sc_hd__mux2_1 _6210_ (.A0(net9),
    .A1(_3357_),
    .S(net197),
    .X(_2585_));
 sky130_fd_sc_hd__and2_1 _6211_ (.A(_2585_),
    .B(_2581_),
    .X(_2586_));
 sky130_fd_sc_hd__clkbuf_1 _6212_ (.A(_2586_),
    .X(_0186_));
 sky130_fd_sc_hd__mux2_1 _6213_ (.A0(net8),
    .A1(_0674_),
    .S(net197),
    .X(_2587_));
 sky130_fd_sc_hd__and2_1 _6214_ (.A(_2587_),
    .B(_2581_),
    .X(_2588_));
 sky130_fd_sc_hd__clkbuf_1 _6215_ (.A(_2588_),
    .X(_0185_));
 sky130_fd_sc_hd__mux2_1 _6216_ (.A0(net1),
    .A1(_0675_),
    .S(net197),
    .X(_2589_));
 sky130_fd_sc_hd__and2_1 _6217_ (.A(_2589_),
    .B(_2581_),
    .X(_2590_));
 sky130_fd_sc_hd__clkbuf_1 _6218_ (.A(_2590_),
    .X(_0184_));
 sky130_fd_sc_hd__or2_1 _6219_ (.A(\egd_top.BitStream_buffer.pc_previous[1] ),
    .B(\egd_top.BitStream_buffer.exp_golomb_len[1] ),
    .X(_2591_));
 sky130_fd_sc_hd__nand2_2 _6220_ (.A(\egd_top.BitStream_buffer.pc_previous[1] ),
    .B(\egd_top.BitStream_buffer.exp_golomb_len[1] ),
    .Y(_2592_));
 sky130_fd_sc_hd__nand2_2 _6221_ (.A(_2591_),
    .B(_2592_),
    .Y(_2593_));
 sky130_fd_sc_hd__o21ai_4 _6222_ (.A1(_2960_),
    .A2(_2593_),
    .B1(_2592_),
    .Y(_2594_));
 sky130_fd_sc_hd__or2_1 _6223_ (.A(\egd_top.BitStream_buffer.pc_previous[2] ),
    .B(\egd_top.BitStream_buffer.exp_golomb_len[2] ),
    .X(_2595_));
 sky130_fd_sc_hd__nand2_1 _6224_ (.A(\egd_top.BitStream_buffer.pc_previous[2] ),
    .B(\egd_top.BitStream_buffer.exp_golomb_len[2] ),
    .Y(_2596_));
 sky130_fd_sc_hd__a21bo_2 _6225_ (.A1(_2594_),
    .A2(_2595_),
    .B1_N(_2596_),
    .X(_2597_));
 sky130_fd_sc_hd__or2_1 _6226_ (.A(\egd_top.BitStream_buffer.pc_previous[3] ),
    .B(\egd_top.BitStream_buffer.exp_golomb_len[3] ),
    .X(_2598_));
 sky130_fd_sc_hd__nand2_1 _6227_ (.A(\egd_top.BitStream_buffer.pc_previous[3] ),
    .B(\egd_top.BitStream_buffer.exp_golomb_len[3] ),
    .Y(_2599_));
 sky130_fd_sc_hd__a21bo_2 _6228_ (.A1(_2597_),
    .A2(_2598_),
    .B1_N(_2599_),
    .X(_2600_));
 sky130_fd_sc_hd__and3_2 _6229_ (.A(_2600_),
    .B(\egd_top.BitStream_buffer.pc_previous[4] ),
    .C(\egd_top.BitStream_buffer.pc_previous[5] ),
    .X(_2601_));
 sky130_fd_sc_hd__xor2_4 _6230_ (.A(\egd_top.BitStream_buffer.pc_previous[6] ),
    .B(_2601_),
    .X(\egd_top.BitStream_buffer.pc[6] ));
 sky130_fd_sc_hd__nand2_1 _6231_ (.A(_2989_),
    .B(\egd_top.BitStream_buffer.pc[6] ),
    .Y(_2602_));
 sky130_fd_sc_hd__inv_2 _6232_ (.A(_2602_),
    .Y(_0183_));
 sky130_fd_sc_hd__a21oi_1 _6233_ (.A1(_2600_),
    .A2(\egd_top.BitStream_buffer.pc_previous[4] ),
    .B1(\egd_top.BitStream_buffer.pc_previous[5] ),
    .Y(_2603_));
 sky130_fd_sc_hd__nor2_2 _6234_ (.A(_2603_),
    .B(_2601_),
    .Y(\egd_top.BitStream_buffer.pc[5] ));
 sky130_fd_sc_hd__nand2_1 _6235_ (.A(_2989_),
    .B(\egd_top.BitStream_buffer.pc[5] ),
    .Y(_2604_));
 sky130_fd_sc_hd__inv_2 _6236_ (.A(_2604_),
    .Y(_0182_));
 sky130_fd_sc_hd__xor2_4 _6237_ (.A(\egd_top.BitStream_buffer.pc_previous[4] ),
    .B(_2600_),
    .X(\egd_top.BitStream_buffer.pc[4] ));
 sky130_fd_sc_hd__nand2_1 _6238_ (.A(_2989_),
    .B(\egd_top.BitStream_buffer.pc[4] ),
    .Y(_2605_));
 sky130_fd_sc_hd__inv_2 _6239_ (.A(_2605_),
    .Y(_0181_));
 sky130_fd_sc_hd__nand2_2 _6240_ (.A(_2598_),
    .B(_2599_),
    .Y(_2606_));
 sky130_fd_sc_hd__xnor2_4 _6241_ (.A(_2606_),
    .B(_2597_),
    .Y(\egd_top.BitStream_buffer.pc[3] ));
 sky130_fd_sc_hd__nand2_1 _6242_ (.A(_2989_),
    .B(\egd_top.BitStream_buffer.pc[3] ),
    .Y(_2607_));
 sky130_fd_sc_hd__inv_2 _6243_ (.A(_2607_),
    .Y(_0180_));
 sky130_fd_sc_hd__nand2_2 _6244_ (.A(_2595_),
    .B(_2596_),
    .Y(_2608_));
 sky130_fd_sc_hd__xnor2_4 _6245_ (.A(_2608_),
    .B(_2594_),
    .Y(\egd_top.BitStream_buffer.pc[2] ));
 sky130_fd_sc_hd__nand2_1 _6246_ (.A(_2989_),
    .B(\egd_top.BitStream_buffer.pc[2] ),
    .Y(_2609_));
 sky130_fd_sc_hd__inv_2 _6247_ (.A(_2609_),
    .Y(_0179_));
 sky130_fd_sc_hd__xor2_4 _6248_ (.A(_2960_),
    .B(_2593_),
    .X(\egd_top.BitStream_buffer.pc[1] ));
 sky130_fd_sc_hd__nand2_1 _6249_ (.A(_2989_),
    .B(\egd_top.BitStream_buffer.pc[1] ),
    .Y(_2610_));
 sky130_fd_sc_hd__inv_2 _6250_ (.A(_2610_),
    .Y(_0178_));
 sky130_fd_sc_hd__nand2_1 _6251_ (.A(_2962_),
    .B(_2989_),
    .Y(_2611_));
 sky130_fd_sc_hd__inv_2 _6252_ (.A(_2611_),
    .Y(_0177_));
 sky130_fd_sc_hd__or4b_4 _6253_ (.A(_2978_),
    .B(net198),
    .C(_2972_),
    .D_N(_3002_),
    .X(_2612_));
 sky130_fd_sc_hd__buf_4 _6254_ (.A(_2612_),
    .X(_2613_));
 sky130_fd_sc_hd__mux2_1 _6255_ (.A0(net7),
    .A1(_3255_),
    .S(_2613_),
    .X(_2614_));
 sky130_fd_sc_hd__and2_1 _6256_ (.A(_2614_),
    .B(_2581_),
    .X(_2615_));
 sky130_fd_sc_hd__clkbuf_1 _6257_ (.A(_2615_),
    .X(_0176_));
 sky130_fd_sc_hd__mux2_1 _6258_ (.A0(net6),
    .A1(_3247_),
    .S(_2613_),
    .X(_2616_));
 sky130_fd_sc_hd__and2_1 _6259_ (.A(_2616_),
    .B(_2581_),
    .X(_2617_));
 sky130_fd_sc_hd__clkbuf_1 _6260_ (.A(_2617_),
    .X(_0175_));
 sky130_fd_sc_hd__mux2_1 _6261_ (.A0(net5),
    .A1(_3259_),
    .S(_2613_),
    .X(_2618_));
 sky130_fd_sc_hd__and2_1 _6262_ (.A(_2618_),
    .B(_2581_),
    .X(_2619_));
 sky130_fd_sc_hd__clkbuf_1 _6263_ (.A(_2619_),
    .X(_0174_));
 sky130_fd_sc_hd__mux2_1 _6264_ (.A0(net4),
    .A1(_3251_),
    .S(_2613_),
    .X(_2620_));
 sky130_fd_sc_hd__and2_1 _6265_ (.A(_2620_),
    .B(_2581_),
    .X(_2621_));
 sky130_fd_sc_hd__clkbuf_1 _6266_ (.A(_2621_),
    .X(_0173_));
 sky130_fd_sc_hd__mux2_1 _6267_ (.A0(net3),
    .A1(_0646_),
    .S(_2613_),
    .X(_2622_));
 sky130_fd_sc_hd__and2_1 _6268_ (.A(_2622_),
    .B(_2581_),
    .X(_2623_));
 sky130_fd_sc_hd__clkbuf_1 _6269_ (.A(_2623_),
    .X(_0172_));
 sky130_fd_sc_hd__mux2_1 _6270_ (.A0(net2),
    .A1(_3265_),
    .S(_2613_),
    .X(_2624_));
 sky130_fd_sc_hd__and2_1 _6271_ (.A(_2624_),
    .B(_2581_),
    .X(_2625_));
 sky130_fd_sc_hd__clkbuf_1 _6272_ (.A(_2625_),
    .X(_0171_));
 sky130_fd_sc_hd__mux2_1 _6273_ (.A0(net16),
    .A1(_3272_),
    .S(_2613_),
    .X(_2626_));
 sky130_fd_sc_hd__and2_1 _6274_ (.A(_2626_),
    .B(_2581_),
    .X(_2627_));
 sky130_fd_sc_hd__clkbuf_1 _6275_ (.A(_2627_),
    .X(_0170_));
 sky130_fd_sc_hd__mux2_1 _6276_ (.A0(net15),
    .A1(_3275_),
    .S(_2613_),
    .X(_2628_));
 sky130_fd_sc_hd__and2_1 _6277_ (.A(_2628_),
    .B(_2372_),
    .X(_2629_));
 sky130_fd_sc_hd__clkbuf_1 _6278_ (.A(_2629_),
    .X(_0169_));
 sky130_fd_sc_hd__mux2_1 _6279_ (.A0(net14),
    .A1(_0653_),
    .S(_2613_),
    .X(_2630_));
 sky130_fd_sc_hd__and2_1 _6280_ (.A(_2630_),
    .B(_2372_),
    .X(_2631_));
 sky130_fd_sc_hd__clkbuf_1 _6281_ (.A(_2631_),
    .X(_0168_));
 sky130_fd_sc_hd__mux2_1 _6282_ (.A0(net13),
    .A1(_0804_),
    .S(_2613_),
    .X(_2632_));
 sky130_fd_sc_hd__and2_1 _6283_ (.A(_2632_),
    .B(_2372_),
    .X(_2633_));
 sky130_fd_sc_hd__clkbuf_1 _6284_ (.A(_2633_),
    .X(_0167_));
 sky130_fd_sc_hd__mux2_1 _6285_ (.A0(net12),
    .A1(_3225_),
    .S(_2613_),
    .X(_2634_));
 sky130_fd_sc_hd__and2_1 _6286_ (.A(_2634_),
    .B(_2372_),
    .X(_2635_));
 sky130_fd_sc_hd__clkbuf_1 _6287_ (.A(_2635_),
    .X(_0166_));
 sky130_fd_sc_hd__mux2_1 _6288_ (.A0(net11),
    .A1(_3232_),
    .S(_2613_),
    .X(_2636_));
 sky130_fd_sc_hd__and2_1 _6289_ (.A(_2636_),
    .B(_2372_),
    .X(_2637_));
 sky130_fd_sc_hd__clkbuf_1 _6290_ (.A(_2637_),
    .X(_0165_));
 sky130_fd_sc_hd__mux2_1 _6291_ (.A0(net10),
    .A1(_3286_),
    .S(net199),
    .X(_2638_));
 sky130_fd_sc_hd__and2_1 _6292_ (.A(_2638_),
    .B(_2372_),
    .X(_2639_));
 sky130_fd_sc_hd__clkbuf_1 _6293_ (.A(_2639_),
    .X(_0164_));
 sky130_fd_sc_hd__mux2_1 _6294_ (.A0(net9),
    .A1(_3290_),
    .S(net199),
    .X(_2640_));
 sky130_fd_sc_hd__and2_1 _6295_ (.A(_2640_),
    .B(_2372_),
    .X(_2641_));
 sky130_fd_sc_hd__clkbuf_1 _6296_ (.A(_2641_),
    .X(_0163_));
 sky130_fd_sc_hd__mux2_1 _6297_ (.A0(net8),
    .A1(_3278_),
    .S(net199),
    .X(_2642_));
 sky130_fd_sc_hd__and2_1 _6298_ (.A(_2642_),
    .B(_2372_),
    .X(_2643_));
 sky130_fd_sc_hd__clkbuf_1 _6299_ (.A(_2643_),
    .X(_0162_));
 sky130_fd_sc_hd__mux2_1 _6300_ (.A0(net1),
    .A1(_3282_),
    .S(net199),
    .X(_2644_));
 sky130_fd_sc_hd__and2_1 _6301_ (.A(_2644_),
    .B(_2372_),
    .X(_2645_));
 sky130_fd_sc_hd__clkbuf_1 _6302_ (.A(_2645_),
    .X(_0161_));
 sky130_fd_sc_hd__nand2_1 _6303_ (.A(net18),
    .B(net17),
    .Y(_2646_));
 sky130_fd_sc_hd__inv_2 _6304_ (.A(_2646_),
    .Y(_2647_));
 sky130_fd_sc_hd__and3b_1 _6305_ (.A_N(net21),
    .B(_2647_),
    .C(net20),
    .X(_2648_));
 sky130_fd_sc_hd__inv_2 _6306_ (.A(\egd_top.exp_golomb_decoding.te_range[2] ),
    .Y(_2649_));
 sky130_fd_sc_hd__and2_2 _6307_ (.A(_2648_),
    .B(_2649_),
    .X(_2650_));
 sky130_fd_sc_hd__nor2_1 _6308_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[15] ),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[14] ),
    .Y(_2651_));
 sky130_fd_sc_hd__nand2_1 _6309_ (.A(_2651_),
    .B(_2997_),
    .Y(_2652_));
 sky130_fd_sc_hd__nand2_1 _6310_ (.A(_1029_),
    .B(_1157_),
    .Y(_2653_));
 sky130_fd_sc_hd__nor2_1 _6311_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[13] ),
    .B(_2653_),
    .Y(_2654_));
 sky130_fd_sc_hd__nand2_1 _6312_ (.A(_2654_),
    .B(_1282_),
    .Y(_2655_));
 sky130_fd_sc_hd__inv_2 _6313_ (.A(_2655_),
    .Y(_2656_));
 sky130_fd_sc_hd__and3_1 _6314_ (.A(_2656_),
    .B(_1406_),
    .C(_1530_),
    .X(_2657_));
 sky130_fd_sc_hd__inv_2 _6315_ (.A(_2657_),
    .Y(_2658_));
 sky130_fd_sc_hd__nor2_1 _6316_ (.A(_2652_),
    .B(_2658_),
    .Y(_2659_));
 sky130_fd_sc_hd__nor2_1 _6317_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[6] ),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[5] ),
    .Y(_2660_));
 sky130_fd_sc_hd__inv_2 _6318_ (.A(_2660_),
    .Y(_2661_));
 sky130_fd_sc_hd__nor2_1 _6319_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[7] ),
    .B(_2661_),
    .Y(_2662_));
 sky130_fd_sc_hd__nand2_1 _6320_ (.A(_2662_),
    .B(_2013_),
    .Y(_2663_));
 sky130_fd_sc_hd__inv_2 _6321_ (.A(_2652_),
    .Y(_2664_));
 sky130_fd_sc_hd__nor2_1 _6322_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[13] ),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[12] ),
    .Y(_2665_));
 sky130_fd_sc_hd__nand2_2 _6323_ (.A(_2664_),
    .B(_2665_),
    .Y(_2666_));
 sky130_fd_sc_hd__a21o_1 _6324_ (.A1(_2657_),
    .A2(_2663_),
    .B1(_2666_),
    .X(_2667_));
 sky130_fd_sc_hd__nor2_2 _6325_ (.A(_2659_),
    .B(_2667_),
    .Y(_2668_));
 sky130_fd_sc_hd__inv_6 _6326_ (.A(_2668_),
    .Y(_2669_));
 sky130_fd_sc_hd__nand2_1 _6327_ (.A(_2251_),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[1] ),
    .Y(_2670_));
 sky130_fd_sc_hd__nand2_1 _6328_ (.A(_2670_),
    .B(_2132_),
    .Y(_2671_));
 sky130_fd_sc_hd__nand2_1 _6329_ (.A(_2671_),
    .B(_2013_),
    .Y(_2672_));
 sky130_fd_sc_hd__nand2_1 _6330_ (.A(_2672_),
    .B(_1894_),
    .Y(_2673_));
 sky130_fd_sc_hd__nand2_1 _6331_ (.A(_2673_),
    .B(_1774_),
    .Y(_2674_));
 sky130_fd_sc_hd__nand2_1 _6332_ (.A(_2674_),
    .B(_1652_),
    .Y(_2675_));
 sky130_fd_sc_hd__nand2_1 _6333_ (.A(_2675_),
    .B(_1530_),
    .Y(_2676_));
 sky130_fd_sc_hd__nand2_1 _6334_ (.A(_2676_),
    .B(_1406_),
    .Y(_2677_));
 sky130_fd_sc_hd__nand2_1 _6335_ (.A(_2677_),
    .B(_2656_),
    .Y(_2678_));
 sky130_fd_sc_hd__a21oi_1 _6336_ (.A1(_1029_),
    .A2(\egd_top.BitStream_buffer.BitStream_buffer_output[11] ),
    .B1(\egd_top.BitStream_buffer.BitStream_buffer_output[13] ),
    .Y(_2679_));
 sky130_fd_sc_hd__nand2_1 _6337_ (.A(_2678_),
    .B(_2679_),
    .Y(_2680_));
 sky130_fd_sc_hd__nand2_2 _6338_ (.A(_2680_),
    .B(_2651_),
    .Y(_2681_));
 sky130_fd_sc_hd__o21ai_1 _6339_ (.A1(\egd_top.BitStream_buffer.BitStream_buffer_output[3] ),
    .A2(\egd_top.BitStream_buffer.BitStream_buffer_output[2] ),
    .B1(_2013_),
    .Y(_2682_));
 sky130_fd_sc_hd__o211a_1 _6340_ (.A1(\egd_top.BitStream_buffer.BitStream_buffer_output[5] ),
    .A2(_2682_),
    .B1(_1652_),
    .C1(_1774_),
    .X(_2683_));
 sky130_fd_sc_hd__a21o_1 _6341_ (.A1(_2655_),
    .A2(_2665_),
    .B1(_2652_),
    .X(_2684_));
 sky130_fd_sc_hd__o21bai_4 _6342_ (.A1(_2683_),
    .A2(_2658_),
    .B1_N(_2684_),
    .Y(_2685_));
 sky130_fd_sc_hd__nor2_2 _6343_ (.A(_2996_),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[15] ),
    .Y(_2686_));
 sky130_fd_sc_hd__nand3_1 _6344_ (.A(_2681_),
    .B(_2685_),
    .C(_2686_),
    .Y(_2687_));
 sky130_fd_sc_hd__nor2_2 _6345_ (.A(_2669_),
    .B(_2687_),
    .Y(_2688_));
 sky130_fd_sc_hd__clkinvlp_2 _6346_ (.A(_2688_),
    .Y(_2689_));
 sky130_fd_sc_hd__nor2_1 _6347_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[5] ),
    .B(_2689_),
    .Y(_2690_));
 sky130_fd_sc_hd__inv_4 _6348_ (.A(_2685_),
    .Y(_2691_));
 sky130_fd_sc_hd__nor2_1 _6349_ (.A(_2691_),
    .B(_2669_),
    .Y(_2692_));
 sky130_fd_sc_hd__nand2_2 _6350_ (.A(_2681_),
    .B(_2686_),
    .Y(_2693_));
 sky130_fd_sc_hd__nand2_1 _6351_ (.A(_2692_),
    .B(_2693_),
    .Y(_2694_));
 sky130_fd_sc_hd__nand2_1 _6352_ (.A(_2691_),
    .B(_2666_),
    .Y(_2695_));
 sky130_fd_sc_hd__inv_2 _6353_ (.A(_2695_),
    .Y(_2696_));
 sky130_fd_sc_hd__nand3_1 _6354_ (.A(_2696_),
    .B(_2693_),
    .C(_1157_),
    .Y(_2697_));
 sky130_fd_sc_hd__o21ai_1 _6355_ (.A1(\egd_top.BitStream_buffer.BitStream_buffer_output[7] ),
    .A2(_2694_),
    .B1(_2697_),
    .Y(_2698_));
 sky130_fd_sc_hd__nor2_1 _6356_ (.A(_2690_),
    .B(_2698_),
    .Y(_2699_));
 sky130_fd_sc_hd__nand3_4 _6357_ (.A(_2681_),
    .B(_2691_),
    .C(_2686_),
    .Y(_2700_));
 sky130_fd_sc_hd__inv_2 _6358_ (.A(_2700_),
    .Y(_2701_));
 sky130_fd_sc_hd__and3_1 _6359_ (.A(_2701_),
    .B(_1406_),
    .C(_2666_),
    .X(_2702_));
 sky130_fd_sc_hd__inv_2 _6360_ (.A(_2687_),
    .Y(_2703_));
 sky130_fd_sc_hd__and3_1 _6361_ (.A(_2703_),
    .B(_0897_),
    .C(_2666_),
    .X(_2704_));
 sky130_fd_sc_hd__nor2_1 _6362_ (.A(_2702_),
    .B(_2704_),
    .Y(_2705_));
 sky130_fd_sc_hd__o21ai_1 _6363_ (.A1(_2669_),
    .A2(_2700_),
    .B1(_2132_),
    .Y(_2706_));
 sky130_fd_sc_hd__nor2_4 _6364_ (.A(_2669_),
    .B(_2700_),
    .Y(_2707_));
 sky130_fd_sc_hd__nand2_1 _6365_ (.A(_2707_),
    .B(_2370_),
    .Y(_2708_));
 sky130_fd_sc_hd__nand2_2 _6366_ (.A(_2706_),
    .B(_2708_),
    .Y(_2709_));
 sky130_fd_sc_hd__nor2_2 _6367_ (.A(_2685_),
    .B(_2669_),
    .Y(_2710_));
 sky130_fd_sc_hd__nand2_1 _6368_ (.A(_2709_),
    .B(_2710_),
    .Y(_2711_));
 sky130_fd_sc_hd__nand3_2 _6369_ (.A(_2699_),
    .B(_2705_),
    .C(_2711_),
    .Y(_2712_));
 sky130_fd_sc_hd__nand2_2 _6370_ (.A(_2712_),
    .B(_2959_),
    .Y(_2713_));
 sky130_fd_sc_hd__inv_2 _6371_ (.A(_2713_),
    .Y(_2714_));
 sky130_fd_sc_hd__or2_1 _6372_ (.A(_2650_),
    .B(_2714_),
    .X(_2715_));
 sky130_fd_sc_hd__inv_2 _6373_ (.A(_2959_),
    .Y(_2716_));
 sky130_fd_sc_hd__a311o_1 _6374_ (.A1(_2693_),
    .A2(_2667_),
    .A3(_2685_),
    .B1(_2716_),
    .C1(_2659_),
    .X(_2717_));
 sky130_fd_sc_hd__nand2_1 _6375_ (.A(_2717_),
    .B(_2650_),
    .Y(_2718_));
 sky130_fd_sc_hd__nor2_1 _6376_ (.A(net18),
    .B(_2956_),
    .Y(_2719_));
 sky130_fd_sc_hd__nand2_1 _6377_ (.A(_2701_),
    .B(_2668_),
    .Y(_2720_));
 sky130_fd_sc_hd__nand2_1 _6378_ (.A(_2720_),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[3] ),
    .Y(_2721_));
 sky130_fd_sc_hd__nand2_1 _6379_ (.A(_2707_),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[1] ),
    .Y(_2722_));
 sky130_fd_sc_hd__nand2_1 _6380_ (.A(_2721_),
    .B(_2722_),
    .Y(_2723_));
 sky130_fd_sc_hd__o21ai_1 _6381_ (.A1(_2669_),
    .A2(_2700_),
    .B1(_2013_),
    .Y(_2724_));
 sky130_fd_sc_hd__nand3_1 _6382_ (.A(_2701_),
    .B(_2251_),
    .C(_2668_),
    .Y(_2725_));
 sky130_fd_sc_hd__nand2_1 _6383_ (.A(_2724_),
    .B(_2725_),
    .Y(_2726_));
 sky130_fd_sc_hd__nand2_1 _6384_ (.A(_2723_),
    .B(_2726_),
    .Y(_2727_));
 sky130_fd_sc_hd__o21ai_1 _6385_ (.A1(_2669_),
    .A2(_2700_),
    .B1(\egd_top.BitStream_buffer.BitStream_buffer_output[4] ),
    .Y(_2728_));
 sky130_fd_sc_hd__nand3_1 _6386_ (.A(_2701_),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[2] ),
    .C(_2668_),
    .Y(_2729_));
 sky130_fd_sc_hd__nand2_1 _6387_ (.A(_2728_),
    .B(_2729_),
    .Y(_2730_));
 sky130_fd_sc_hd__nand2_1 _6388_ (.A(_2709_),
    .B(_2730_),
    .Y(_2731_));
 sky130_fd_sc_hd__nand3_1 _6389_ (.A(_2727_),
    .B(_2731_),
    .C(_2710_),
    .Y(_2732_));
 sky130_fd_sc_hd__and2_1 _6390_ (.A(_2701_),
    .B(_2666_),
    .X(_2733_));
 sky130_fd_sc_hd__nor2_1 _6391_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[10] ),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[9] ),
    .Y(_2734_));
 sky130_fd_sc_hd__inv_2 _6392_ (.A(_2734_),
    .Y(_2735_));
 sky130_fd_sc_hd__nand2_1 _6393_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[10] ),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[9] ),
    .Y(_2736_));
 sky130_fd_sc_hd__nand2_1 _6394_ (.A(_2735_),
    .B(_2736_),
    .Y(_2737_));
 sky130_fd_sc_hd__nand2_1 _6395_ (.A(_2733_),
    .B(_2737_),
    .Y(_2738_));
 sky130_fd_sc_hd__xnor2_1 _6396_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[14] ),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[13] ),
    .Y(_2739_));
 sky130_fd_sc_hd__nand3_1 _6397_ (.A(_2703_),
    .B(_2666_),
    .C(_2739_),
    .Y(_2740_));
 sky130_fd_sc_hd__nand2_1 _6398_ (.A(_2738_),
    .B(_2740_),
    .Y(_2741_));
 sky130_fd_sc_hd__xor2_1 _6399_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[12] ),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[11] ),
    .X(_2742_));
 sky130_fd_sc_hd__nand2_1 _6400_ (.A(_2696_),
    .B(_2693_),
    .Y(_2743_));
 sky130_fd_sc_hd__nor2_1 _6401_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[8] ),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[7] ),
    .Y(_2744_));
 sky130_fd_sc_hd__inv_2 _6402_ (.A(_2744_),
    .Y(_2745_));
 sky130_fd_sc_hd__nand2_1 _6403_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[8] ),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[7] ),
    .Y(_2746_));
 sky130_fd_sc_hd__nand2_1 _6404_ (.A(_2745_),
    .B(_2746_),
    .Y(_2747_));
 sky130_fd_sc_hd__nand3_1 _6405_ (.A(_2692_),
    .B(_2693_),
    .C(_2747_),
    .Y(_2748_));
 sky130_fd_sc_hd__nand2_1 _6406_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[6] ),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[5] ),
    .Y(_2749_));
 sky130_fd_sc_hd__nand2_1 _6407_ (.A(_2661_),
    .B(_2749_),
    .Y(_2750_));
 sky130_fd_sc_hd__nand2_1 _6408_ (.A(_2688_),
    .B(_2750_),
    .Y(_2751_));
 sky130_fd_sc_hd__o211ai_1 _6409_ (.A1(_2742_),
    .A2(_2743_),
    .B1(_2748_),
    .C1(_2751_),
    .Y(_2752_));
 sky130_fd_sc_hd__nor2_1 _6410_ (.A(_2741_),
    .B(_2752_),
    .Y(_2753_));
 sky130_fd_sc_hd__nand2_1 _6411_ (.A(_2732_),
    .B(_2753_),
    .Y(_2754_));
 sky130_fd_sc_hd__nand3_1 _6412_ (.A(_2754_),
    .B(_2959_),
    .C(_2712_),
    .Y(_2755_));
 sky130_fd_sc_hd__nor2_2 _6413_ (.A(net17),
    .B(_2955_),
    .Y(_2756_));
 sky130_fd_sc_hd__a22o_1 _6414_ (.A1(_2714_),
    .A2(_2719_),
    .B1(_2755_),
    .B2(_2756_),
    .X(_2757_));
 sky130_fd_sc_hd__nand2_2 _6415_ (.A(_2754_),
    .B(_2959_),
    .Y(_2758_));
 sky130_fd_sc_hd__nand2_1 _6416_ (.A(_2758_),
    .B(_2713_),
    .Y(_2759_));
 sky130_fd_sc_hd__a32o_2 _6417_ (.A1(_2647_),
    .A2(_2715_),
    .A3(_2718_),
    .B1(_2757_),
    .B2(_2759_),
    .X(net20));
 sky130_fd_sc_hd__a31o_1 _6418_ (.A1(_2648_),
    .A2(net18),
    .A3(_2649_),
    .B1(_2956_),
    .X(_2760_));
 sky130_fd_sc_hd__nand2_1 _6419_ (.A(_2709_),
    .B(_2726_),
    .Y(_2761_));
 sky130_fd_sc_hd__o21ai_1 _6420_ (.A1(_2669_),
    .A2(_2700_),
    .B1(_1894_),
    .Y(_2762_));
 sky130_fd_sc_hd__nand2_1 _6421_ (.A(_2707_),
    .B(_2132_),
    .Y(_2763_));
 sky130_fd_sc_hd__nand2_1 _6422_ (.A(_2762_),
    .B(_2763_),
    .Y(_2764_));
 sky130_fd_sc_hd__nand2_1 _6423_ (.A(_2761_),
    .B(_2764_),
    .Y(_2765_));
 sky130_fd_sc_hd__o21ai_1 _6424_ (.A1(_2669_),
    .A2(_2700_),
    .B1(\egd_top.BitStream_buffer.BitStream_buffer_output[5] ),
    .Y(_2766_));
 sky130_fd_sc_hd__nand2_1 _6425_ (.A(_2707_),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[3] ),
    .Y(_2767_));
 sky130_fd_sc_hd__nand2_1 _6426_ (.A(_2766_),
    .B(_2767_),
    .Y(_2768_));
 sky130_fd_sc_hd__nand3_1 _6427_ (.A(_2709_),
    .B(_2768_),
    .C(_2726_),
    .Y(_2769_));
 sky130_fd_sc_hd__nand3_1 _6428_ (.A(_2765_),
    .B(_2769_),
    .C(_2710_),
    .Y(_2770_));
 sky130_fd_sc_hd__nor2_1 _6429_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[11] ),
    .B(_2735_),
    .Y(_2771_));
 sky130_fd_sc_hd__nor2_1 _6430_ (.A(_1157_),
    .B(_2734_),
    .Y(_2772_));
 sky130_fd_sc_hd__o21ai_1 _6431_ (.A1(_2771_),
    .A2(_2772_),
    .B1(_2733_),
    .Y(_2773_));
 sky130_fd_sc_hd__nor2_1 _6432_ (.A(_1652_),
    .B(_2660_),
    .Y(_2774_));
 sky130_fd_sc_hd__o21ai_1 _6433_ (.A1(_2662_),
    .A2(_2774_),
    .B1(_2688_),
    .Y(_2775_));
 sky130_fd_sc_hd__nand2_1 _6434_ (.A(_2773_),
    .B(_2775_),
    .Y(_2776_));
 sky130_fd_sc_hd__and2_1 _6435_ (.A(_2653_),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[13] ),
    .X(_2777_));
 sky130_fd_sc_hd__nor2_1 _6436_ (.A(_2654_),
    .B(_2777_),
    .Y(_2778_));
 sky130_fd_sc_hd__nor2_1 _6437_ (.A(_1406_),
    .B(_2744_),
    .Y(_2779_));
 sky130_fd_sc_hd__nor2_1 _6438_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[9] ),
    .B(_2745_),
    .Y(_2780_));
 sky130_fd_sc_hd__inv_2 _6439_ (.A(_2694_),
    .Y(_2781_));
 sky130_fd_sc_hd__o21ai_1 _6440_ (.A1(_2779_),
    .A2(_2780_),
    .B1(_2781_),
    .Y(_2782_));
 sky130_fd_sc_hd__o21ai_1 _6441_ (.A1(_2743_),
    .A2(_2778_),
    .B1(_2782_),
    .Y(_2783_));
 sky130_fd_sc_hd__nor2_1 _6442_ (.A(_2776_),
    .B(_2783_),
    .Y(_2784_));
 sky130_fd_sc_hd__nand2_1 _6443_ (.A(_2770_),
    .B(_2784_),
    .Y(_2785_));
 sky130_fd_sc_hd__nand2_2 _6444_ (.A(_2785_),
    .B(_2959_),
    .Y(_2786_));
 sky130_fd_sc_hd__or2_1 _6445_ (.A(_2758_),
    .B(_2786_),
    .X(_2787_));
 sky130_fd_sc_hd__nand2_2 _6446_ (.A(_2786_),
    .B(_2758_),
    .Y(_2788_));
 sky130_fd_sc_hd__nand3_1 _6447_ (.A(_2787_),
    .B(_2788_),
    .C(_2756_),
    .Y(_2789_));
 sky130_fd_sc_hd__o21ai_2 _6448_ (.A1(_2758_),
    .A2(_2760_),
    .B1(_2789_),
    .Y(net21));
 sky130_fd_sc_hd__o21ai_1 _6449_ (.A1(_2758_),
    .A2(_2786_),
    .B1(_2714_),
    .Y(_2790_));
 sky130_fd_sc_hd__nand2_1 _6450_ (.A(_2790_),
    .B(_2788_),
    .Y(_2791_));
 sky130_fd_sc_hd__nor2_1 _6451_ (.A(_2730_),
    .B(_2723_),
    .Y(_2792_));
 sky130_fd_sc_hd__nand2_1 _6452_ (.A(_2707_),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[4] ),
    .Y(_2793_));
 sky130_fd_sc_hd__o21ai_1 _6453_ (.A1(_1774_),
    .A2(_2707_),
    .B1(_2793_),
    .Y(_2794_));
 sky130_fd_sc_hd__nand3_1 _6454_ (.A(_2792_),
    .B(_2794_),
    .C(_2764_),
    .Y(_2795_));
 sky130_fd_sc_hd__nand3_1 _6455_ (.A(_2709_),
    .B(_2764_),
    .C(_2726_),
    .Y(_2796_));
 sky130_fd_sc_hd__nand2_1 _6456_ (.A(_2707_),
    .B(_2013_),
    .Y(_2797_));
 sky130_fd_sc_hd__o21ai_1 _6457_ (.A1(\egd_top.BitStream_buffer.BitStream_buffer_output[6] ),
    .A2(_2707_),
    .B1(_2797_),
    .Y(_2798_));
 sky130_fd_sc_hd__nand2_1 _6458_ (.A(_2796_),
    .B(_2798_),
    .Y(_2799_));
 sky130_fd_sc_hd__nand3_1 _6459_ (.A(_2795_),
    .B(_2799_),
    .C(_2710_),
    .Y(_2800_));
 sky130_fd_sc_hd__nand2_1 _6460_ (.A(_2771_),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[12] ),
    .Y(_2801_));
 sky130_fd_sc_hd__or2_1 _6461_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[12] ),
    .B(_2771_),
    .X(_2802_));
 sky130_fd_sc_hd__and3_1 _6462_ (.A(_2733_),
    .B(_2801_),
    .C(_2802_),
    .X(_2803_));
 sky130_fd_sc_hd__or2_1 _6463_ (.A(_1530_),
    .B(_2662_),
    .X(_2804_));
 sky130_fd_sc_hd__nor2_1 _6464_ (.A(_2661_),
    .B(_2745_),
    .Y(_2805_));
 sky130_fd_sc_hd__inv_2 _6465_ (.A(_2805_),
    .Y(_2806_));
 sky130_fd_sc_hd__nand2_1 _6466_ (.A(_2804_),
    .B(_2806_),
    .Y(_2807_));
 sky130_fd_sc_hd__mux2_1 _6467_ (.A0(\egd_top.BitStream_buffer.BitStream_buffer_output[10] ),
    .A1(_2737_),
    .S(_2744_),
    .X(_2808_));
 sky130_fd_sc_hd__a22o_1 _6468_ (.A1(_2688_),
    .A2(_2807_),
    .B1(_2781_),
    .B2(_2808_),
    .X(_2809_));
 sky130_fd_sc_hd__nor2_1 _6469_ (.A(_2803_),
    .B(_2809_),
    .Y(_2810_));
 sky130_fd_sc_hd__a21oi_1 _6470_ (.A1(_2800_),
    .A2(_2810_),
    .B1(_2716_),
    .Y(_2811_));
 sky130_fd_sc_hd__nand2_1 _6471_ (.A(_2791_),
    .B(_2811_),
    .Y(_2812_));
 sky130_fd_sc_hd__nand2_1 _6472_ (.A(_2800_),
    .B(_2810_),
    .Y(_2813_));
 sky130_fd_sc_hd__nand2_1 _6473_ (.A(_2813_),
    .B(_2959_),
    .Y(_2814_));
 sky130_fd_sc_hd__nand3_1 _6474_ (.A(_2790_),
    .B(_2788_),
    .C(_2814_),
    .Y(_2815_));
 sky130_fd_sc_hd__nand2_1 _6475_ (.A(_2812_),
    .B(_2815_),
    .Y(_2816_));
 sky130_fd_sc_hd__nand2_1 _6476_ (.A(_2816_),
    .B(_2756_),
    .Y(_2817_));
 sky130_fd_sc_hd__or2_1 _6477_ (.A(_2760_),
    .B(_2786_),
    .X(_2818_));
 sky130_fd_sc_hd__nand2_1 _6478_ (.A(net20),
    .B(net21),
    .Y(_2819_));
 sky130_fd_sc_hd__a21oi_1 _6479_ (.A1(_2817_),
    .A2(_2818_),
    .B1(_2819_),
    .Y(_2820_));
 sky130_fd_sc_hd__nand3_1 _6480_ (.A(_2817_),
    .B(_2819_),
    .C(_2818_),
    .Y(_2821_));
 sky130_fd_sc_hd__nand2_1 _6481_ (.A(_2821_),
    .B(_2647_),
    .Y(_2822_));
 sky130_fd_sc_hd__nor2_1 _6482_ (.A(_2820_),
    .B(_2822_),
    .Y(\egd_top.exp_golomb_decoding.te_range[2] ));
 sky130_fd_sc_hd__or3_1 _6483_ (.A(_2716_),
    .B(_2650_),
    .C(_2693_),
    .X(_2823_));
 sky130_fd_sc_hd__inv_2 _6484_ (.A(_2823_),
    .Y(\egd_top.BitStream_buffer.exp_golomb_len[1] ));
 sky130_fd_sc_hd__or3_1 _6485_ (.A(_2716_),
    .B(_2650_),
    .C(_2685_),
    .X(_2824_));
 sky130_fd_sc_hd__inv_2 _6486_ (.A(_2824_),
    .Y(\egd_top.BitStream_buffer.exp_golomb_len[2] ));
 sky130_fd_sc_hd__or3_1 _6487_ (.A(_2716_),
    .B(_2650_),
    .C(_2667_),
    .X(_2825_));
 sky130_fd_sc_hd__inv_2 _6488_ (.A(_2825_),
    .Y(\egd_top.BitStream_buffer.exp_golomb_len[3] ));
 sky130_fd_sc_hd__nand2_1 _6489_ (.A(_2817_),
    .B(_2818_),
    .Y(net22));
 sky130_fd_sc_hd__nand2_1 _6490_ (.A(_2798_),
    .B(_2764_),
    .Y(_2826_));
 sky130_fd_sc_hd__nand2_1 _6491_ (.A(_2707_),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[5] ),
    .Y(_2827_));
 sky130_fd_sc_hd__o21ai_2 _6492_ (.A1(_1652_),
    .A2(_2707_),
    .B1(_2827_),
    .Y(_2828_));
 sky130_fd_sc_hd__inv_2 _6493_ (.A(_2828_),
    .Y(_2829_));
 sky130_fd_sc_hd__o21ai_1 _6494_ (.A1(_2761_),
    .A2(_2826_),
    .B1(_2829_),
    .Y(_2830_));
 sky130_fd_sc_hd__nor2_1 _6495_ (.A(_2761_),
    .B(_2826_),
    .Y(_2831_));
 sky130_fd_sc_hd__nand2_1 _6496_ (.A(_2831_),
    .B(_2828_),
    .Y(_2832_));
 sky130_fd_sc_hd__nand3_1 _6497_ (.A(_2830_),
    .B(_2832_),
    .C(_2710_),
    .Y(_2833_));
 sky130_fd_sc_hd__nor2_1 _6498_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[9] ),
    .B(_2805_),
    .Y(_2834_));
 sky130_fd_sc_hd__nor2_1 _6499_ (.A(_1406_),
    .B(_2806_),
    .Y(_2835_));
 sky130_fd_sc_hd__nand2_1 _6500_ (.A(_2744_),
    .B(_2734_),
    .Y(_2836_));
 sky130_fd_sc_hd__xor2_1 _6501_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[11] ),
    .B(_2836_),
    .X(_2837_));
 sky130_fd_sc_hd__o32a_1 _6502_ (.A1(_2834_),
    .A2(_2835_),
    .A3(_2689_),
    .B1(_2694_),
    .B2(_2837_),
    .X(_2838_));
 sky130_fd_sc_hd__nand2_1 _6503_ (.A(_2833_),
    .B(_2838_),
    .Y(_2839_));
 sky130_fd_sc_hd__nand2_2 _6504_ (.A(_2839_),
    .B(_2959_),
    .Y(_2840_));
 sky130_fd_sc_hd__nor2_1 _6505_ (.A(_2788_),
    .B(_2811_),
    .Y(_2841_));
 sky130_fd_sc_hd__nor2_1 _6506_ (.A(_2840_),
    .B(_2841_),
    .Y(_2842_));
 sky130_fd_sc_hd__nand2_1 _6507_ (.A(_2840_),
    .B(_2814_),
    .Y(_2843_));
 sky130_fd_sc_hd__nor2_1 _6508_ (.A(_2788_),
    .B(_2843_),
    .Y(_2844_));
 sky130_fd_sc_hd__o21a_1 _6509_ (.A1(_2842_),
    .A2(_2844_),
    .B1(_2713_),
    .X(_2845_));
 sky130_fd_sc_hd__nor2_1 _6510_ (.A(_2755_),
    .B(_2786_),
    .Y(_2846_));
 sky130_fd_sc_hd__nand2_1 _6511_ (.A(_2811_),
    .B(_2846_),
    .Y(_2847_));
 sky130_fd_sc_hd__nor2_1 _6512_ (.A(_2840_),
    .B(_2847_),
    .Y(_2848_));
 sky130_fd_sc_hd__and2_1 _6513_ (.A(_2847_),
    .B(_2840_),
    .X(_2849_));
 sky130_fd_sc_hd__o21ai_1 _6514_ (.A1(_2848_),
    .A2(_2849_),
    .B1(_2714_),
    .Y(_2850_));
 sky130_fd_sc_hd__nand2_1 _6515_ (.A(_2850_),
    .B(_2756_),
    .Y(_2851_));
 sky130_fd_sc_hd__inv_2 _6516_ (.A(_2760_),
    .Y(_2852_));
 sky130_fd_sc_hd__nand2_1 _6517_ (.A(_2813_),
    .B(_2852_),
    .Y(_2853_));
 sky130_fd_sc_hd__o21ai_2 _6518_ (.A1(_2845_),
    .A2(_2851_),
    .B1(_2853_),
    .Y(net23));
 sky130_fd_sc_hd__nand2_1 _6519_ (.A(_2844_),
    .B(_2713_),
    .Y(_2854_));
 sky130_fd_sc_hd__o21ai_1 _6520_ (.A1(_2840_),
    .A2(_2847_),
    .B1(_2714_),
    .Y(_2855_));
 sky130_fd_sc_hd__nand2_1 _6521_ (.A(_2854_),
    .B(_2855_),
    .Y(_2856_));
 sky130_fd_sc_hd__nor2_1 _6522_ (.A(_2768_),
    .B(_2794_),
    .Y(_2857_));
 sky130_fd_sc_hd__nand3_1 _6523_ (.A(_2857_),
    .B(_2792_),
    .C(_2829_),
    .Y(_2858_));
 sky130_fd_sc_hd__a21oi_2 _6524_ (.A1(_2707_),
    .A2(_1774_),
    .B1(_1530_),
    .Y(_2859_));
 sky130_fd_sc_hd__inv_2 _6525_ (.A(_2859_),
    .Y(_2860_));
 sky130_fd_sc_hd__nand2_1 _6526_ (.A(_2858_),
    .B(_2860_),
    .Y(_2861_));
 sky130_fd_sc_hd__nand3_1 _6527_ (.A(_2831_),
    .B(_2859_),
    .C(_2829_),
    .Y(_2862_));
 sky130_fd_sc_hd__nand3_1 _6528_ (.A(_2861_),
    .B(_2862_),
    .C(_2710_),
    .Y(_2863_));
 sky130_fd_sc_hd__nor2_1 _6529_ (.A(_2737_),
    .B(_2806_),
    .Y(_2864_));
 sky130_fd_sc_hd__a211o_1 _6530_ (.A1(_1282_),
    .A2(_2806_),
    .B1(_2864_),
    .C1(_2689_),
    .X(_2865_));
 sky130_fd_sc_hd__nand2_1 _6531_ (.A(_2863_),
    .B(_2865_),
    .Y(_2866_));
 sky130_fd_sc_hd__nand2_1 _6532_ (.A(_2866_),
    .B(_2959_),
    .Y(_2867_));
 sky130_fd_sc_hd__nand2_1 _6533_ (.A(_2856_),
    .B(_2867_),
    .Y(_2868_));
 sky130_fd_sc_hd__inv_2 _6534_ (.A(_2867_),
    .Y(_2869_));
 sky130_fd_sc_hd__nand3_1 _6535_ (.A(_2854_),
    .B(_2855_),
    .C(_2869_),
    .Y(_2870_));
 sky130_fd_sc_hd__nand3_1 _6536_ (.A(_2868_),
    .B(_2870_),
    .C(_2756_),
    .Y(_2871_));
 sky130_fd_sc_hd__nand2_1 _6537_ (.A(_2839_),
    .B(_2852_),
    .Y(_2872_));
 sky130_fd_sc_hd__nand2_1 _6538_ (.A(_2871_),
    .B(_2872_),
    .Y(net24));
 sky130_fd_sc_hd__nand3_1 _6539_ (.A(_2866_),
    .B(_2959_),
    .C(_2839_),
    .Y(_2873_));
 sky130_fd_sc_hd__inv_2 _6540_ (.A(_2873_),
    .Y(_2874_));
 sky130_fd_sc_hd__nor3_1 _6541_ (.A(_2786_),
    .B(_2755_),
    .C(_2814_),
    .Y(_2875_));
 sky130_fd_sc_hd__nand2_1 _6542_ (.A(_2874_),
    .B(_2875_),
    .Y(_2876_));
 sky130_fd_sc_hd__nor2_1 _6543_ (.A(_2859_),
    .B(_2828_),
    .Y(_2877_));
 sky130_fd_sc_hd__nand2_1 _6544_ (.A(_2831_),
    .B(_2877_),
    .Y(_2878_));
 sky130_fd_sc_hd__o21ai_2 _6545_ (.A1(_1652_),
    .A2(_2720_),
    .B1(_1406_),
    .Y(_2879_));
 sky130_fd_sc_hd__inv_2 _6546_ (.A(_2879_),
    .Y(_2880_));
 sky130_fd_sc_hd__nand2_1 _6547_ (.A(_2878_),
    .B(_2880_),
    .Y(_2881_));
 sky130_fd_sc_hd__nand3_1 _6548_ (.A(_2831_),
    .B(_2877_),
    .C(_2879_),
    .Y(_2882_));
 sky130_fd_sc_hd__nand3_1 _6549_ (.A(_2881_),
    .B(_2710_),
    .C(_2882_),
    .Y(_2883_));
 sky130_fd_sc_hd__nor2_2 _6550_ (.A(_2716_),
    .B(_2883_),
    .Y(_2884_));
 sky130_fd_sc_hd__inv_2 _6551_ (.A(_2884_),
    .Y(_2885_));
 sky130_fd_sc_hd__nand2_1 _6552_ (.A(_2876_),
    .B(_2885_),
    .Y(_2886_));
 sky130_fd_sc_hd__nand3_1 _6553_ (.A(_2874_),
    .B(_2875_),
    .C(_2884_),
    .Y(_2887_));
 sky130_fd_sc_hd__nand2_1 _6554_ (.A(_2886_),
    .B(_2887_),
    .Y(_2888_));
 sky130_fd_sc_hd__nand2_1 _6555_ (.A(_2888_),
    .B(_2714_),
    .Y(_2889_));
 sky130_fd_sc_hd__nand3_1 _6556_ (.A(_2841_),
    .B(_2840_),
    .C(_2867_),
    .Y(_2890_));
 sky130_fd_sc_hd__nand2_1 _6557_ (.A(_2890_),
    .B(_2884_),
    .Y(_2891_));
 sky130_fd_sc_hd__a21oi_1 _6558_ (.A1(_2866_),
    .A2(_2959_),
    .B1(_2884_),
    .Y(_2892_));
 sky130_fd_sc_hd__nand2_1 _6559_ (.A(_2844_),
    .B(_2892_),
    .Y(_2893_));
 sky130_fd_sc_hd__nand2_1 _6560_ (.A(_2891_),
    .B(_2893_),
    .Y(_2894_));
 sky130_fd_sc_hd__nand2_1 _6561_ (.A(_2894_),
    .B(_2713_),
    .Y(_2895_));
 sky130_fd_sc_hd__nand3_1 _6562_ (.A(_2889_),
    .B(_2895_),
    .C(_2756_),
    .Y(_2896_));
 sky130_fd_sc_hd__nand2_1 _6563_ (.A(_2866_),
    .B(_2852_),
    .Y(_2897_));
 sky130_fd_sc_hd__nand2_1 _6564_ (.A(_2896_),
    .B(_2897_),
    .Y(net25));
 sky130_fd_sc_hd__nand3_1 _6565_ (.A(_2848_),
    .B(_2884_),
    .C(_2869_),
    .Y(_2898_));
 sky130_fd_sc_hd__or2_1 _6566_ (.A(_2879_),
    .B(_2878_),
    .X(_2899_));
 sky130_fd_sc_hd__nand2_1 _6567_ (.A(_2899_),
    .B(_2707_),
    .Y(_2900_));
 sky130_fd_sc_hd__inv_2 _6568_ (.A(_2900_),
    .Y(_2901_));
 sky130_fd_sc_hd__nand2_1 _6569_ (.A(_2901_),
    .B(_2959_),
    .Y(_2902_));
 sky130_fd_sc_hd__nand2_1 _6570_ (.A(_2898_),
    .B(_2902_),
    .Y(_2903_));
 sky130_fd_sc_hd__nand2_1 _6571_ (.A(_2903_),
    .B(_2714_),
    .Y(_2904_));
 sky130_fd_sc_hd__inv_2 _6572_ (.A(_2902_),
    .Y(_2905_));
 sky130_fd_sc_hd__nand2_1 _6573_ (.A(_2893_),
    .B(_2905_),
    .Y(_2906_));
 sky130_fd_sc_hd__nor2_1 _6574_ (.A(_2717_),
    .B(_2712_),
    .Y(_2907_));
 sky130_fd_sc_hd__nand2_1 _6575_ (.A(_2906_),
    .B(_2907_),
    .Y(_2908_));
 sky130_fd_sc_hd__nand2_1 _6576_ (.A(_2904_),
    .B(_2908_),
    .Y(_2909_));
 sky130_fd_sc_hd__nand2_1 _6577_ (.A(_2909_),
    .B(_2756_),
    .Y(_2910_));
 sky130_fd_sc_hd__a211o_1 _6578_ (.A1(net18),
    .A2(_2650_),
    .B1(_2956_),
    .C1(_2883_),
    .X(_2911_));
 sky130_fd_sc_hd__nand2_1 _6579_ (.A(_2910_),
    .B(_2911_),
    .Y(net26));
 sky130_fd_sc_hd__a211o_1 _6580_ (.A1(net18),
    .A2(_2650_),
    .B1(_2956_),
    .C1(_2900_),
    .X(_2912_));
 sky130_fd_sc_hd__a21bo_1 _6581_ (.A1(_2756_),
    .A2(_2907_),
    .B1_N(_2912_),
    .X(net27));
 sky130_fd_sc_hd__buf_1 _6582_ (.A(wb_clk_i),
    .X(_2913_));
 sky130_fd_sc_hd__buf_1 _6583_ (.A(clknet_1_1__leaf__2913_),
    .X(_2914_));
 sky130_fd_sc_hd__buf_1 _6584_ (.A(clknet_1_1__leaf__2914_),
    .X(_2915_));
 sky130_fd_sc_hd__inv_2 _6585__78 (.A(clknet_1_0__leaf__2915_),
    .Y(net112));
 sky130_fd_sc_hd__inv_2 _6586__79 (.A(clknet_1_0__leaf__2915_),
    .Y(net113));
 sky130_fd_sc_hd__inv_2 _6587__80 (.A(clknet_1_0__leaf__2915_),
    .Y(net114));
 sky130_fd_sc_hd__inv_2 _6588__81 (.A(clknet_1_0__leaf__2915_),
    .Y(net115));
 sky130_fd_sc_hd__inv_2 _6589__82 (.A(clknet_1_0__leaf__2915_),
    .Y(net116));
 sky130_fd_sc_hd__inv_2 _6590__83 (.A(clknet_1_0__leaf__2915_),
    .Y(net117));
 sky130_fd_sc_hd__inv_2 _6591__84 (.A(clknet_1_1__leaf__2915_),
    .Y(net118));
 sky130_fd_sc_hd__inv_2 _6592__85 (.A(clknet_1_1__leaf__2915_),
    .Y(net119));
 sky130_fd_sc_hd__inv_2 _6593__86 (.A(clknet_1_1__leaf__2915_),
    .Y(net120));
 sky130_fd_sc_hd__inv_2 _6594__87 (.A(clknet_1_1__leaf__2915_),
    .Y(net121));
 sky130_fd_sc_hd__inv_2 _6595__88 (.A(clknet_1_0__leaf__2915_),
    .Y(net122));
 sky130_fd_sc_hd__inv_2 _6596__89 (.A(clknet_1_1__leaf__2915_),
    .Y(net123));
 sky130_fd_sc_hd__buf_1 _6597_ (.A(clknet_1_0__leaf__2914_),
    .X(_2916_));
 sky130_fd_sc_hd__inv_2 _6598__90 (.A(clknet_1_1__leaf__2916_),
    .Y(net124));
 sky130_fd_sc_hd__inv_2 _6599__91 (.A(clknet_1_1__leaf__2916_),
    .Y(net125));
 sky130_fd_sc_hd__inv_2 _6600__92 (.A(clknet_1_1__leaf__2916_),
    .Y(net126));
 sky130_fd_sc_hd__inv_2 _6601__93 (.A(clknet_1_1__leaf__2916_),
    .Y(net127));
 sky130_fd_sc_hd__inv_2 _6602__94 (.A(clknet_1_0__leaf__2916_),
    .Y(net128));
 sky130_fd_sc_hd__inv_2 _6603__95 (.A(clknet_1_0__leaf__2916_),
    .Y(net129));
 sky130_fd_sc_hd__inv_2 _6604__96 (.A(clknet_1_0__leaf__2916_),
    .Y(net130));
 sky130_fd_sc_hd__inv_2 _6605__97 (.A(clknet_1_0__leaf__2916_),
    .Y(net131));
 sky130_fd_sc_hd__inv_2 _6606__98 (.A(clknet_1_0__leaf__2916_),
    .Y(net132));
 sky130_fd_sc_hd__inv_2 _6607__99 (.A(clknet_1_0__leaf__2916_),
    .Y(net133));
 sky130_fd_sc_hd__inv_2 _6608__100 (.A(clknet_1_1__leaf__2916_),
    .Y(net134));
 sky130_fd_sc_hd__inv_2 _6609__101 (.A(clknet_1_0__leaf__2916_),
    .Y(net135));
 sky130_fd_sc_hd__buf_1 _6610_ (.A(clknet_1_1__leaf__2914_),
    .X(_2917_));
 sky130_fd_sc_hd__inv_2 _6611__102 (.A(clknet_1_0__leaf__2917_),
    .Y(net136));
 sky130_fd_sc_hd__inv_2 _6612__103 (.A(clknet_1_0__leaf__2917_),
    .Y(net137));
 sky130_fd_sc_hd__inv_2 _6613__104 (.A(clknet_1_0__leaf__2917_),
    .Y(net138));
 sky130_fd_sc_hd__inv_2 _6614__105 (.A(clknet_1_0__leaf__2917_),
    .Y(net139));
 sky130_fd_sc_hd__inv_2 _6615__106 (.A(clknet_1_0__leaf__2917_),
    .Y(net140));
 sky130_fd_sc_hd__inv_2 _6616__107 (.A(clknet_1_1__leaf__2917_),
    .Y(net141));
 sky130_fd_sc_hd__inv_2 _6617__108 (.A(clknet_1_1__leaf__2917_),
    .Y(net142));
 sky130_fd_sc_hd__inv_2 _6618__109 (.A(clknet_1_1__leaf__2917_),
    .Y(net143));
 sky130_fd_sc_hd__inv_2 _6619__110 (.A(clknet_1_1__leaf__2917_),
    .Y(net144));
 sky130_fd_sc_hd__inv_2 _6620__111 (.A(clknet_1_1__leaf__2917_),
    .Y(net145));
 sky130_fd_sc_hd__inv_2 _6621__112 (.A(clknet_1_1__leaf__2917_),
    .Y(net146));
 sky130_fd_sc_hd__inv_2 _6622__113 (.A(clknet_1_1__leaf__2917_),
    .Y(net147));
 sky130_fd_sc_hd__buf_1 _6623_ (.A(clknet_1_1__leaf__2914_),
    .X(_2918_));
 sky130_fd_sc_hd__inv_2 _6624__114 (.A(clknet_1_0__leaf__2918_),
    .Y(net148));
 sky130_fd_sc_hd__inv_2 _6625__115 (.A(clknet_1_0__leaf__2918_),
    .Y(net149));
 sky130_fd_sc_hd__inv_2 _6626__116 (.A(clknet_1_0__leaf__2918_),
    .Y(net150));
 sky130_fd_sc_hd__inv_2 _6627__117 (.A(clknet_1_1__leaf__2918_),
    .Y(net151));
 sky130_fd_sc_hd__inv_2 _6628__118 (.A(clknet_1_0__leaf__2918_),
    .Y(net152));
 sky130_fd_sc_hd__inv_2 _6629__119 (.A(clknet_1_0__leaf__2918_),
    .Y(net153));
 sky130_fd_sc_hd__inv_2 _6630__120 (.A(clknet_1_1__leaf__2918_),
    .Y(net154));
 sky130_fd_sc_hd__inv_2 _6631__121 (.A(clknet_1_1__leaf__2918_),
    .Y(net155));
 sky130_fd_sc_hd__inv_2 _6632__122 (.A(clknet_1_1__leaf__2918_),
    .Y(net156));
 sky130_fd_sc_hd__inv_2 _6633__123 (.A(clknet_1_1__leaf__2918_),
    .Y(net157));
 sky130_fd_sc_hd__inv_2 _6634__124 (.A(clknet_1_1__leaf__2918_),
    .Y(net158));
 sky130_fd_sc_hd__inv_2 _6635__125 (.A(clknet_1_1__leaf__2918_),
    .Y(net159));
 sky130_fd_sc_hd__buf_1 _6636_ (.A(clknet_1_1__leaf__2914_),
    .X(_2919_));
 sky130_fd_sc_hd__inv_2 _6637__126 (.A(clknet_1_0__leaf__2919_),
    .Y(net160));
 sky130_fd_sc_hd__inv_2 _6638__127 (.A(clknet_1_0__leaf__2919_),
    .Y(net161));
 sky130_fd_sc_hd__inv_2 _6639__128 (.A(clknet_1_0__leaf__2919_),
    .Y(net162));
 sky130_fd_sc_hd__inv_2 _6640__129 (.A(clknet_1_0__leaf__2919_),
    .Y(net163));
 sky130_fd_sc_hd__inv_2 _6641__130 (.A(clknet_1_0__leaf__2919_),
    .Y(net164));
 sky130_fd_sc_hd__inv_2 _6642__131 (.A(clknet_1_0__leaf__2919_),
    .Y(net165));
 sky130_fd_sc_hd__inv_2 _6643__132 (.A(clknet_1_1__leaf__2919_),
    .Y(net166));
 sky130_fd_sc_hd__inv_2 _6644__133 (.A(clknet_1_1__leaf__2919_),
    .Y(net167));
 sky130_fd_sc_hd__inv_2 _6645__134 (.A(clknet_1_1__leaf__2919_),
    .Y(net168));
 sky130_fd_sc_hd__inv_2 _6646__135 (.A(clknet_1_1__leaf__2919_),
    .Y(net169));
 sky130_fd_sc_hd__inv_2 _6647__136 (.A(clknet_1_1__leaf__2919_),
    .Y(net170));
 sky130_fd_sc_hd__inv_2 _6648__137 (.A(clknet_1_1__leaf__2919_),
    .Y(net171));
 sky130_fd_sc_hd__buf_1 _6649_ (.A(clknet_1_1__leaf__2914_),
    .X(_2920_));
 sky130_fd_sc_hd__inv_2 _6650__138 (.A(clknet_1_0__leaf__2920_),
    .Y(net172));
 sky130_fd_sc_hd__inv_2 _6651__139 (.A(clknet_1_0__leaf__2920_),
    .Y(net173));
 sky130_fd_sc_hd__inv_2 _6652__140 (.A(clknet_1_0__leaf__2920_),
    .Y(net174));
 sky130_fd_sc_hd__inv_2 _6653__141 (.A(clknet_1_0__leaf__2920_),
    .Y(net175));
 sky130_fd_sc_hd__inv_2 _6654__142 (.A(clknet_1_0__leaf__2920_),
    .Y(net176));
 sky130_fd_sc_hd__inv_2 _6655__143 (.A(clknet_1_0__leaf__2920_),
    .Y(net177));
 sky130_fd_sc_hd__inv_2 _6656__144 (.A(clknet_1_0__leaf__2920_),
    .Y(net178));
 sky130_fd_sc_hd__inv_2 _6657__145 (.A(clknet_1_1__leaf__2920_),
    .Y(net179));
 sky130_fd_sc_hd__inv_2 _6658__146 (.A(clknet_1_1__leaf__2920_),
    .Y(net180));
 sky130_fd_sc_hd__inv_2 _6659__147 (.A(clknet_1_1__leaf__2920_),
    .Y(net181));
 sky130_fd_sc_hd__inv_2 _6660__148 (.A(clknet_1_1__leaf__2920_),
    .Y(net182));
 sky130_fd_sc_hd__inv_2 _6661__149 (.A(clknet_1_1__leaf__2920_),
    .Y(net183));
 sky130_fd_sc_hd__buf_1 _6662_ (.A(clknet_1_0__leaf__2914_),
    .X(_2921_));
 sky130_fd_sc_hd__inv_2 _6663__150 (.A(clknet_1_1__leaf__2921_),
    .Y(net184));
 sky130_fd_sc_hd__inv_2 _6664__151 (.A(clknet_1_1__leaf__2921_),
    .Y(net185));
 sky130_fd_sc_hd__inv_2 _6665__152 (.A(clknet_1_1__leaf__2921_),
    .Y(net186));
 sky130_fd_sc_hd__inv_2 _6666__153 (.A(clknet_1_1__leaf__2921_),
    .Y(net187));
 sky130_fd_sc_hd__inv_2 _6667__154 (.A(clknet_1_1__leaf__2921_),
    .Y(net188));
 sky130_fd_sc_hd__inv_2 _6668__155 (.A(clknet_1_0__leaf__2921_),
    .Y(net189));
 sky130_fd_sc_hd__inv_2 _6669__156 (.A(clknet_1_0__leaf__2921_),
    .Y(net190));
 sky130_fd_sc_hd__inv_2 _6670__157 (.A(clknet_1_0__leaf__2921_),
    .Y(net191));
 sky130_fd_sc_hd__inv_2 _6671__158 (.A(clknet_1_0__leaf__2921_),
    .Y(net192));
 sky130_fd_sc_hd__inv_2 _6672__159 (.A(clknet_1_0__leaf__2921_),
    .Y(net193));
 sky130_fd_sc_hd__inv_2 _6673__160 (.A(clknet_1_0__leaf__2921_),
    .Y(net194));
 sky130_fd_sc_hd__inv_2 _6674__161 (.A(clknet_1_0__leaf__2921_),
    .Y(net195));
 sky130_fd_sc_hd__buf_1 _6675_ (.A(clknet_1_1__leaf__2913_),
    .X(_2922_));
 sky130_fd_sc_hd__inv_2 _6676__6 (.A(clknet_1_1__leaf__2922_),
    .Y(net40));
 sky130_fd_sc_hd__inv_2 _6677__7 (.A(clknet_1_1__leaf__2922_),
    .Y(net41));
 sky130_fd_sc_hd__inv_2 _6678__8 (.A(clknet_1_1__leaf__2922_),
    .Y(net42));
 sky130_fd_sc_hd__inv_2 _6679__9 (.A(clknet_1_1__leaf__2922_),
    .Y(net43));
 sky130_fd_sc_hd__inv_2 _6680__10 (.A(clknet_1_1__leaf__2922_),
    .Y(net44));
 sky130_fd_sc_hd__inv_2 _6681__11 (.A(clknet_1_0__leaf__2922_),
    .Y(net45));
 sky130_fd_sc_hd__inv_2 _6682__12 (.A(clknet_1_0__leaf__2922_),
    .Y(net46));
 sky130_fd_sc_hd__inv_2 _6683__13 (.A(clknet_1_0__leaf__2922_),
    .Y(net47));
 sky130_fd_sc_hd__inv_2 _6684__14 (.A(clknet_1_0__leaf__2922_),
    .Y(net48));
 sky130_fd_sc_hd__inv_2 _6685__15 (.A(clknet_1_0__leaf__2922_),
    .Y(net49));
 sky130_fd_sc_hd__inv_2 _6686__16 (.A(clknet_1_0__leaf__2922_),
    .Y(net50));
 sky130_fd_sc_hd__inv_2 _6687__17 (.A(clknet_1_0__leaf__2922_),
    .Y(net51));
 sky130_fd_sc_hd__buf_1 _6688_ (.A(clknet_1_1__leaf__2913_),
    .X(_2923_));
 sky130_fd_sc_hd__inv_2 _6689__18 (.A(clknet_1_1__leaf__2923_),
    .Y(net52));
 sky130_fd_sc_hd__inv_2 _6690__19 (.A(clknet_1_1__leaf__2923_),
    .Y(net53));
 sky130_fd_sc_hd__inv_2 _6691__20 (.A(clknet_1_1__leaf__2923_),
    .Y(net54));
 sky130_fd_sc_hd__inv_2 _6692__21 (.A(clknet_1_1__leaf__2923_),
    .Y(net55));
 sky130_fd_sc_hd__inv_2 _6693__22 (.A(clknet_1_1__leaf__2923_),
    .Y(net56));
 sky130_fd_sc_hd__inv_2 _6694__23 (.A(clknet_1_0__leaf__2923_),
    .Y(net57));
 sky130_fd_sc_hd__inv_2 _6695__24 (.A(clknet_1_1__leaf__2923_),
    .Y(net58));
 sky130_fd_sc_hd__inv_2 _6696__25 (.A(clknet_1_0__leaf__2923_),
    .Y(net59));
 sky130_fd_sc_hd__inv_2 _6697__26 (.A(clknet_1_0__leaf__2923_),
    .Y(net60));
 sky130_fd_sc_hd__inv_2 _6698__27 (.A(clknet_1_0__leaf__2923_),
    .Y(net61));
 sky130_fd_sc_hd__inv_2 _6699__28 (.A(clknet_1_0__leaf__2923_),
    .Y(net62));
 sky130_fd_sc_hd__inv_2 _6700__29 (.A(clknet_1_0__leaf__2923_),
    .Y(net63));
 sky130_fd_sc_hd__buf_1 _6701_ (.A(clknet_1_0__leaf__2913_),
    .X(_2924_));
 sky130_fd_sc_hd__inv_2 _6702__30 (.A(clknet_1_1__leaf__2924_),
    .Y(net64));
 sky130_fd_sc_hd__inv_2 _6703__31 (.A(clknet_1_1__leaf__2924_),
    .Y(net65));
 sky130_fd_sc_hd__inv_2 _6704__32 (.A(clknet_1_1__leaf__2924_),
    .Y(net66));
 sky130_fd_sc_hd__inv_2 _6705__33 (.A(clknet_1_1__leaf__2924_),
    .Y(net67));
 sky130_fd_sc_hd__inv_2 _6706__34 (.A(clknet_1_0__leaf__2924_),
    .Y(net68));
 sky130_fd_sc_hd__inv_2 _6707__35 (.A(clknet_1_0__leaf__2924_),
    .Y(net69));
 sky130_fd_sc_hd__inv_2 _6708__36 (.A(clknet_1_0__leaf__2924_),
    .Y(net70));
 sky130_fd_sc_hd__inv_2 _6709__37 (.A(clknet_1_0__leaf__2924_),
    .Y(net71));
 sky130_fd_sc_hd__inv_2 _6710__38 (.A(clknet_1_0__leaf__2924_),
    .Y(net72));
 sky130_fd_sc_hd__inv_2 _6711__39 (.A(clknet_1_0__leaf__2924_),
    .Y(net73));
 sky130_fd_sc_hd__inv_2 _6712__40 (.A(clknet_1_0__leaf__2924_),
    .Y(net74));
 sky130_fd_sc_hd__inv_2 _6713__41 (.A(clknet_1_1__leaf__2924_),
    .Y(net75));
 sky130_fd_sc_hd__buf_1 _6714_ (.A(clknet_1_0__leaf__2913_),
    .X(_2925_));
 sky130_fd_sc_hd__inv_2 _6715__42 (.A(clknet_1_1__leaf__2925_),
    .Y(net76));
 sky130_fd_sc_hd__inv_2 _6716__43 (.A(clknet_1_1__leaf__2925_),
    .Y(net77));
 sky130_fd_sc_hd__inv_2 _6717__44 (.A(clknet_1_0__leaf__2925_),
    .Y(net78));
 sky130_fd_sc_hd__inv_2 _6718__45 (.A(clknet_1_0__leaf__2925_),
    .Y(net79));
 sky130_fd_sc_hd__inv_2 _6719__46 (.A(clknet_1_0__leaf__2925_),
    .Y(net80));
 sky130_fd_sc_hd__inv_2 _6720__47 (.A(clknet_1_1__leaf__2925_),
    .Y(net81));
 sky130_fd_sc_hd__inv_2 _6721__48 (.A(clknet_1_0__leaf__2925_),
    .Y(net82));
 sky130_fd_sc_hd__inv_2 _6722__49 (.A(clknet_1_0__leaf__2925_),
    .Y(net83));
 sky130_fd_sc_hd__inv_2 _6723__50 (.A(clknet_1_1__leaf__2925_),
    .Y(net84));
 sky130_fd_sc_hd__inv_2 _6724__51 (.A(clknet_1_1__leaf__2925_),
    .Y(net85));
 sky130_fd_sc_hd__inv_2 _6725__52 (.A(clknet_1_1__leaf__2925_),
    .Y(net86));
 sky130_fd_sc_hd__inv_2 _6726__53 (.A(clknet_1_1__leaf__2925_),
    .Y(net87));
 sky130_fd_sc_hd__buf_1 _6727_ (.A(clknet_1_0__leaf__2913_),
    .X(_2926_));
 sky130_fd_sc_hd__inv_2 _6728__54 (.A(clknet_1_1__leaf__2926_),
    .Y(net88));
 sky130_fd_sc_hd__inv_2 _6729__55 (.A(clknet_1_1__leaf__2926_),
    .Y(net89));
 sky130_fd_sc_hd__inv_2 _6730__56 (.A(clknet_1_1__leaf__2926_),
    .Y(net90));
 sky130_fd_sc_hd__inv_2 _6731__57 (.A(clknet_1_1__leaf__2926_),
    .Y(net91));
 sky130_fd_sc_hd__inv_2 _6732__58 (.A(clknet_1_1__leaf__2926_),
    .Y(net92));
 sky130_fd_sc_hd__inv_2 _6733__59 (.A(clknet_1_1__leaf__2926_),
    .Y(net93));
 sky130_fd_sc_hd__inv_2 _6734__60 (.A(clknet_1_1__leaf__2926_),
    .Y(net94));
 sky130_fd_sc_hd__inv_2 _6735__61 (.A(clknet_1_0__leaf__2926_),
    .Y(net95));
 sky130_fd_sc_hd__inv_2 _6736__62 (.A(clknet_1_0__leaf__2926_),
    .Y(net96));
 sky130_fd_sc_hd__inv_2 _6737__63 (.A(clknet_1_0__leaf__2926_),
    .Y(net97));
 sky130_fd_sc_hd__inv_2 _6738__64 (.A(clknet_1_0__leaf__2926_),
    .Y(net98));
 sky130_fd_sc_hd__inv_2 _6739__65 (.A(clknet_1_0__leaf__2926_),
    .Y(net99));
 sky130_fd_sc_hd__buf_1 _6740_ (.A(clknet_1_0__leaf__2913_),
    .X(_2927_));
 sky130_fd_sc_hd__inv_2 _6741__66 (.A(clknet_1_1__leaf__2927_),
    .Y(net100));
 sky130_fd_sc_hd__inv_2 _6742__67 (.A(clknet_1_1__leaf__2927_),
    .Y(net101));
 sky130_fd_sc_hd__inv_2 _6743__68 (.A(clknet_1_0__leaf__2927_),
    .Y(net102));
 sky130_fd_sc_hd__inv_2 _6744__69 (.A(clknet_1_0__leaf__2927_),
    .Y(net103));
 sky130_fd_sc_hd__inv_2 _6745__70 (.A(clknet_1_0__leaf__2927_),
    .Y(net104));
 sky130_fd_sc_hd__inv_2 _6746__71 (.A(clknet_1_0__leaf__2927_),
    .Y(net105));
 sky130_fd_sc_hd__inv_2 _6747__72 (.A(clknet_1_0__leaf__2927_),
    .Y(net106));
 sky130_fd_sc_hd__inv_2 _6748__73 (.A(clknet_1_0__leaf__2927_),
    .Y(net107));
 sky130_fd_sc_hd__inv_2 _6749__74 (.A(clknet_1_0__leaf__2927_),
    .Y(net108));
 sky130_fd_sc_hd__inv_2 _6750__75 (.A(clknet_1_1__leaf__2927_),
    .Y(net109));
 sky130_fd_sc_hd__inv_2 _6751__76 (.A(clknet_1_1__leaf__2927_),
    .Y(net110));
 sky130_fd_sc_hd__inv_2 _6752__77 (.A(clknet_1_1__leaf__2927_),
    .Y(net111));
 sky130_fd_sc_hd__inv_2 _6753__1 (.A(clknet_1_0__leaf__2914_),
    .Y(net35));
 sky130_fd_sc_hd__inv_2 _6754__2 (.A(clknet_1_0__leaf__2914_),
    .Y(net36));
 sky130_fd_sc_hd__inv_2 _6755__3 (.A(clknet_1_0__leaf__2914_),
    .Y(net37));
 sky130_fd_sc_hd__inv_2 _6756__4 (.A(clknet_1_0__leaf__2914_),
    .Y(net38));
 sky130_fd_sc_hd__inv_2 _6757__5 (.A(clknet_1_0__leaf__2914_),
    .Y(net39));
 sky130_fd_sc_hd__dfxtp_1 _6758_ (.CLK(net112),
    .D(_0161_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[95] ));
 sky130_fd_sc_hd__dfxtp_1 _6759_ (.CLK(net113),
    .D(_0162_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[94] ));
 sky130_fd_sc_hd__dfxtp_1 _6760_ (.CLK(net114),
    .D(_0163_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[93] ));
 sky130_fd_sc_hd__dfxtp_1 _6761_ (.CLK(net115),
    .D(_0164_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[92] ));
 sky130_fd_sc_hd__dfxtp_1 _6762_ (.CLK(net116),
    .D(_0165_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[91] ));
 sky130_fd_sc_hd__dfxtp_1 _6763_ (.CLK(net117),
    .D(_0166_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[90] ));
 sky130_fd_sc_hd__dfxtp_1 _6764_ (.CLK(net118),
    .D(_0167_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[89] ));
 sky130_fd_sc_hd__dfxtp_1 _6765_ (.CLK(net119),
    .D(_0168_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[88] ));
 sky130_fd_sc_hd__dfxtp_1 _6766_ (.CLK(net120),
    .D(_0169_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[87] ));
 sky130_fd_sc_hd__dfxtp_1 _6767_ (.CLK(net121),
    .D(_0170_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[86] ));
 sky130_fd_sc_hd__dfxtp_1 _6768_ (.CLK(net122),
    .D(_0171_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[85] ));
 sky130_fd_sc_hd__dfxtp_1 _6769_ (.CLK(net123),
    .D(_0172_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[84] ));
 sky130_fd_sc_hd__dfxtp_1 _6770_ (.CLK(net124),
    .D(_0173_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[83] ));
 sky130_fd_sc_hd__dfxtp_1 _6771_ (.CLK(net125),
    .D(_0174_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[82] ));
 sky130_fd_sc_hd__dfxtp_1 _6772_ (.CLK(net126),
    .D(_0175_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[81] ));
 sky130_fd_sc_hd__dfxtp_1 _6773_ (.CLK(net127),
    .D(_0176_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[80] ));
 sky130_fd_sc_hd__dfxtp_1 _6774_ (.CLK(net128),
    .D(_0177_),
    .Q(\egd_top.BitStream_buffer.pc_previous[0] ));
 sky130_fd_sc_hd__dfxtp_1 _6775_ (.CLK(net129),
    .D(_0178_),
    .Q(\egd_top.BitStream_buffer.pc_previous[1] ));
 sky130_fd_sc_hd__dfxtp_1 _6776_ (.CLK(net130),
    .D(_0179_),
    .Q(\egd_top.BitStream_buffer.pc_previous[2] ));
 sky130_fd_sc_hd__dfxtp_1 _6777_ (.CLK(net131),
    .D(_0180_),
    .Q(\egd_top.BitStream_buffer.pc_previous[3] ));
 sky130_fd_sc_hd__dfxtp_2 _6778_ (.CLK(net132),
    .D(_0181_),
    .Q(\egd_top.BitStream_buffer.pc_previous[4] ));
 sky130_fd_sc_hd__dfxtp_1 _6779_ (.CLK(net133),
    .D(_0182_),
    .Q(\egd_top.BitStream_buffer.pc_previous[5] ));
 sky130_fd_sc_hd__dfxtp_2 _6780_ (.CLK(net134),
    .D(_0183_),
    .Q(\egd_top.BitStream_buffer.pc_previous[6] ));
 sky130_fd_sc_hd__dfxtp_1 _6781_ (.CLK(net135),
    .D(_0184_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[111] ));
 sky130_fd_sc_hd__dfxtp_1 _6782_ (.CLK(net136),
    .D(_0185_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[110] ));
 sky130_fd_sc_hd__dfxtp_1 _6783_ (.CLK(net137),
    .D(_0186_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[109] ));
 sky130_fd_sc_hd__dfxtp_1 _6784_ (.CLK(net138),
    .D(_0187_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[108] ));
 sky130_fd_sc_hd__dfxtp_1 _6785_ (.CLK(net139),
    .D(_0188_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[107] ));
 sky130_fd_sc_hd__dfxtp_1 _6786_ (.CLK(net140),
    .D(_0189_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[106] ));
 sky130_fd_sc_hd__dfxtp_1 _6787_ (.CLK(net141),
    .D(_0190_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[105] ));
 sky130_fd_sc_hd__dfxtp_1 _6788_ (.CLK(net142),
    .D(_0191_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[104] ));
 sky130_fd_sc_hd__dfxtp_1 _6789_ (.CLK(net143),
    .D(_0192_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[103] ));
 sky130_fd_sc_hd__dfxtp_1 _6790_ (.CLK(net144),
    .D(_0193_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[102] ));
 sky130_fd_sc_hd__dfxtp_1 _6791_ (.CLK(net145),
    .D(_0194_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[101] ));
 sky130_fd_sc_hd__dfxtp_1 _6792_ (.CLK(net146),
    .D(_0195_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[100] ));
 sky130_fd_sc_hd__dfxtp_1 _6793_ (.CLK(net147),
    .D(_0196_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[99] ));
 sky130_fd_sc_hd__dfxtp_1 _6794_ (.CLK(net148),
    .D(_0197_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[98] ));
 sky130_fd_sc_hd__dfxtp_1 _6795_ (.CLK(net149),
    .D(_0198_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[97] ));
 sky130_fd_sc_hd__dfxtp_1 _6796_ (.CLK(net150),
    .D(_0199_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[96] ));
 sky130_fd_sc_hd__dfxtp_1 _6797_ (.CLK(net151),
    .D(_0200_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[79] ));
 sky130_fd_sc_hd__dfxtp_1 _6798_ (.CLK(net152),
    .D(_0201_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[78] ));
 sky130_fd_sc_hd__dfxtp_1 _6799_ (.CLK(net153),
    .D(_0202_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[77] ));
 sky130_fd_sc_hd__dfxtp_1 _6800_ (.CLK(net154),
    .D(_0203_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[76] ));
 sky130_fd_sc_hd__dfxtp_1 _6801_ (.CLK(net155),
    .D(_0204_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[75] ));
 sky130_fd_sc_hd__dfxtp_1 _6802_ (.CLK(net156),
    .D(_0205_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[74] ));
 sky130_fd_sc_hd__dfxtp_1 _6803_ (.CLK(net157),
    .D(_0206_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[73] ));
 sky130_fd_sc_hd__dfxtp_1 _6804_ (.CLK(net158),
    .D(_0207_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[72] ));
 sky130_fd_sc_hd__dfxtp_1 _6805_ (.CLK(net159),
    .D(_0208_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[71] ));
 sky130_fd_sc_hd__dfxtp_1 _6806_ (.CLK(net160),
    .D(_0209_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[70] ));
 sky130_fd_sc_hd__dfxtp_1 _6807_ (.CLK(net161),
    .D(_0210_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[69] ));
 sky130_fd_sc_hd__dfxtp_1 _6808_ (.CLK(net162),
    .D(_0211_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[68] ));
 sky130_fd_sc_hd__dfxtp_1 _6809_ (.CLK(net163),
    .D(_0212_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[67] ));
 sky130_fd_sc_hd__dfxtp_1 _6810_ (.CLK(net164),
    .D(_0213_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[66] ));
 sky130_fd_sc_hd__dfxtp_1 _6811_ (.CLK(net165),
    .D(_0214_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[65] ));
 sky130_fd_sc_hd__dfxtp_1 _6812_ (.CLK(net166),
    .D(_0215_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[64] ));
 sky130_fd_sc_hd__dfxtp_1 _6813_ (.CLK(net167),
    .D(_0216_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[63] ));
 sky130_fd_sc_hd__dfxtp_1 _6814_ (.CLK(net168),
    .D(_0217_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[62] ));
 sky130_fd_sc_hd__dfxtp_1 _6815_ (.CLK(net169),
    .D(_0218_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[61] ));
 sky130_fd_sc_hd__dfxtp_1 _6816_ (.CLK(net170),
    .D(_0219_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[60] ));
 sky130_fd_sc_hd__dfxtp_1 _6817_ (.CLK(net171),
    .D(_0220_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[59] ));
 sky130_fd_sc_hd__dfxtp_1 _6818_ (.CLK(net172),
    .D(_0221_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[58] ));
 sky130_fd_sc_hd__dfxtp_1 _6819_ (.CLK(net173),
    .D(_0222_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[57] ));
 sky130_fd_sc_hd__dfxtp_1 _6820_ (.CLK(net174),
    .D(_0223_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[56] ));
 sky130_fd_sc_hd__dfxtp_1 _6821_ (.CLK(net175),
    .D(_0224_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[55] ));
 sky130_fd_sc_hd__dfxtp_1 _6822_ (.CLK(net176),
    .D(_0225_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[54] ));
 sky130_fd_sc_hd__dfxtp_1 _6823_ (.CLK(net177),
    .D(_0226_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[53] ));
 sky130_fd_sc_hd__dfxtp_1 _6824_ (.CLK(net178),
    .D(_0227_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[52] ));
 sky130_fd_sc_hd__dfxtp_1 _6825_ (.CLK(net179),
    .D(_0228_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[51] ));
 sky130_fd_sc_hd__dfxtp_1 _6826_ (.CLK(net180),
    .D(_0229_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[50] ));
 sky130_fd_sc_hd__dfxtp_1 _6827_ (.CLK(net181),
    .D(_0230_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[49] ));
 sky130_fd_sc_hd__dfxtp_1 _6828_ (.CLK(net182),
    .D(_0231_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[48] ));
 sky130_fd_sc_hd__dfxtp_1 _6829_ (.CLK(net183),
    .D(_0232_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[47] ));
 sky130_fd_sc_hd__dfxtp_1 _6830_ (.CLK(net184),
    .D(_0233_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[46] ));
 sky130_fd_sc_hd__dfxtp_1 _6831_ (.CLK(net185),
    .D(_0234_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[45] ));
 sky130_fd_sc_hd__dfxtp_1 _6832_ (.CLK(net186),
    .D(_0235_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[44] ));
 sky130_fd_sc_hd__dfxtp_1 _6833_ (.CLK(net187),
    .D(_0236_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[43] ));
 sky130_fd_sc_hd__dfxtp_1 _6834_ (.CLK(net188),
    .D(_0237_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[42] ));
 sky130_fd_sc_hd__dfxtp_1 _6835_ (.CLK(net189),
    .D(_0238_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[41] ));
 sky130_fd_sc_hd__dfxtp_1 _6836_ (.CLK(net190),
    .D(_0239_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[40] ));
 sky130_fd_sc_hd__dfxtp_1 _6837_ (.CLK(net191),
    .D(_0240_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[39] ));
 sky130_fd_sc_hd__dfxtp_1 _6838_ (.CLK(net192),
    .D(_0241_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[38] ));
 sky130_fd_sc_hd__dfxtp_1 _6839_ (.CLK(net193),
    .D(_0242_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[37] ));
 sky130_fd_sc_hd__dfxtp_1 _6840_ (.CLK(net194),
    .D(_0243_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[36] ));
 sky130_fd_sc_hd__dfxtp_1 _6841_ (.CLK(net195),
    .D(_0244_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[35] ));
 sky130_fd_sc_hd__dfxtp_1 _6842_ (.CLK(net40),
    .D(_0245_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[34] ));
 sky130_fd_sc_hd__dfxtp_1 _6843_ (.CLK(net41),
    .D(_0246_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[33] ));
 sky130_fd_sc_hd__dfxtp_1 _6844_ (.CLK(net42),
    .D(_0247_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[32] ));
 sky130_fd_sc_hd__dfxtp_1 _6845_ (.CLK(net43),
    .D(_0248_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[31] ));
 sky130_fd_sc_hd__dfxtp_1 _6846_ (.CLK(net44),
    .D(_0249_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[30] ));
 sky130_fd_sc_hd__dfxtp_1 _6847_ (.CLK(net45),
    .D(_0250_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[29] ));
 sky130_fd_sc_hd__dfxtp_1 _6848_ (.CLK(net46),
    .D(_0251_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[28] ));
 sky130_fd_sc_hd__dfxtp_1 _6849_ (.CLK(net47),
    .D(_0252_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[27] ));
 sky130_fd_sc_hd__dfxtp_1 _6850_ (.CLK(net48),
    .D(_0253_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[26] ));
 sky130_fd_sc_hd__dfxtp_1 _6851_ (.CLK(net49),
    .D(_0254_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[25] ));
 sky130_fd_sc_hd__dfxtp_1 _6852_ (.CLK(net50),
    .D(_0255_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[24] ));
 sky130_fd_sc_hd__dfxtp_1 _6853_ (.CLK(net51),
    .D(_0256_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[23] ));
 sky130_fd_sc_hd__dfxtp_1 _6854_ (.CLK(net52),
    .D(_0257_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[22] ));
 sky130_fd_sc_hd__dfxtp_1 _6855_ (.CLK(net53),
    .D(_0258_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[21] ));
 sky130_fd_sc_hd__dfxtp_1 _6856_ (.CLK(net54),
    .D(_0259_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[20] ));
 sky130_fd_sc_hd__dfxtp_1 _6857_ (.CLK(net55),
    .D(_0260_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[19] ));
 sky130_fd_sc_hd__dfxtp_1 _6858_ (.CLK(net56),
    .D(_0261_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[18] ));
 sky130_fd_sc_hd__dfxtp_1 _6859_ (.CLK(net57),
    .D(_0262_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[17] ));
 sky130_fd_sc_hd__dfxtp_2 _6860_ (.CLK(net58),
    .D(_0263_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[16] ));
 sky130_fd_sc_hd__dfxtp_2 _6861_ (.CLK(net59),
    .D(_0264_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[15] ));
 sky130_fd_sc_hd__dfxtp_2 _6862_ (.CLK(net60),
    .D(_0265_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[14] ));
 sky130_fd_sc_hd__dfxtp_2 _6863_ (.CLK(net61),
    .D(_0266_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[13] ));
 sky130_fd_sc_hd__dfxtp_4 _6864_ (.CLK(net62),
    .D(_0267_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[12] ));
 sky130_fd_sc_hd__dfxtp_2 _6865_ (.CLK(net63),
    .D(_0268_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[11] ));
 sky130_fd_sc_hd__dfxtp_4 _6866_ (.CLK(net64),
    .D(_0269_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[10] ));
 sky130_fd_sc_hd__dfxtp_2 _6867_ (.CLK(net65),
    .D(_0270_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[9] ));
 sky130_fd_sc_hd__dfxtp_2 _6868_ (.CLK(net66),
    .D(_0271_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[8] ));
 sky130_fd_sc_hd__dfxtp_2 _6869_ (.CLK(net67),
    .D(_0272_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[7] ));
 sky130_fd_sc_hd__dfxtp_1 _6870_ (.CLK(net68),
    .D(_0273_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[6] ));
 sky130_fd_sc_hd__dfxtp_1 _6871_ (.CLK(net69),
    .D(_0274_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[5] ));
 sky130_fd_sc_hd__dfxtp_1 _6872_ (.CLK(net70),
    .D(_0275_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[4] ));
 sky130_fd_sc_hd__dfxtp_1 _6873_ (.CLK(net71),
    .D(_0276_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[3] ));
 sky130_fd_sc_hd__dfxtp_1 _6874_ (.CLK(net72),
    .D(_0277_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[2] ));
 sky130_fd_sc_hd__dfxtp_1 _6875_ (.CLK(net73),
    .D(_0278_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[1] ));
 sky130_fd_sc_hd__dfxtp_1 _6876_ (.CLK(net74),
    .D(_0279_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _6877_ (.CLK(net75),
    .D(_0280_),
    .Q(\egd_top.BitStream_buffer.buffer_index[4] ));
 sky130_fd_sc_hd__dfxtp_1 _6878_ (.CLK(net76),
    .D(_0281_),
    .Q(\egd_top.BitStream_buffer.buffer_index[5] ));
 sky130_fd_sc_hd__dfxtp_1 _6879_ (.CLK(net77),
    .D(_0282_),
    .Q(\egd_top.BitStream_buffer.buffer_index[6] ));
 sky130_fd_sc_hd__dfxtp_1 _6880_ (.CLK(net78),
    .D(_0283_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[1] ));
 sky130_fd_sc_hd__dfxtp_1 _6881_ (.CLK(net79),
    .D(_0284_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[2] ));
 sky130_fd_sc_hd__dfxtp_1 _6882_ (.CLK(net80),
    .D(_0285_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[3] ));
 sky130_fd_sc_hd__dfxtp_1 _6883_ (.CLK(net81),
    .D(_0286_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[4] ));
 sky130_fd_sc_hd__dfxtp_2 _6884_ (.CLK(net82),
    .D(_0287_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[5] ));
 sky130_fd_sc_hd__dfxtp_1 _6885_ (.CLK(net83),
    .D(_0288_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[6] ));
 sky130_fd_sc_hd__dfxtp_1 _6886_ (.CLK(net84),
    .D(_0289_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[7] ));
 sky130_fd_sc_hd__dfxtp_1 _6887_ (.CLK(net85),
    .D(_0290_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[8] ));
 sky130_fd_sc_hd__dfxtp_1 _6888_ (.CLK(net86),
    .D(_0291_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[9] ));
 sky130_fd_sc_hd__dfxtp_1 _6889_ (.CLK(net87),
    .D(_0292_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[10] ));
 sky130_fd_sc_hd__dfxtp_2 _6890_ (.CLK(net88),
    .D(_0293_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[11] ));
 sky130_fd_sc_hd__dfxtp_1 _6891_ (.CLK(net89),
    .D(_0294_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[12] ));
 sky130_fd_sc_hd__dfxtp_2 _6892_ (.CLK(net90),
    .D(_0295_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[13] ));
 sky130_fd_sc_hd__dfxtp_1 _6893_ (.CLK(net91),
    .D(_0296_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[14] ));
 sky130_fd_sc_hd__dfxtp_1 _6894_ (.CLK(net92),
    .D(_0297_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[15] ));
 sky130_fd_sc_hd__dfxtp_1 _6895_ (.CLK(net93),
    .D(_0298_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[127] ));
 sky130_fd_sc_hd__dfxtp_1 _6896_ (.CLK(net94),
    .D(_0299_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[126] ));
 sky130_fd_sc_hd__dfxtp_1 _6897_ (.CLK(net95),
    .D(_0300_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[125] ));
 sky130_fd_sc_hd__dfxtp_1 _6898_ (.CLK(net96),
    .D(_0301_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[124] ));
 sky130_fd_sc_hd__dfxtp_1 _6899_ (.CLK(net97),
    .D(_0302_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[123] ));
 sky130_fd_sc_hd__dfxtp_1 _6900_ (.CLK(net98),
    .D(_0303_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[122] ));
 sky130_fd_sc_hd__dfxtp_1 _6901_ (.CLK(net99),
    .D(_0304_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[121] ));
 sky130_fd_sc_hd__dfxtp_1 _6902_ (.CLK(net100),
    .D(_0305_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[120] ));
 sky130_fd_sc_hd__dfxtp_1 _6903_ (.CLK(net101),
    .D(_0306_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[119] ));
 sky130_fd_sc_hd__dfxtp_1 _6904_ (.CLK(net102),
    .D(_0307_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[118] ));
 sky130_fd_sc_hd__dfxtp_1 _6905_ (.CLK(net103),
    .D(_0308_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[117] ));
 sky130_fd_sc_hd__dfxtp_1 _6906_ (.CLK(net104),
    .D(_0309_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[116] ));
 sky130_fd_sc_hd__dfxtp_1 _6907_ (.CLK(net105),
    .D(_0310_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[115] ));
 sky130_fd_sc_hd__dfxtp_1 _6908_ (.CLK(net106),
    .D(_0311_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[114] ));
 sky130_fd_sc_hd__dfxtp_1 _6909_ (.CLK(net107),
    .D(_0312_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[113] ));
 sky130_fd_sc_hd__dfxtp_1 _6910_ (.CLK(net108),
    .D(_0313_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[112] ));
 sky130_fd_sc_hd__dfxtp_1 _6911_ (.CLK(net109),
    .D(_0314_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_valid_n ));
 sky130_fd_sc_hd__dfxtp_2 _6912_ (.CLK(net110),
    .D(_0315_),
    .Q(net28));
 sky130_fd_sc_hd__dfxtp_2 _6913_ (.CLK(net111),
    .D(_0316_),
    .Q(net29));
 sky130_fd_sc_hd__dfxtp_2 _6914_ (.CLK(net35),
    .D(_0317_),
    .Q(net30));
 sky130_fd_sc_hd__dfxtp_1 _6915_ (.CLK(net36),
    .D(_0318_),
    .Q(net31));
 sky130_fd_sc_hd__dfxtp_2 _6916_ (.CLK(net37),
    .D(_0319_),
    .Q(net32));
 sky130_fd_sc_hd__dfxtp_2 _6917_ (.CLK(net38),
    .D(_0320_),
    .Q(net33));
 sky130_fd_sc_hd__dfxtp_2 _6918_ (.CLK(net39),
    .D(_0321_),
    .Q(net34));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2913_ (.A(_2913_),
    .X(clknet_0__2913_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2914_ (.A(_2914_),
    .X(clknet_0__2914_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2915_ (.A(_2915_),
    .X(clknet_0__2915_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2916_ (.A(_2916_),
    .X(clknet_0__2916_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2917_ (.A(_2917_),
    .X(clknet_0__2917_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2918_ (.A(_2918_),
    .X(clknet_0__2918_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2919_ (.A(_2919_),
    .X(clknet_0__2919_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2920_ (.A(_2920_),
    .X(clknet_0__2920_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2921_ (.A(_2921_),
    .X(clknet_0__2921_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2922_ (.A(_2922_),
    .X(clknet_0__2922_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2923_ (.A(_2923_),
    .X(clknet_0__2923_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2924_ (.A(_2924_),
    .X(clknet_0__2924_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2925_ (.A(_2925_),
    .X(clknet_0__2925_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2926_ (.A(_2926_),
    .X(clknet_0__2926_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2927_ (.A(_2927_),
    .X(clknet_0__2927_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2913_ (.A(clknet_0__2913_),
    .X(clknet_1_0__leaf__2913_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2914_ (.A(clknet_0__2914_),
    .X(clknet_1_0__leaf__2914_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2915_ (.A(clknet_0__2915_),
    .X(clknet_1_0__leaf__2915_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2916_ (.A(clknet_0__2916_),
    .X(clknet_1_0__leaf__2916_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2917_ (.A(clknet_0__2917_),
    .X(clknet_1_0__leaf__2917_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2918_ (.A(clknet_0__2918_),
    .X(clknet_1_0__leaf__2918_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2919_ (.A(clknet_0__2919_),
    .X(clknet_1_0__leaf__2919_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2920_ (.A(clknet_0__2920_),
    .X(clknet_1_0__leaf__2920_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2921_ (.A(clknet_0__2921_),
    .X(clknet_1_0__leaf__2921_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2922_ (.A(clknet_0__2922_),
    .X(clknet_1_0__leaf__2922_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2923_ (.A(clknet_0__2923_),
    .X(clknet_1_0__leaf__2923_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2924_ (.A(clknet_0__2924_),
    .X(clknet_1_0__leaf__2924_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2925_ (.A(clknet_0__2925_),
    .X(clknet_1_0__leaf__2925_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2926_ (.A(clknet_0__2926_),
    .X(clknet_1_0__leaf__2926_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2927_ (.A(clknet_0__2927_),
    .X(clknet_1_0__leaf__2927_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2913_ (.A(clknet_0__2913_),
    .X(clknet_1_1__leaf__2913_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2914_ (.A(clknet_0__2914_),
    .X(clknet_1_1__leaf__2914_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2915_ (.A(clknet_0__2915_),
    .X(clknet_1_1__leaf__2915_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2916_ (.A(clknet_0__2916_),
    .X(clknet_1_1__leaf__2916_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2917_ (.A(clknet_0__2917_),
    .X(clknet_1_1__leaf__2917_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2918_ (.A(clknet_0__2918_),
    .X(clknet_1_1__leaf__2918_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2919_ (.A(clknet_0__2919_),
    .X(clknet_1_1__leaf__2919_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2920_ (.A(clknet_0__2920_),
    .X(clknet_1_1__leaf__2920_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2921_ (.A(clknet_0__2921_),
    .X(clknet_1_1__leaf__2921_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2922_ (.A(clknet_0__2922_),
    .X(clknet_1_1__leaf__2922_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2923_ (.A(clknet_0__2923_),
    .X(clknet_1_1__leaf__2923_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2924_ (.A(clknet_0__2924_),
    .X(clknet_1_1__leaf__2924_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2925_ (.A(clknet_0__2925_),
    .X(clknet_1_1__leaf__2925_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2926_ (.A(clknet_0__2926_),
    .X(clknet_1_1__leaf__2926_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2927_ (.A(clknet_0__2927_),
    .X(clknet_1_1__leaf__2927_));
 sky130_fd_sc_hd__buf_1 hold1 (.A(net202),
    .X(net196));
 sky130_fd_sc_hd__clkbuf_2 hold2 (.A(_2556_),
    .X(net197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\egd_top.BitStream_buffer.buffer_index[5] ),
    .X(net198));
 sky130_fd_sc_hd__clkbuf_2 hold4 (.A(_2612_),
    .X(net199));
 sky130_fd_sc_hd__buf_1 hold5 (.A(\egd_top.BitStream_buffer.buffer_index[6] ),
    .X(net200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(\egd_top.BitStream_buffer.buffer_index[4] ),
    .X(net201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\egd_top.BitStream_buffer.buffer_index[4] ),
    .X(net202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(_2450_),
    .X(net203));
 sky130_fd_sc_hd__clkbuf_8 input1 (.A(la_data_in_58_43[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_8 input10 (.A(la_data_in_58_43[3]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_8 input11 (.A(la_data_in_58_43[4]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_8 input12 (.A(la_data_in_58_43[5]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_8 input13 (.A(la_data_in_58_43[6]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_8 input14 (.A(la_data_in_58_43[7]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_8 input15 (.A(la_data_in_58_43[8]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_8 input16 (.A(la_data_in_58_43[9]),
    .X(net16));
 sky130_fd_sc_hd__buf_2 input17 (.A(la_data_in_60_59[0]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_4 input18 (.A(la_data_in_60_59[1]),
    .X(net18));
 sky130_fd_sc_hd__buf_1 input19 (.A(la_data_in_65),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_8 input2 (.A(la_data_in_58_43[10]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_8 input3 (.A(la_data_in_58_43[11]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_8 input4 (.A(la_data_in_58_43[12]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_8 input5 (.A(la_data_in_58_43[13]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_8 input6 (.A(la_data_in_58_43[14]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_8 input7 (.A(la_data_in_58_43[15]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_8 input8 (.A(la_data_in_58_43[1]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_8 input9 (.A(la_data_in_58_43[2]),
    .X(net9));
 sky130_fd_sc_hd__buf_12 output20 (.A(net20),
    .X(la_data_out_23_16[0]));
 sky130_fd_sc_hd__buf_12 output21 (.A(net21),
    .X(la_data_out_23_16[1]));
 sky130_fd_sc_hd__buf_12 output22 (.A(net22),
    .X(la_data_out_23_16[2]));
 sky130_fd_sc_hd__buf_12 output23 (.A(net23),
    .X(la_data_out_23_16[3]));
 sky130_fd_sc_hd__buf_12 output24 (.A(net24),
    .X(la_data_out_23_16[4]));
 sky130_fd_sc_hd__buf_12 output25 (.A(net25),
    .X(la_data_out_23_16[5]));
 sky130_fd_sc_hd__buf_12 output26 (.A(net26),
    .X(la_data_out_23_16[6]));
 sky130_fd_sc_hd__buf_12 output27 (.A(net27),
    .X(la_data_out_23_16[7]));
 sky130_fd_sc_hd__buf_12 output28 (.A(net28),
    .X(la_data_out_26_24[0]));
 sky130_fd_sc_hd__buf_12 output29 (.A(net29),
    .X(la_data_out_26_24[1]));
 sky130_fd_sc_hd__buf_12 output30 (.A(net30),
    .X(la_data_out_26_24[2]));
 sky130_fd_sc_hd__buf_12 output31 (.A(net31),
    .X(la_data_out_30_27[0]));
 sky130_fd_sc_hd__buf_12 output32 (.A(net32),
    .X(la_data_out_30_27[1]));
 sky130_fd_sc_hd__buf_12 output33 (.A(net33),
    .X(la_data_out_30_27[2]));
 sky130_fd_sc_hd__buf_12 output34 (.A(net34),
    .X(la_data_out_30_27[3]));
endmodule

