magic
tech sky130A
timestamp 1676037725
<< properties >>
string GDS_END 34244
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sram_1rw1r_32_256_8_sky130.gds
string GDS_START 33920
<< end >>
