magic
tech sky130A
magscale 1 2
timestamp 1676037725
<< nwell >>
rect -38 261 1878 582
<< pwell >>
rect 42 201 1525 203
rect 42 23 1831 201
rect 42 21 339 23
rect 836 21 1028 23
rect 1440 21 1831 23
rect 42 17 63 21
rect 29 -17 63 17
<< scnmos >>
rect 120 47 150 177
rect 204 47 234 177
rect 328 93 358 177
rect 550 49 580 177
rect 660 49 690 177
rect 922 47 952 177
rect 1108 49 1138 177
rect 1260 49 1290 133
rect 1419 49 1449 177
rect 1539 47 1569 167
rect 1639 47 1669 175
rect 1723 47 1753 175
<< scpmoshvt >>
rect 124 297 154 497
rect 208 297 238 497
rect 328 297 358 425
rect 542 325 572 493
rect 648 325 678 493
rect 889 297 919 497
rect 1108 297 1138 465
rect 1260 297 1290 425
rect 1435 329 1465 457
rect 1538 329 1568 497
rect 1639 297 1669 497
rect 1723 297 1753 497
<< ndiff >>
rect 68 93 120 177
rect 68 59 76 93
rect 110 59 120 93
rect 68 47 120 59
rect 150 129 204 177
rect 150 95 160 129
rect 194 95 204 129
rect 150 47 204 95
rect 234 93 328 177
rect 358 169 442 177
rect 358 135 396 169
rect 430 135 442 169
rect 358 93 442 135
rect 496 165 550 177
rect 496 131 506 165
rect 540 131 550 165
rect 234 89 313 93
rect 234 55 260 89
rect 294 55 313 89
rect 234 47 313 55
rect 496 49 550 131
rect 580 91 660 177
rect 580 57 590 91
rect 624 57 660 91
rect 580 49 660 57
rect 690 169 789 177
rect 690 135 742 169
rect 776 135 789 169
rect 690 49 789 135
rect 862 157 922 177
rect 862 123 878 157
rect 912 123 922 157
rect 862 89 922 123
rect 862 55 878 89
rect 912 55 922 89
rect 862 47 922 55
rect 952 161 1004 177
rect 952 127 962 161
rect 996 127 1004 161
rect 952 121 1004 127
rect 952 47 1002 121
rect 1058 105 1108 177
rect 1056 97 1108 105
rect 1056 63 1064 97
rect 1098 63 1108 97
rect 1056 49 1108 63
rect 1138 133 1239 177
rect 1315 169 1419 177
rect 1315 135 1361 169
rect 1395 135 1419 169
rect 1315 133 1419 135
rect 1138 126 1260 133
rect 1138 92 1148 126
rect 1182 92 1260 126
rect 1138 49 1260 92
rect 1290 49 1419 133
rect 1449 167 1499 177
rect 1589 167 1639 175
rect 1449 93 1539 167
rect 1449 59 1461 93
rect 1495 59 1539 93
rect 1449 49 1539 59
rect 1466 47 1539 49
rect 1569 142 1639 167
rect 1569 108 1595 142
rect 1629 108 1639 142
rect 1569 47 1639 108
rect 1669 97 1723 175
rect 1669 63 1679 97
rect 1713 63 1723 97
rect 1669 47 1723 63
rect 1753 101 1805 175
rect 1753 67 1763 101
rect 1797 67 1805 101
rect 1753 47 1805 67
<< pdiff >>
rect 72 477 124 497
rect 72 443 80 477
rect 114 443 124 477
rect 72 297 124 443
rect 154 477 208 497
rect 154 443 164 477
rect 198 443 208 477
rect 154 409 208 443
rect 154 375 164 409
rect 198 375 208 409
rect 154 341 208 375
rect 154 307 164 341
rect 198 307 208 341
rect 154 297 208 307
rect 238 477 313 497
rect 238 443 265 477
rect 299 443 313 477
rect 238 425 313 443
rect 238 297 328 425
rect 358 341 414 425
rect 358 307 368 341
rect 402 307 414 341
rect 478 413 542 493
rect 478 379 498 413
rect 532 379 542 413
rect 478 325 542 379
rect 572 481 648 493
rect 572 447 591 481
rect 625 447 648 481
rect 572 325 648 447
rect 678 481 783 493
rect 678 447 738 481
rect 772 447 783 481
rect 678 325 783 447
rect 837 481 889 497
rect 837 447 845 481
rect 879 447 889 481
rect 358 297 414 307
rect 837 297 889 447
rect 919 349 969 497
rect 1023 405 1108 465
rect 1023 371 1031 405
rect 1065 371 1108 405
rect 1023 365 1108 371
rect 919 343 971 349
rect 919 309 929 343
rect 963 309 971 343
rect 919 297 971 309
rect 1025 297 1108 365
rect 1138 425 1238 465
rect 1480 489 1538 497
rect 1480 457 1492 489
rect 1350 425 1435 457
rect 1138 409 1260 425
rect 1138 375 1189 409
rect 1223 375 1260 409
rect 1138 341 1260 375
rect 1138 307 1189 341
rect 1223 307 1260 341
rect 1138 297 1260 307
rect 1290 421 1435 425
rect 1290 387 1391 421
rect 1425 387 1435 421
rect 1290 329 1435 387
rect 1465 455 1492 457
rect 1526 455 1538 489
rect 1465 329 1538 455
rect 1568 341 1639 497
rect 1568 329 1595 341
rect 1290 297 1385 329
rect 1583 307 1595 329
rect 1629 307 1639 341
rect 1583 297 1639 307
rect 1669 489 1723 497
rect 1669 455 1679 489
rect 1713 455 1723 489
rect 1669 297 1723 455
rect 1753 477 1806 497
rect 1753 443 1764 477
rect 1798 443 1806 477
rect 1753 409 1806 443
rect 1753 375 1764 409
rect 1798 375 1806 409
rect 1753 297 1806 375
<< ndiffc >>
rect 76 59 110 93
rect 160 95 194 129
rect 396 135 430 169
rect 506 131 540 165
rect 260 55 294 89
rect 590 57 624 91
rect 742 135 776 169
rect 878 123 912 157
rect 878 55 912 89
rect 962 127 996 161
rect 1064 63 1098 97
rect 1361 135 1395 169
rect 1148 92 1182 126
rect 1461 59 1495 93
rect 1595 108 1629 142
rect 1679 63 1713 97
rect 1763 67 1797 101
<< pdiffc >>
rect 80 443 114 477
rect 164 443 198 477
rect 164 375 198 409
rect 164 307 198 341
rect 265 443 299 477
rect 368 307 402 341
rect 498 379 532 413
rect 591 447 625 481
rect 738 447 772 481
rect 845 447 879 481
rect 1031 371 1065 405
rect 929 309 963 343
rect 1189 375 1223 409
rect 1189 307 1223 341
rect 1391 387 1425 421
rect 1492 455 1526 489
rect 1595 307 1629 341
rect 1679 455 1713 489
rect 1764 443 1798 477
rect 1764 375 1798 409
<< poly >>
rect 124 497 154 523
rect 208 497 238 523
rect 542 493 572 519
rect 648 493 678 519
rect 889 497 919 523
rect 328 425 358 483
rect 124 265 154 297
rect 208 265 238 297
rect 328 265 358 297
rect 542 271 572 325
rect 542 265 581 271
rect 648 265 678 325
rect 1108 493 1465 523
rect 1538 497 1568 523
rect 1639 497 1669 523
rect 1723 497 1753 523
rect 1108 465 1138 493
rect 1435 457 1465 493
rect 1260 425 1290 451
rect 120 249 286 265
rect 120 215 242 249
rect 276 215 286 249
rect 120 199 286 215
rect 328 249 581 265
rect 328 215 469 249
rect 503 215 537 249
rect 571 215 581 249
rect 328 199 581 215
rect 636 249 690 265
rect 636 215 646 249
rect 680 215 690 249
rect 889 247 919 297
rect 1108 247 1138 297
rect 1260 265 1290 297
rect 1435 265 1465 329
rect 889 217 1138 247
rect 636 199 690 215
rect 120 177 150 199
rect 204 177 234 199
rect 328 177 358 199
rect 550 197 581 199
rect 550 177 580 197
rect 660 177 690 199
rect 922 177 952 217
rect 1108 177 1138 217
rect 1180 249 1290 265
rect 1180 215 1190 249
rect 1224 215 1290 249
rect 1180 199 1290 215
rect 328 67 358 93
rect 120 21 150 47
rect 204 21 234 47
rect 550 21 580 49
rect 660 21 690 49
rect 1260 133 1290 199
rect 1419 249 1473 265
rect 1538 256 1568 329
rect 1639 265 1669 297
rect 1723 265 1753 297
rect 1538 255 1569 256
rect 1419 215 1429 249
rect 1463 215 1473 249
rect 1419 199 1473 215
rect 1515 239 1569 255
rect 1515 205 1525 239
rect 1559 205 1569 239
rect 1419 177 1449 199
rect 1515 189 1569 205
rect 1611 249 1669 265
rect 1611 215 1621 249
rect 1655 215 1669 249
rect 1611 199 1669 215
rect 1711 249 1765 265
rect 1711 215 1721 249
rect 1755 215 1765 249
rect 1711 199 1765 215
rect 1539 167 1569 189
rect 1639 175 1669 199
rect 1723 175 1753 199
rect 922 21 952 47
rect 1108 21 1138 49
rect 1260 23 1290 49
rect 1419 21 1449 49
rect 1539 21 1569 47
rect 1639 21 1669 47
rect 1723 21 1753 47
<< polycont >>
rect 242 215 276 249
rect 469 215 503 249
rect 537 215 571 249
rect 646 215 680 249
rect 1190 215 1224 249
rect 1429 215 1463 249
rect 1525 205 1559 239
rect 1621 215 1655 249
rect 1721 215 1755 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1840 561
rect 60 477 130 527
rect 60 443 80 477
rect 114 443 130 477
rect 164 477 214 493
rect 198 443 214 477
rect 248 477 315 527
rect 829 481 895 527
rect 1663 489 1730 527
rect 248 443 265 477
rect 299 443 315 477
rect 352 447 591 481
rect 625 447 671 481
rect 714 447 738 481
rect 772 447 795 481
rect 829 447 845 481
rect 879 447 895 481
rect 962 455 1492 489
rect 1526 455 1581 489
rect 1663 455 1679 489
rect 1713 455 1730 489
rect 1764 477 1823 493
rect 164 409 214 443
rect 352 409 386 447
rect 761 413 795 447
rect 962 413 996 455
rect 109 375 164 409
rect 198 375 214 409
rect 109 341 214 375
rect 109 307 164 341
rect 198 307 214 341
rect 109 288 214 307
rect 248 375 386 409
rect 466 379 498 413
rect 532 379 727 413
rect 761 379 996 413
rect 1031 405 1065 421
rect 109 185 172 288
rect 248 265 282 375
rect 329 307 368 341
rect 402 307 659 341
rect 242 249 282 265
rect 276 215 282 249
rect 242 199 282 215
rect 109 132 210 185
rect 248 173 282 199
rect 248 139 362 173
rect 160 129 210 132
rect 194 95 210 129
rect 60 59 76 93
rect 110 59 126 93
rect 160 70 210 95
rect 244 89 294 105
rect 60 17 126 59
rect 244 55 260 89
rect 244 17 294 55
rect 328 85 362 139
rect 396 169 430 307
rect 625 265 659 307
rect 693 339 727 379
rect 693 323 799 339
rect 693 305 765 323
rect 742 289 765 305
rect 742 275 799 289
rect 464 249 591 265
rect 464 215 469 249
rect 503 215 537 249
rect 571 215 591 249
rect 464 199 591 215
rect 625 249 680 265
rect 625 215 646 249
rect 625 199 680 215
rect 742 169 776 275
rect 833 241 867 379
rect 913 309 929 343
rect 963 309 996 343
rect 913 289 996 309
rect 396 119 430 135
rect 486 131 506 165
rect 540 131 708 165
rect 570 85 590 91
rect 328 57 590 85
rect 624 57 640 91
rect 328 51 640 57
rect 674 85 708 131
rect 742 119 776 135
rect 810 207 867 241
rect 810 85 844 207
rect 948 187 996 289
rect 674 51 844 85
rect 878 157 912 173
rect 878 89 912 123
rect 948 153 949 187
rect 983 161 996 187
rect 948 127 962 153
rect 948 83 996 127
rect 1031 119 1065 371
rect 1099 178 1133 455
rect 1798 443 1823 477
rect 1764 421 1823 443
rect 1171 375 1189 409
rect 1223 375 1254 409
rect 1171 341 1254 375
rect 1171 307 1189 341
rect 1223 323 1254 341
rect 1361 387 1391 421
rect 1425 409 1823 421
rect 1425 387 1764 409
rect 1223 307 1225 323
rect 1171 289 1225 307
rect 1259 289 1327 323
rect 1174 249 1259 254
rect 1174 215 1190 249
rect 1224 215 1259 249
rect 1174 199 1259 215
rect 1216 187 1259 199
rect 1099 165 1143 178
rect 1099 144 1182 165
rect 1109 131 1182 144
rect 1148 126 1182 131
rect 1216 153 1225 187
rect 1216 126 1259 153
rect 1031 85 1041 119
rect 878 17 912 55
rect 1031 63 1064 85
rect 1098 63 1114 97
rect 1148 64 1182 92
rect 1293 85 1327 289
rect 1361 169 1395 387
rect 1726 375 1764 387
rect 1798 375 1823 409
rect 1429 289 1545 323
rect 1579 307 1595 341
rect 1629 307 1743 341
rect 1579 299 1743 307
rect 1429 249 1463 289
rect 1709 265 1743 299
rect 1429 199 1463 215
rect 1497 239 1559 255
rect 1497 205 1525 239
rect 1593 249 1675 265
rect 1593 215 1621 249
rect 1655 215 1675 249
rect 1709 249 1755 265
rect 1709 215 1721 249
rect 1497 189 1559 205
rect 1709 199 1755 215
rect 1497 187 1538 189
rect 1497 153 1501 187
rect 1535 153 1538 187
rect 1709 181 1743 199
rect 1497 146 1538 153
rect 1595 150 1743 181
rect 1587 147 1743 150
rect 1361 119 1395 135
rect 1587 142 1645 147
rect 1587 119 1595 142
rect 1429 85 1461 93
rect 1031 53 1114 63
rect 1293 59 1461 85
rect 1495 59 1522 93
rect 1587 85 1593 119
rect 1629 108 1645 142
rect 1789 117 1823 375
rect 1627 85 1645 108
rect 1587 59 1645 85
rect 1679 97 1713 113
rect 1293 51 1522 59
rect 1679 17 1713 63
rect 1763 101 1823 117
rect 1797 67 1823 101
rect 1763 51 1823 67
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1840 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 765 289 799 323
rect 949 161 983 187
rect 949 153 962 161
rect 962 153 983 161
rect 1225 289 1259 323
rect 1225 153 1259 187
rect 1041 97 1075 119
rect 1041 85 1064 97
rect 1064 85 1075 97
rect 1501 153 1535 187
rect 1593 108 1595 119
rect 1595 108 1627 119
rect 1593 85 1627 108
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
<< metal1 >>
rect 0 561 1840 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1840 561
rect 0 496 1840 527
rect 753 323 811 329
rect 753 289 765 323
rect 799 320 811 323
rect 1213 323 1271 329
rect 1213 320 1225 323
rect 799 292 1225 320
rect 799 289 811 292
rect 753 283 811 289
rect 1213 289 1225 292
rect 1259 289 1271 323
rect 1213 283 1271 289
rect 937 187 995 193
rect 937 153 949 187
rect 983 184 995 187
rect 1213 187 1271 193
rect 1213 184 1225 187
rect 983 156 1225 184
rect 983 153 995 156
rect 937 147 995 153
rect 1213 153 1225 156
rect 1259 184 1271 187
rect 1489 187 1547 193
rect 1489 184 1501 187
rect 1259 156 1501 184
rect 1259 153 1271 156
rect 1213 147 1271 153
rect 1489 153 1501 156
rect 1535 153 1547 187
rect 1489 147 1547 153
rect 1029 119 1087 125
rect 1029 85 1041 119
rect 1075 116 1087 119
rect 1581 119 1639 125
rect 1581 116 1593 119
rect 1075 88 1593 116
rect 1075 85 1087 88
rect 1029 79 1087 85
rect 1581 85 1593 88
rect 1627 85 1639 119
rect 1581 79 1639 85
rect 0 17 1840 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1840 17
rect 0 -48 1840 -17
<< labels >>
flabel locali s 121 357 155 391 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 489 221 523 255 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 1501 289 1535 323 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 1593 221 1627 255 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 hkscl5hdv1_xor3_1
flabel comment s 0 544 0 544 3 FreeSans 200 0 0 0 HHNEC
rlabel metal1 s 0 -48 1840 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1840 592 1 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1840 544
string GDS_END 685594
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 673288
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 9.200 0.000 
<< end >>
