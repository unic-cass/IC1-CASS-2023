magic
tech sky130A
magscale 1 2
timestamp 1699127393
<< obsli1 >>
rect 1104 2159 98808 97393
<< obsm1 >>
rect 934 76 98808 99136
<< metal2 >>
rect 2502 99200 2558 100000
rect 6458 99200 6514 100000
rect 10414 99200 10470 100000
rect 14370 99200 14426 100000
rect 18326 99200 18382 100000
rect 22282 99200 22338 100000
rect 26238 99200 26294 100000
rect 30194 99200 30250 100000
rect 34150 99200 34206 100000
rect 38106 99200 38162 100000
rect 42062 99200 42118 100000
rect 46018 99200 46074 100000
rect 49974 99200 50030 100000
rect 53930 99200 53986 100000
rect 57886 99200 57942 100000
rect 61842 99200 61898 100000
rect 65798 99200 65854 100000
rect 69754 99200 69810 100000
rect 73710 99200 73766 100000
rect 77666 99200 77722 100000
rect 81622 99200 81678 100000
rect 85578 99200 85634 100000
rect 89534 99200 89590 100000
rect 93490 99200 93546 100000
rect 97446 99200 97502 100000
rect 3054 0 3110 800
rect 4434 0 4490 800
rect 5814 0 5870 800
rect 7194 0 7250 800
rect 8574 0 8630 800
rect 9954 0 10010 800
rect 11334 0 11390 800
rect 12714 0 12770 800
rect 14094 0 14150 800
rect 15474 0 15530 800
rect 16854 0 16910 800
rect 18234 0 18290 800
rect 19614 0 19670 800
rect 20994 0 21050 800
rect 22374 0 22430 800
rect 23754 0 23810 800
rect 25134 0 25190 800
rect 26514 0 26570 800
rect 27894 0 27950 800
rect 29274 0 29330 800
rect 30654 0 30710 800
rect 32034 0 32090 800
rect 33414 0 33470 800
rect 34794 0 34850 800
rect 36174 0 36230 800
rect 37554 0 37610 800
rect 38934 0 38990 800
rect 40314 0 40370 800
rect 41694 0 41750 800
rect 43074 0 43130 800
rect 44454 0 44510 800
rect 45834 0 45890 800
rect 47214 0 47270 800
rect 48594 0 48650 800
rect 49974 0 50030 800
rect 51354 0 51410 800
rect 52734 0 52790 800
rect 54114 0 54170 800
rect 55494 0 55550 800
rect 56874 0 56930 800
rect 58254 0 58310 800
rect 59634 0 59690 800
rect 61014 0 61070 800
rect 62394 0 62450 800
rect 63774 0 63830 800
rect 65154 0 65210 800
rect 66534 0 66590 800
rect 67914 0 67970 800
rect 69294 0 69350 800
rect 70674 0 70730 800
rect 72054 0 72110 800
rect 73434 0 73490 800
rect 74814 0 74870 800
rect 76194 0 76250 800
rect 77574 0 77630 800
rect 78954 0 79010 800
rect 80334 0 80390 800
rect 81714 0 81770 800
rect 83094 0 83150 800
rect 84474 0 84530 800
rect 85854 0 85910 800
rect 87234 0 87290 800
rect 88614 0 88670 800
rect 89994 0 90050 800
rect 91374 0 91430 800
rect 92754 0 92810 800
rect 94134 0 94190 800
rect 95514 0 95570 800
rect 96894 0 96950 800
<< obsm2 >>
rect 938 99144 2446 99362
rect 2614 99144 6402 99362
rect 6570 99144 10358 99362
rect 10526 99144 14314 99362
rect 14482 99144 18270 99362
rect 18438 99144 22226 99362
rect 22394 99144 26182 99362
rect 26350 99144 30138 99362
rect 30306 99144 34094 99362
rect 34262 99144 38050 99362
rect 38218 99144 42006 99362
rect 42174 99144 45962 99362
rect 46130 99144 49918 99362
rect 50086 99144 53874 99362
rect 54042 99144 57830 99362
rect 57998 99144 61786 99362
rect 61954 99144 65742 99362
rect 65910 99144 69698 99362
rect 69866 99144 73654 99362
rect 73822 99144 77610 99362
rect 77778 99144 81566 99362
rect 81734 99144 85522 99362
rect 85690 99144 89478 99362
rect 89646 99144 93434 99362
rect 93602 99144 97390 99362
rect 97558 99144 98144 99362
rect 938 856 98144 99144
rect 938 70 2998 856
rect 3166 70 4378 856
rect 4546 70 5758 856
rect 5926 70 7138 856
rect 7306 70 8518 856
rect 8686 70 9898 856
rect 10066 70 11278 856
rect 11446 70 12658 856
rect 12826 70 14038 856
rect 14206 70 15418 856
rect 15586 70 16798 856
rect 16966 70 18178 856
rect 18346 70 19558 856
rect 19726 70 20938 856
rect 21106 70 22318 856
rect 22486 70 23698 856
rect 23866 70 25078 856
rect 25246 70 26458 856
rect 26626 70 27838 856
rect 28006 70 29218 856
rect 29386 70 30598 856
rect 30766 70 31978 856
rect 32146 70 33358 856
rect 33526 70 34738 856
rect 34906 70 36118 856
rect 36286 70 37498 856
rect 37666 70 38878 856
rect 39046 70 40258 856
rect 40426 70 41638 856
rect 41806 70 43018 856
rect 43186 70 44398 856
rect 44566 70 45778 856
rect 45946 70 47158 856
rect 47326 70 48538 856
rect 48706 70 49918 856
rect 50086 70 51298 856
rect 51466 70 52678 856
rect 52846 70 54058 856
rect 54226 70 55438 856
rect 55606 70 56818 856
rect 56986 70 58198 856
rect 58366 70 59578 856
rect 59746 70 60958 856
rect 61126 70 62338 856
rect 62506 70 63718 856
rect 63886 70 65098 856
rect 65266 70 66478 856
rect 66646 70 67858 856
rect 68026 70 69238 856
rect 69406 70 70618 856
rect 70786 70 71998 856
rect 72166 70 73378 856
rect 73546 70 74758 856
rect 74926 70 76138 856
rect 76306 70 77518 856
rect 77686 70 78898 856
rect 79066 70 80278 856
rect 80446 70 81658 856
rect 81826 70 83038 856
rect 83206 70 84418 856
rect 84586 70 85798 856
rect 85966 70 87178 856
rect 87346 70 88558 856
rect 88726 70 89938 856
rect 90106 70 91318 856
rect 91486 70 92698 856
rect 92866 70 94078 856
rect 94246 70 95458 856
rect 95626 70 96838 856
rect 97006 70 98144 856
<< metal3 >>
rect 0 96976 800 97096
rect 0 94120 800 94240
rect 0 91264 800 91384
rect 0 88408 800 88528
rect 0 85552 800 85672
rect 0 82696 800 82816
rect 0 79840 800 79960
rect 0 76984 800 77104
rect 0 74128 800 74248
rect 0 71272 800 71392
rect 0 68416 800 68536
rect 0 65560 800 65680
rect 0 62704 800 62824
rect 0 59848 800 59968
rect 0 56992 800 57112
rect 0 54136 800 54256
rect 0 51280 800 51400
rect 0 48424 800 48544
rect 0 45568 800 45688
rect 0 42712 800 42832
rect 0 39856 800 39976
rect 0 37000 800 37120
rect 0 34144 800 34264
rect 0 31288 800 31408
rect 0 28432 800 28552
rect 0 25576 800 25696
rect 0 22720 800 22840
rect 0 19864 800 19984
rect 0 17008 800 17128
rect 0 14152 800 14272
rect 0 11296 800 11416
rect 0 8440 800 8560
rect 0 5584 800 5704
rect 0 2728 800 2848
<< obsm3 >>
rect 800 97176 98059 97409
rect 880 96896 98059 97176
rect 800 94320 98059 96896
rect 880 94040 98059 94320
rect 800 91464 98059 94040
rect 880 91184 98059 91464
rect 800 88608 98059 91184
rect 880 88328 98059 88608
rect 800 85752 98059 88328
rect 880 85472 98059 85752
rect 800 82896 98059 85472
rect 880 82616 98059 82896
rect 800 80040 98059 82616
rect 880 79760 98059 80040
rect 800 77184 98059 79760
rect 880 76904 98059 77184
rect 800 74328 98059 76904
rect 880 74048 98059 74328
rect 800 71472 98059 74048
rect 880 71192 98059 71472
rect 800 68616 98059 71192
rect 880 68336 98059 68616
rect 800 65760 98059 68336
rect 880 65480 98059 65760
rect 800 62904 98059 65480
rect 880 62624 98059 62904
rect 800 60048 98059 62624
rect 880 59768 98059 60048
rect 800 57192 98059 59768
rect 880 56912 98059 57192
rect 800 54336 98059 56912
rect 880 54056 98059 54336
rect 800 51480 98059 54056
rect 880 51200 98059 51480
rect 800 48624 98059 51200
rect 880 48344 98059 48624
rect 800 45768 98059 48344
rect 880 45488 98059 45768
rect 800 42912 98059 45488
rect 880 42632 98059 42912
rect 800 40056 98059 42632
rect 880 39776 98059 40056
rect 800 37200 98059 39776
rect 880 36920 98059 37200
rect 800 34344 98059 36920
rect 880 34064 98059 34344
rect 800 31488 98059 34064
rect 880 31208 98059 31488
rect 800 28632 98059 31208
rect 880 28352 98059 28632
rect 800 25776 98059 28352
rect 880 25496 98059 25776
rect 800 22920 98059 25496
rect 880 22640 98059 22920
rect 800 20064 98059 22640
rect 880 19784 98059 20064
rect 800 17208 98059 19784
rect 880 16928 98059 17208
rect 800 14352 98059 16928
rect 880 14072 98059 14352
rect 800 11496 98059 14072
rect 880 11216 98059 11496
rect 800 8640 98059 11216
rect 880 8360 98059 8640
rect 800 5784 98059 8360
rect 880 5504 98059 5784
rect 800 2928 98059 5504
rect 880 2648 98059 2928
rect 800 1667 98059 2648
<< metal4 >>
rect 4208 2128 4528 97424
rect 19568 2128 19888 97424
rect 34928 2128 35248 97424
rect 50288 2128 50608 97424
rect 65648 2128 65968 97424
rect 81008 2128 81328 97424
rect 96368 2128 96688 97424
<< obsm4 >>
rect 13675 2347 19488 96933
rect 19968 2347 34848 96933
rect 35328 2347 50208 96933
rect 50688 2347 65568 96933
rect 66048 2347 80928 96933
rect 81408 2347 96288 96933
rect 96768 2347 97829 96933
<< labels >>
rlabel metal2 s 2502 99200 2558 100000 6 buttons
port 1 nsew signal input
rlabel metal2 s 3054 0 3110 800 6 clk
port 2 nsew signal input
rlabel metal2 s 9954 0 10010 800 6 i_wb_addr[0]
port 3 nsew signal input
rlabel metal2 s 23754 0 23810 800 6 i_wb_addr[10]
port 4 nsew signal input
rlabel metal2 s 25134 0 25190 800 6 i_wb_addr[11]
port 5 nsew signal input
rlabel metal2 s 26514 0 26570 800 6 i_wb_addr[12]
port 6 nsew signal input
rlabel metal2 s 27894 0 27950 800 6 i_wb_addr[13]
port 7 nsew signal input
rlabel metal2 s 29274 0 29330 800 6 i_wb_addr[14]
port 8 nsew signal input
rlabel metal2 s 30654 0 30710 800 6 i_wb_addr[15]
port 9 nsew signal input
rlabel metal2 s 32034 0 32090 800 6 i_wb_addr[16]
port 10 nsew signal input
rlabel metal2 s 33414 0 33470 800 6 i_wb_addr[17]
port 11 nsew signal input
rlabel metal2 s 34794 0 34850 800 6 i_wb_addr[18]
port 12 nsew signal input
rlabel metal2 s 36174 0 36230 800 6 i_wb_addr[19]
port 13 nsew signal input
rlabel metal2 s 11334 0 11390 800 6 i_wb_addr[1]
port 14 nsew signal input
rlabel metal2 s 37554 0 37610 800 6 i_wb_addr[20]
port 15 nsew signal input
rlabel metal2 s 38934 0 38990 800 6 i_wb_addr[21]
port 16 nsew signal input
rlabel metal2 s 40314 0 40370 800 6 i_wb_addr[22]
port 17 nsew signal input
rlabel metal2 s 41694 0 41750 800 6 i_wb_addr[23]
port 18 nsew signal input
rlabel metal2 s 43074 0 43130 800 6 i_wb_addr[24]
port 19 nsew signal input
rlabel metal2 s 44454 0 44510 800 6 i_wb_addr[25]
port 20 nsew signal input
rlabel metal2 s 45834 0 45890 800 6 i_wb_addr[26]
port 21 nsew signal input
rlabel metal2 s 47214 0 47270 800 6 i_wb_addr[27]
port 22 nsew signal input
rlabel metal2 s 48594 0 48650 800 6 i_wb_addr[28]
port 23 nsew signal input
rlabel metal2 s 49974 0 50030 800 6 i_wb_addr[29]
port 24 nsew signal input
rlabel metal2 s 12714 0 12770 800 6 i_wb_addr[2]
port 25 nsew signal input
rlabel metal2 s 51354 0 51410 800 6 i_wb_addr[30]
port 26 nsew signal input
rlabel metal2 s 52734 0 52790 800 6 i_wb_addr[31]
port 27 nsew signal input
rlabel metal2 s 14094 0 14150 800 6 i_wb_addr[3]
port 28 nsew signal input
rlabel metal2 s 15474 0 15530 800 6 i_wb_addr[4]
port 29 nsew signal input
rlabel metal2 s 16854 0 16910 800 6 i_wb_addr[5]
port 30 nsew signal input
rlabel metal2 s 18234 0 18290 800 6 i_wb_addr[6]
port 31 nsew signal input
rlabel metal2 s 19614 0 19670 800 6 i_wb_addr[7]
port 32 nsew signal input
rlabel metal2 s 20994 0 21050 800 6 i_wb_addr[8]
port 33 nsew signal input
rlabel metal2 s 22374 0 22430 800 6 i_wb_addr[9]
port 34 nsew signal input
rlabel metal2 s 5814 0 5870 800 6 i_wb_cyc
port 35 nsew signal input
rlabel metal2 s 54114 0 54170 800 6 i_wb_data[0]
port 36 nsew signal input
rlabel metal2 s 67914 0 67970 800 6 i_wb_data[10]
port 37 nsew signal input
rlabel metal2 s 69294 0 69350 800 6 i_wb_data[11]
port 38 nsew signal input
rlabel metal2 s 70674 0 70730 800 6 i_wb_data[12]
port 39 nsew signal input
rlabel metal2 s 72054 0 72110 800 6 i_wb_data[13]
port 40 nsew signal input
rlabel metal2 s 73434 0 73490 800 6 i_wb_data[14]
port 41 nsew signal input
rlabel metal2 s 74814 0 74870 800 6 i_wb_data[15]
port 42 nsew signal input
rlabel metal2 s 76194 0 76250 800 6 i_wb_data[16]
port 43 nsew signal input
rlabel metal2 s 77574 0 77630 800 6 i_wb_data[17]
port 44 nsew signal input
rlabel metal2 s 78954 0 79010 800 6 i_wb_data[18]
port 45 nsew signal input
rlabel metal2 s 80334 0 80390 800 6 i_wb_data[19]
port 46 nsew signal input
rlabel metal2 s 55494 0 55550 800 6 i_wb_data[1]
port 47 nsew signal input
rlabel metal2 s 81714 0 81770 800 6 i_wb_data[20]
port 48 nsew signal input
rlabel metal2 s 83094 0 83150 800 6 i_wb_data[21]
port 49 nsew signal input
rlabel metal2 s 84474 0 84530 800 6 i_wb_data[22]
port 50 nsew signal input
rlabel metal2 s 85854 0 85910 800 6 i_wb_data[23]
port 51 nsew signal input
rlabel metal2 s 87234 0 87290 800 6 i_wb_data[24]
port 52 nsew signal input
rlabel metal2 s 88614 0 88670 800 6 i_wb_data[25]
port 53 nsew signal input
rlabel metal2 s 89994 0 90050 800 6 i_wb_data[26]
port 54 nsew signal input
rlabel metal2 s 91374 0 91430 800 6 i_wb_data[27]
port 55 nsew signal input
rlabel metal2 s 92754 0 92810 800 6 i_wb_data[28]
port 56 nsew signal input
rlabel metal2 s 94134 0 94190 800 6 i_wb_data[29]
port 57 nsew signal input
rlabel metal2 s 56874 0 56930 800 6 i_wb_data[2]
port 58 nsew signal input
rlabel metal2 s 95514 0 95570 800 6 i_wb_data[30]
port 59 nsew signal input
rlabel metal2 s 96894 0 96950 800 6 i_wb_data[31]
port 60 nsew signal input
rlabel metal2 s 58254 0 58310 800 6 i_wb_data[3]
port 61 nsew signal input
rlabel metal2 s 59634 0 59690 800 6 i_wb_data[4]
port 62 nsew signal input
rlabel metal2 s 61014 0 61070 800 6 i_wb_data[5]
port 63 nsew signal input
rlabel metal2 s 62394 0 62450 800 6 i_wb_data[6]
port 64 nsew signal input
rlabel metal2 s 63774 0 63830 800 6 i_wb_data[7]
port 65 nsew signal input
rlabel metal2 s 65154 0 65210 800 6 i_wb_data[8]
port 66 nsew signal input
rlabel metal2 s 66534 0 66590 800 6 i_wb_data[9]
port 67 nsew signal input
rlabel metal2 s 7194 0 7250 800 6 i_wb_stb
port 68 nsew signal input
rlabel metal2 s 8574 0 8630 800 6 i_wb_we
port 69 nsew signal input
rlabel metal2 s 6458 99200 6514 100000 6 led_enb[0]
port 70 nsew signal output
rlabel metal2 s 46018 99200 46074 100000 6 led_enb[10]
port 71 nsew signal output
rlabel metal2 s 49974 99200 50030 100000 6 led_enb[11]
port 72 nsew signal output
rlabel metal2 s 10414 99200 10470 100000 6 led_enb[1]
port 73 nsew signal output
rlabel metal2 s 14370 99200 14426 100000 6 led_enb[2]
port 74 nsew signal output
rlabel metal2 s 18326 99200 18382 100000 6 led_enb[3]
port 75 nsew signal output
rlabel metal2 s 22282 99200 22338 100000 6 led_enb[4]
port 76 nsew signal output
rlabel metal2 s 26238 99200 26294 100000 6 led_enb[5]
port 77 nsew signal output
rlabel metal2 s 30194 99200 30250 100000 6 led_enb[6]
port 78 nsew signal output
rlabel metal2 s 34150 99200 34206 100000 6 led_enb[7]
port 79 nsew signal output
rlabel metal2 s 38106 99200 38162 100000 6 led_enb[8]
port 80 nsew signal output
rlabel metal2 s 42062 99200 42118 100000 6 led_enb[9]
port 81 nsew signal output
rlabel metal2 s 53930 99200 53986 100000 6 leds[0]
port 82 nsew signal output
rlabel metal2 s 93490 99200 93546 100000 6 leds[10]
port 83 nsew signal output
rlabel metal2 s 97446 99200 97502 100000 6 leds[11]
port 84 nsew signal output
rlabel metal2 s 57886 99200 57942 100000 6 leds[1]
port 85 nsew signal output
rlabel metal2 s 61842 99200 61898 100000 6 leds[2]
port 86 nsew signal output
rlabel metal2 s 65798 99200 65854 100000 6 leds[3]
port 87 nsew signal output
rlabel metal2 s 69754 99200 69810 100000 6 leds[4]
port 88 nsew signal output
rlabel metal2 s 73710 99200 73766 100000 6 leds[5]
port 89 nsew signal output
rlabel metal2 s 77666 99200 77722 100000 6 leds[6]
port 90 nsew signal output
rlabel metal2 s 81622 99200 81678 100000 6 leds[7]
port 91 nsew signal output
rlabel metal2 s 85578 99200 85634 100000 6 leds[8]
port 92 nsew signal output
rlabel metal2 s 89534 99200 89590 100000 6 leds[9]
port 93 nsew signal output
rlabel metal3 s 0 2728 800 2848 6 o_wb_ack
port 94 nsew signal output
rlabel metal3 s 0 8440 800 8560 6 o_wb_data[0]
port 95 nsew signal output
rlabel metal3 s 0 37000 800 37120 6 o_wb_data[10]
port 96 nsew signal output
rlabel metal3 s 0 39856 800 39976 6 o_wb_data[11]
port 97 nsew signal output
rlabel metal3 s 0 42712 800 42832 6 o_wb_data[12]
port 98 nsew signal output
rlabel metal3 s 0 45568 800 45688 6 o_wb_data[13]
port 99 nsew signal output
rlabel metal3 s 0 48424 800 48544 6 o_wb_data[14]
port 100 nsew signal output
rlabel metal3 s 0 51280 800 51400 6 o_wb_data[15]
port 101 nsew signal output
rlabel metal3 s 0 54136 800 54256 6 o_wb_data[16]
port 102 nsew signal output
rlabel metal3 s 0 56992 800 57112 6 o_wb_data[17]
port 103 nsew signal output
rlabel metal3 s 0 59848 800 59968 6 o_wb_data[18]
port 104 nsew signal output
rlabel metal3 s 0 62704 800 62824 6 o_wb_data[19]
port 105 nsew signal output
rlabel metal3 s 0 11296 800 11416 6 o_wb_data[1]
port 106 nsew signal output
rlabel metal3 s 0 65560 800 65680 6 o_wb_data[20]
port 107 nsew signal output
rlabel metal3 s 0 68416 800 68536 6 o_wb_data[21]
port 108 nsew signal output
rlabel metal3 s 0 71272 800 71392 6 o_wb_data[22]
port 109 nsew signal output
rlabel metal3 s 0 74128 800 74248 6 o_wb_data[23]
port 110 nsew signal output
rlabel metal3 s 0 76984 800 77104 6 o_wb_data[24]
port 111 nsew signal output
rlabel metal3 s 0 79840 800 79960 6 o_wb_data[25]
port 112 nsew signal output
rlabel metal3 s 0 82696 800 82816 6 o_wb_data[26]
port 113 nsew signal output
rlabel metal3 s 0 85552 800 85672 6 o_wb_data[27]
port 114 nsew signal output
rlabel metal3 s 0 88408 800 88528 6 o_wb_data[28]
port 115 nsew signal output
rlabel metal3 s 0 91264 800 91384 6 o_wb_data[29]
port 116 nsew signal output
rlabel metal3 s 0 14152 800 14272 6 o_wb_data[2]
port 117 nsew signal output
rlabel metal3 s 0 94120 800 94240 6 o_wb_data[30]
port 118 nsew signal output
rlabel metal3 s 0 96976 800 97096 6 o_wb_data[31]
port 119 nsew signal output
rlabel metal3 s 0 17008 800 17128 6 o_wb_data[3]
port 120 nsew signal output
rlabel metal3 s 0 19864 800 19984 6 o_wb_data[4]
port 121 nsew signal output
rlabel metal3 s 0 22720 800 22840 6 o_wb_data[5]
port 122 nsew signal output
rlabel metal3 s 0 25576 800 25696 6 o_wb_data[6]
port 123 nsew signal output
rlabel metal3 s 0 28432 800 28552 6 o_wb_data[7]
port 124 nsew signal output
rlabel metal3 s 0 31288 800 31408 6 o_wb_data[8]
port 125 nsew signal output
rlabel metal3 s 0 34144 800 34264 6 o_wb_data[9]
port 126 nsew signal output
rlabel metal3 s 0 5584 800 5704 6 o_wb_stall
port 127 nsew signal output
rlabel metal2 s 4434 0 4490 800 6 reset
port 128 nsew signal input
rlabel metal4 s 4208 2128 4528 97424 6 vccd1
port 129 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 97424 6 vccd1
port 129 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 97424 6 vccd1
port 129 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 97424 6 vccd1
port 129 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 97424 6 vssd1
port 130 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 97424 6 vssd1
port 130 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 97424 6 vssd1
port 130 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 100000 100000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 26653208
string GDS_FILE /home/rodrigowue/test/IC1-CASS-2023/openlane/wb_buttons_leds/runs/23_11_04_16_42/results/signoff/wb_buttons_leds.magic.gds
string GDS_START 1162660
<< end >>

