magic
tech sky130B
magscale 1 2
timestamp 1676037725
<< nwell >>
rect -38 261 774 582
<< pwell >>
rect 1 21 734 203
rect 30 -17 64 21
<< locali >>
rect 580 357 632 493
rect 18 215 115 255
rect 153 215 248 257
rect 204 135 248 215
rect 302 215 368 257
rect 402 215 483 255
rect 302 135 344 215
rect 598 117 632 357
rect 580 51 632 117
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 19 459 253 493
rect 19 325 85 459
rect 187 451 253 459
rect 291 443 362 527
rect 119 407 165 425
rect 396 407 446 493
rect 119 359 446 407
rect 480 375 546 527
rect 19 291 563 325
rect 19 17 109 170
rect 529 181 563 291
rect 395 147 563 181
rect 395 101 429 147
rect 666 289 700 527
rect 164 51 429 101
rect 471 17 537 113
rect 666 17 700 197
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
rlabel locali s 302 135 344 215 6 A1
port 1 nsew signal input
rlabel locali s 302 215 368 257 6 A1
port 1 nsew signal input
rlabel locali s 402 215 483 255 6 A2
port 2 nsew signal input
rlabel locali s 204 135 248 215 6 B1
port 3 nsew signal input
rlabel locali s 153 215 248 257 6 B1
port 3 nsew signal input
rlabel locali s 18 215 115 255 6 B2
port 4 nsew signal input
rlabel metal1 s 0 -48 736 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 1 21 734 203 6 VNB
port 6 nsew ground bidirectional
rlabel nwell s -38 261 774 582 6 VPB
port 7 nsew power bidirectional
rlabel metal1 s 0 496 736 592 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 580 51 632 117 6 X
port 9 nsew signal output
rlabel locali s 598 117 632 357 6 X
port 9 nsew signal output
rlabel locali s 580 357 632 493 6 X
port 9 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 736 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 4059210
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 4052462
<< end >>
