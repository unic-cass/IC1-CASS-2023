// This is the unpowered netlist.
module R4_butter (c1,
    c2,
    c3,
    Xio,
    Xro,
    la_oenb,
    xi0,
    xi1,
    xi2,
    xi3,
    xr0,
    xr1,
    xr2,
    xr3);
 input c1;
 input c2;
 input c3;
 output [3:0] Xio;
 output [3:0] Xro;
 output [7:0] la_oenb;
 input [3:0] xi0;
 input [3:0] xi1;
 input [3:0] xi2;
 input [3:0] xi3;
 input [3:0] xr0;
 input [3:0] xr1;
 input [3:0] xr2;
 input [3:0] xr3;

 wire net23;
 wire net24;
 wire net25;
 wire net20;
 wire net21;
 wire net22;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire _00_;
 wire _01_;
 wire _02_;
 wire _03_;
 wire _04_;
 wire _05_;
 wire net1;
 wire net10;
 wire net11;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;

 sky130_fd_sc_hd__decap_3 FILLER_0_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_93 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__conb_1 R4_butter_12 (.LO(net12));
 sky130_fd_sc_hd__conb_1 R4_butter_13 (.LO(net13));
 sky130_fd_sc_hd__conb_1 R4_butter_14 (.LO(net14));
 sky130_fd_sc_hd__conb_1 R4_butter_15 (.LO(net15));
 sky130_fd_sc_hd__conb_1 R4_butter_16 (.LO(net16));
 sky130_fd_sc_hd__conb_1 R4_butter_17 (.LO(net17));
 sky130_fd_sc_hd__conb_1 R4_butter_18 (.LO(net18));
 sky130_fd_sc_hd__conb_1 R4_butter_19 (.LO(net19));
 sky130_fd_sc_hd__conb_1 R4_butter_20 (.LO(net20));
 sky130_fd_sc_hd__conb_1 R4_butter_21 (.LO(net21));
 sky130_fd_sc_hd__conb_1 R4_butter_22 (.LO(net22));
 sky130_fd_sc_hd__conb_1 R4_butter_23 (.LO(net23));
 sky130_fd_sc_hd__conb_1 R4_butter_24 (.LO(net24));
 sky130_fd_sc_hd__conb_1 R4_butter_25 (.LO(net25));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__xnor2_1 _06_ (.A(net9),
    .B(net7),
    .Y(_00_));
 sky130_fd_sc_hd__xnor2_1 _07_ (.A(net8),
    .B(net6),
    .Y(_01_));
 sky130_fd_sc_hd__xnor2_1 _08_ (.A(net4),
    .B(net2),
    .Y(_02_));
 sky130_fd_sc_hd__mux2i_1 _09_ (.A0(_01_),
    .A1(_02_),
    .S(net1),
    .Y(_03_));
 sky130_fd_sc_hd__xnor2_1 _10_ (.A(_00_),
    .B(_03_),
    .Y(net11));
 sky130_fd_sc_hd__xnor2_1 _11_ (.A(net5),
    .B(net3),
    .Y(_04_));
 sky130_fd_sc_hd__mux2i_1 _12_ (.A0(_02_),
    .A1(_01_),
    .S(net1),
    .Y(_05_));
 sky130_fd_sc_hd__xnor2_1 _13_ (.A(_04_),
    .B(_05_),
    .Y(net10));
 sky130_fd_sc_hd__buf_2 input1 (.A(c1),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(xi0[0]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(xi1[0]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(xi2[0]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(xi3[0]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(xr0[0]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(xr1[0]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(xr2[0]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(xr3[0]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 output10 (.A(net10),
    .X(Xio[0]));
 sky130_fd_sc_hd__clkbuf_1 output11 (.A(net11),
    .X(Xro[0]));
 assign Xio[1] = net23;
 assign Xio[2] = net24;
 assign Xio[3] = net25;
 assign Xro[1] = net20;
 assign Xro[2] = net21;
 assign Xro[3] = net22;
 assign la_oenb[0] = net12;
 assign la_oenb[1] = net13;
 assign la_oenb[2] = net14;
 assign la_oenb[3] = net15;
 assign la_oenb[4] = net16;
 assign la_oenb[5] = net17;
 assign la_oenb[6] = net18;
 assign la_oenb[7] = net19;
endmodule

