magic
tech sky130B
magscale 1 2
timestamp 1676037725
<< locali >>
rect 185 1160 192 1194
rect 226 1160 264 1194
rect 298 1160 336 1194
rect 370 1160 408 1194
rect 442 1160 480 1194
rect 514 1160 552 1194
rect 586 1160 591 1194
rect 185 20 192 54
rect 226 20 264 54
rect 298 20 336 54
rect 370 20 408 54
rect 442 20 480 54
rect 514 20 552 54
rect 586 20 591 54
<< viali >>
rect 192 1160 226 1194
rect 264 1160 298 1194
rect 336 1160 370 1194
rect 408 1160 442 1194
rect 480 1160 514 1194
rect 552 1160 586 1194
rect 192 20 226 54
rect 264 20 298 54
rect 336 20 370 54
rect 408 20 442 54
rect 480 20 514 54
rect 552 20 586 54
<< obsli1 >>
rect 48 1020 82 1058
rect 48 948 82 986
rect 48 876 82 914
rect 48 804 82 842
rect 48 732 82 770
rect 48 660 82 698
rect 48 588 82 626
rect 48 516 82 554
rect 48 444 82 482
rect 48 372 82 410
rect 48 300 82 338
rect 48 228 82 266
rect 48 122 82 194
rect 159 98 193 1116
rect 265 98 299 1116
rect 371 98 405 1116
rect 477 98 511 1116
rect 583 98 617 1116
rect 694 1020 728 1058
rect 694 948 728 986
rect 694 876 728 914
rect 694 804 728 842
rect 694 732 728 770
rect 694 660 728 698
rect 694 588 728 626
rect 694 516 728 554
rect 694 444 728 482
rect 694 372 728 410
rect 694 300 728 338
rect 694 228 728 266
rect 694 122 728 194
<< obsli1c >>
rect 48 1058 82 1092
rect 48 986 82 1020
rect 48 914 82 948
rect 48 842 82 876
rect 48 770 82 804
rect 48 698 82 732
rect 48 626 82 660
rect 48 554 82 588
rect 48 482 82 516
rect 48 410 82 444
rect 48 338 82 372
rect 48 266 82 300
rect 48 194 82 228
rect 694 1058 728 1092
rect 694 986 728 1020
rect 694 914 728 948
rect 694 842 728 876
rect 694 770 728 804
rect 694 698 728 732
rect 694 626 728 660
rect 694 554 728 588
rect 694 482 728 516
rect 694 410 728 444
rect 694 338 728 372
rect 694 266 728 300
rect 694 194 728 228
<< metal1 >>
rect 180 1194 598 1214
rect 180 1160 192 1194
rect 226 1160 264 1194
rect 298 1160 336 1194
rect 370 1160 408 1194
rect 442 1160 480 1194
rect 514 1160 552 1194
rect 586 1160 598 1194
rect 180 1148 598 1160
rect 36 1092 94 1104
rect 36 1058 48 1092
rect 82 1058 94 1092
rect 36 1020 94 1058
rect 36 986 48 1020
rect 82 986 94 1020
rect 36 948 94 986
rect 36 914 48 948
rect 82 914 94 948
rect 36 876 94 914
rect 36 842 48 876
rect 82 842 94 876
rect 36 804 94 842
rect 36 770 48 804
rect 82 770 94 804
rect 36 732 94 770
rect 36 698 48 732
rect 82 698 94 732
rect 36 660 94 698
rect 36 626 48 660
rect 82 626 94 660
rect 36 588 94 626
rect 36 554 48 588
rect 82 554 94 588
rect 36 516 94 554
rect 36 482 48 516
rect 82 482 94 516
rect 36 444 94 482
rect 36 410 48 444
rect 82 410 94 444
rect 36 372 94 410
rect 36 338 48 372
rect 82 338 94 372
rect 36 300 94 338
rect 36 266 48 300
rect 82 266 94 300
rect 36 228 94 266
rect 36 194 48 228
rect 82 194 94 228
rect 36 110 94 194
rect 682 1092 740 1104
rect 682 1058 694 1092
rect 728 1058 740 1092
rect 682 1020 740 1058
rect 682 986 694 1020
rect 728 986 740 1020
rect 682 948 740 986
rect 682 914 694 948
rect 728 914 740 948
rect 682 876 740 914
rect 682 842 694 876
rect 728 842 740 876
rect 682 804 740 842
rect 682 770 694 804
rect 728 770 740 804
rect 682 732 740 770
rect 682 698 694 732
rect 728 698 740 732
rect 682 660 740 698
rect 682 626 694 660
rect 728 626 740 660
rect 682 588 740 626
rect 682 554 694 588
rect 728 554 740 588
rect 682 516 740 554
rect 682 482 694 516
rect 728 482 740 516
rect 682 444 740 482
rect 682 410 694 444
rect 728 410 740 444
rect 682 372 740 410
rect 682 338 694 372
rect 728 338 740 372
rect 682 300 740 338
rect 682 266 694 300
rect 728 266 740 300
rect 682 228 740 266
rect 682 194 694 228
rect 728 194 740 228
rect 682 110 740 194
rect 180 54 598 66
rect 180 20 192 54
rect 226 20 264 54
rect 298 20 336 54
rect 370 20 408 54
rect 442 20 480 54
rect 514 20 552 54
rect 586 20 598 54
rect 180 0 598 20
<< obsm1 >>
rect 150 110 202 1104
rect 256 110 308 1104
rect 362 110 414 1104
rect 468 110 520 1104
rect 574 110 626 1104
<< metal2 >>
rect 10 632 766 1104
rect 10 110 766 582
<< labels >>
rlabel metal1 s 682 110 740 1104 6 BULK
port 1 nsew
rlabel metal1 s 36 110 94 1104 6 BULK
port 1 nsew
rlabel metal2 s 10 632 766 1104 6 DRAIN
port 2 nsew
rlabel viali s 552 1160 586 1194 6 GATE
port 3 nsew
rlabel viali s 552 20 586 54 6 GATE
port 3 nsew
rlabel viali s 480 1160 514 1194 6 GATE
port 3 nsew
rlabel viali s 480 20 514 54 6 GATE
port 3 nsew
rlabel viali s 408 1160 442 1194 6 GATE
port 3 nsew
rlabel viali s 408 20 442 54 6 GATE
port 3 nsew
rlabel viali s 336 1160 370 1194 6 GATE
port 3 nsew
rlabel viali s 336 20 370 54 6 GATE
port 3 nsew
rlabel viali s 264 1160 298 1194 6 GATE
port 3 nsew
rlabel viali s 264 20 298 54 6 GATE
port 3 nsew
rlabel viali s 192 1160 226 1194 6 GATE
port 3 nsew
rlabel viali s 192 20 226 54 6 GATE
port 3 nsew
rlabel locali s 185 1160 591 1194 6 GATE
port 3 nsew
rlabel locali s 185 20 591 54 6 GATE
port 3 nsew
rlabel metal1 s 180 1148 598 1214 6 GATE
port 3 nsew
rlabel metal1 s 180 0 598 66 6 GATE
port 3 nsew
rlabel metal2 s 10 110 766 582 6 SOURCE
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 776 1214
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 9448112
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 9425826
<< end >>
