VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wb_buttons_leds
  CLASS BLOCK ;
  FOREIGN wb_buttons_leds ;
  ORIGIN 0.000 0.000 ;
  SIZE 434.190 BY 444.910 ;
  PIN buttons
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 430.190 9.560 434.190 10.160 ;
    END
  END buttons
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 12.050 440.910 12.330 444.910 ;
    END
  END clk
  PIN i_wb_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 36.890 440.910 37.170 444.910 ;
    END
  END i_wb_addr[0]
  PIN i_wb_addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 161.090 440.910 161.370 444.910 ;
    END
  END i_wb_addr[10]
  PIN i_wb_addr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 173.510 440.910 173.790 444.910 ;
    END
  END i_wb_addr[11]
  PIN i_wb_addr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 185.930 440.910 186.210 444.910 ;
    END
  END i_wb_addr[12]
  PIN i_wb_addr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 198.350 440.910 198.630 444.910 ;
    END
  END i_wb_addr[13]
  PIN i_wb_addr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 210.770 440.910 211.050 444.910 ;
    END
  END i_wb_addr[14]
  PIN i_wb_addr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 223.190 440.910 223.470 444.910 ;
    END
  END i_wb_addr[15]
  PIN i_wb_addr[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 235.610 440.910 235.890 444.910 ;
    END
  END i_wb_addr[16]
  PIN i_wb_addr[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 248.030 440.910 248.310 444.910 ;
    END
  END i_wb_addr[17]
  PIN i_wb_addr[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 260.450 440.910 260.730 444.910 ;
    END
  END i_wb_addr[18]
  PIN i_wb_addr[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 272.870 440.910 273.150 444.910 ;
    END
  END i_wb_addr[19]
  PIN i_wb_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 49.310 440.910 49.590 444.910 ;
    END
  END i_wb_addr[1]
  PIN i_wb_addr[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 285.290 440.910 285.570 444.910 ;
    END
  END i_wb_addr[20]
  PIN i_wb_addr[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 297.710 440.910 297.990 444.910 ;
    END
  END i_wb_addr[21]
  PIN i_wb_addr[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 310.130 440.910 310.410 444.910 ;
    END
  END i_wb_addr[22]
  PIN i_wb_addr[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 322.550 440.910 322.830 444.910 ;
    END
  END i_wb_addr[23]
  PIN i_wb_addr[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 334.970 440.910 335.250 444.910 ;
    END
  END i_wb_addr[24]
  PIN i_wb_addr[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 347.390 440.910 347.670 444.910 ;
    END
  END i_wb_addr[25]
  PIN i_wb_addr[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 359.810 440.910 360.090 444.910 ;
    END
  END i_wb_addr[26]
  PIN i_wb_addr[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 372.230 440.910 372.510 444.910 ;
    END
  END i_wb_addr[27]
  PIN i_wb_addr[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 384.650 440.910 384.930 444.910 ;
    END
  END i_wb_addr[28]
  PIN i_wb_addr[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 397.070 440.910 397.350 444.910 ;
    END
  END i_wb_addr[29]
  PIN i_wb_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 61.730 440.910 62.010 444.910 ;
    END
  END i_wb_addr[2]
  PIN i_wb_addr[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 409.490 440.910 409.770 444.910 ;
    END
  END i_wb_addr[30]
  PIN i_wb_addr[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 421.910 440.910 422.190 444.910 ;
    END
  END i_wb_addr[31]
  PIN i_wb_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 74.150 440.910 74.430 444.910 ;
    END
  END i_wb_addr[3]
  PIN i_wb_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 86.570 440.910 86.850 444.910 ;
    END
  END i_wb_addr[4]
  PIN i_wb_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 98.990 440.910 99.270 444.910 ;
    END
  END i_wb_addr[5]
  PIN i_wb_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 111.410 440.910 111.690 444.910 ;
    END
  END i_wb_addr[6]
  PIN i_wb_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 123.830 440.910 124.110 444.910 ;
    END
  END i_wb_addr[7]
  PIN i_wb_addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 136.250 440.910 136.530 444.910 ;
    END
  END i_wb_addr[8]
  PIN i_wb_addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 148.670 440.910 148.950 444.910 ;
    END
  END i_wb_addr[9]
  PIN i_wb_cyc
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 43.790 0.000 44.070 4.000 ;
    END
  END i_wb_cyc
  PIN i_wb_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END i_wb_data[0]
  PIN i_wb_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END i_wb_data[10]
  PIN i_wb_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END i_wb_data[11]
  PIN i_wb_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END i_wb_data[12]
  PIN i_wb_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END i_wb_data[13]
  PIN i_wb_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END i_wb_data[14]
  PIN i_wb_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END i_wb_data[15]
  PIN i_wb_data[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END i_wb_data[16]
  PIN i_wb_data[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 4.000 123.040 ;
    END
  END i_wb_data[17]
  PIN i_wb_data[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END i_wb_data[18]
  PIN i_wb_data[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 4.000 136.640 ;
    END
  END i_wb_data[19]
  PIN i_wb_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END i_wb_data[1]
  PIN i_wb_data[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END i_wb_data[20]
  PIN i_wb_data[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 4.000 150.240 ;
    END
  END i_wb_data[21]
  PIN i_wb_data[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END i_wb_data[22]
  PIN i_wb_data[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 4.000 163.840 ;
    END
  END i_wb_data[23]
  PIN i_wb_data[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 4.000 170.640 ;
    END
  END i_wb_data[24]
  PIN i_wb_data[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END i_wb_data[25]
  PIN i_wb_data[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 4.000 184.240 ;
    END
  END i_wb_data[26]
  PIN i_wb_data[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 190.440 4.000 191.040 ;
    END
  END i_wb_data[27]
  PIN i_wb_data[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.240 4.000 197.840 ;
    END
  END i_wb_data[28]
  PIN i_wb_data[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.040 4.000 204.640 ;
    END
  END i_wb_data[29]
  PIN i_wb_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END i_wb_data[2]
  PIN i_wb_data[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.840 4.000 211.440 ;
    END
  END i_wb_data[30]
  PIN i_wb_data[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 217.640 4.000 218.240 ;
    END
  END i_wb_data[31]
  PIN i_wb_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END i_wb_data[3]
  PIN i_wb_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END i_wb_data[4]
  PIN i_wb_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END i_wb_data[5]
  PIN i_wb_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END i_wb_data[6]
  PIN i_wb_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END i_wb_data[7]
  PIN i_wb_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END i_wb_data[8]
  PIN i_wb_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END i_wb_data[9]
  PIN i_wb_stb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 130.270 0.000 130.550 4.000 ;
    END
  END i_wb_stb
  PIN i_wb_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 216.750 0.000 217.030 4.000 ;
    END
  END i_wb_we
  PIN led_enb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 430.190 27.240 434.190 27.840 ;
    END
  END led_enb[0]
  PIN led_enb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 430.190 204.040 434.190 204.640 ;
    END
  END led_enb[10]
  PIN led_enb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 430.190 221.720 434.190 222.320 ;
    END
  END led_enb[11]
  PIN led_enb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 430.190 44.920 434.190 45.520 ;
    END
  END led_enb[1]
  PIN led_enb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 430.190 62.600 434.190 63.200 ;
    END
  END led_enb[2]
  PIN led_enb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 430.190 80.280 434.190 80.880 ;
    END
  END led_enb[3]
  PIN led_enb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 430.190 97.960 434.190 98.560 ;
    END
  END led_enb[4]
  PIN led_enb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 430.190 115.640 434.190 116.240 ;
    END
  END led_enb[5]
  PIN led_enb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 430.190 133.320 434.190 133.920 ;
    END
  END led_enb[6]
  PIN led_enb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 430.190 151.000 434.190 151.600 ;
    END
  END led_enb[7]
  PIN led_enb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 430.190 168.680 434.190 169.280 ;
    END
  END led_enb[8]
  PIN led_enb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 430.190 186.360 434.190 186.960 ;
    END
  END led_enb[9]
  PIN leds[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 430.190 239.400 434.190 240.000 ;
    END
  END leds[0]
  PIN leds[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 430.190 416.200 434.190 416.800 ;
    END
  END leds[10]
  PIN leds[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 430.190 433.880 434.190 434.480 ;
    END
  END leds[11]
  PIN leds[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 430.190 257.080 434.190 257.680 ;
    END
  END leds[1]
  PIN leds[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 430.190 274.760 434.190 275.360 ;
    END
  END leds[2]
  PIN leds[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 430.190 292.440 434.190 293.040 ;
    END
  END leds[3]
  PIN leds[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 430.190 310.120 434.190 310.720 ;
    END
  END leds[4]
  PIN leds[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 430.190 327.800 434.190 328.400 ;
    END
  END leds[5]
  PIN leds[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 430.190 345.480 434.190 346.080 ;
    END
  END leds[6]
  PIN leds[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 430.190 363.160 434.190 363.760 ;
    END
  END leds[7]
  PIN leds[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 430.190 380.840 434.190 381.440 ;
    END
  END leds[8]
  PIN leds[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 430.190 398.520 434.190 399.120 ;
    END
  END leds[9]
  PIN o_wb_ack
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 303.230 0.000 303.510 4.000 ;
    END
  END o_wb_ack
  PIN o_wb_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 224.440 4.000 225.040 ;
    END
  END o_wb_data[0]
  PIN o_wb_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 292.440 4.000 293.040 ;
    END
  END o_wb_data[10]
  PIN o_wb_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.240 4.000 299.840 ;
    END
  END o_wb_data[11]
  PIN o_wb_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 306.040 4.000 306.640 ;
    END
  END o_wb_data[12]
  PIN o_wb_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.840 4.000 313.440 ;
    END
  END o_wb_data[13]
  PIN o_wb_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 319.640 4.000 320.240 ;
    END
  END o_wb_data[14]
  PIN o_wb_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 326.440 4.000 327.040 ;
    END
  END o_wb_data[15]
  PIN o_wb_data[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 333.240 4.000 333.840 ;
    END
  END o_wb_data[16]
  PIN o_wb_data[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 340.040 4.000 340.640 ;
    END
  END o_wb_data[17]
  PIN o_wb_data[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.840 4.000 347.440 ;
    END
  END o_wb_data[18]
  PIN o_wb_data[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 353.640 4.000 354.240 ;
    END
  END o_wb_data[19]
  PIN o_wb_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.240 4.000 231.840 ;
    END
  END o_wb_data[1]
  PIN o_wb_data[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 360.440 4.000 361.040 ;
    END
  END o_wb_data[20]
  PIN o_wb_data[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 367.240 4.000 367.840 ;
    END
  END o_wb_data[21]
  PIN o_wb_data[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 374.040 4.000 374.640 ;
    END
  END o_wb_data[22]
  PIN o_wb_data[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 380.840 4.000 381.440 ;
    END
  END o_wb_data[23]
  PIN o_wb_data[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 387.640 4.000 388.240 ;
    END
  END o_wb_data[24]
  PIN o_wb_data[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 394.440 4.000 395.040 ;
    END
  END o_wb_data[25]
  PIN o_wb_data[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 401.240 4.000 401.840 ;
    END
  END o_wb_data[26]
  PIN o_wb_data[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 408.040 4.000 408.640 ;
    END
  END o_wb_data[27]
  PIN o_wb_data[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 414.840 4.000 415.440 ;
    END
  END o_wb_data[28]
  PIN o_wb_data[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 421.640 4.000 422.240 ;
    END
  END o_wb_data[29]
  PIN o_wb_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.040 4.000 238.640 ;
    END
  END o_wb_data[2]
  PIN o_wb_data[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 428.440 4.000 429.040 ;
    END
  END o_wb_data[30]
  PIN o_wb_data[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 435.240 4.000 435.840 ;
    END
  END o_wb_data[31]
  PIN o_wb_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.840 4.000 245.440 ;
    END
  END o_wb_data[3]
  PIN o_wb_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 251.640 4.000 252.240 ;
    END
  END o_wb_data[4]
  PIN o_wb_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 258.440 4.000 259.040 ;
    END
  END o_wb_data[5]
  PIN o_wb_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 265.240 4.000 265.840 ;
    END
  END o_wb_data[6]
  PIN o_wb_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.040 4.000 272.640 ;
    END
  END o_wb_data[7]
  PIN o_wb_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.840 4.000 279.440 ;
    END
  END o_wb_data[8]
  PIN o_wb_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 285.640 4.000 286.240 ;
    END
  END o_wb_data[9]
  PIN o_wb_stall
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.710 0.000 389.990 4.000 ;
    END
  END o_wb_stall
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 24.470 440.910 24.750 444.910 ;
    END
  END reset
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 11.720 10.640 13.320 432.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 165.320 10.640 166.920 432.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 318.920 10.640 320.520 432.720 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 88.520 10.640 90.120 432.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 242.120 10.640 243.720 432.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 395.720 10.640 397.320 432.720 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 428.260 432.565 ;
      LAYER met1 ;
        RECT 2.370 7.860 428.560 433.800 ;
      LAYER met2 ;
        RECT 2.400 440.630 11.770 441.050 ;
        RECT 12.610 440.630 24.190 441.050 ;
        RECT 25.030 440.630 36.610 441.050 ;
        RECT 37.450 440.630 49.030 441.050 ;
        RECT 49.870 440.630 61.450 441.050 ;
        RECT 62.290 440.630 73.870 441.050 ;
        RECT 74.710 440.630 86.290 441.050 ;
        RECT 87.130 440.630 98.710 441.050 ;
        RECT 99.550 440.630 111.130 441.050 ;
        RECT 111.970 440.630 123.550 441.050 ;
        RECT 124.390 440.630 135.970 441.050 ;
        RECT 136.810 440.630 148.390 441.050 ;
        RECT 149.230 440.630 160.810 441.050 ;
        RECT 161.650 440.630 173.230 441.050 ;
        RECT 174.070 440.630 185.650 441.050 ;
        RECT 186.490 440.630 198.070 441.050 ;
        RECT 198.910 440.630 210.490 441.050 ;
        RECT 211.330 440.630 222.910 441.050 ;
        RECT 223.750 440.630 235.330 441.050 ;
        RECT 236.170 440.630 247.750 441.050 ;
        RECT 248.590 440.630 260.170 441.050 ;
        RECT 261.010 440.630 272.590 441.050 ;
        RECT 273.430 440.630 285.010 441.050 ;
        RECT 285.850 440.630 297.430 441.050 ;
        RECT 298.270 440.630 309.850 441.050 ;
        RECT 310.690 440.630 322.270 441.050 ;
        RECT 323.110 440.630 334.690 441.050 ;
        RECT 335.530 440.630 347.110 441.050 ;
        RECT 347.950 440.630 359.530 441.050 ;
        RECT 360.370 440.630 371.950 441.050 ;
        RECT 372.790 440.630 384.370 441.050 ;
        RECT 385.210 440.630 396.790 441.050 ;
        RECT 397.630 440.630 409.210 441.050 ;
        RECT 410.050 440.630 421.630 441.050 ;
        RECT 422.470 440.630 427.710 441.050 ;
        RECT 2.400 4.280 427.710 440.630 ;
        RECT 2.400 3.670 43.510 4.280 ;
        RECT 44.350 3.670 129.990 4.280 ;
        RECT 130.830 3.670 216.470 4.280 ;
        RECT 217.310 3.670 302.950 4.280 ;
        RECT 303.790 3.670 389.430 4.280 ;
        RECT 390.270 3.670 427.710 4.280 ;
      LAYER met3 ;
        RECT 4.400 434.880 430.190 435.690 ;
        RECT 4.400 434.840 429.790 434.880 ;
        RECT 3.030 433.480 429.790 434.840 ;
        RECT 3.030 429.440 430.190 433.480 ;
        RECT 4.400 428.040 430.190 429.440 ;
        RECT 3.030 422.640 430.190 428.040 ;
        RECT 4.400 421.240 430.190 422.640 ;
        RECT 3.030 417.200 430.190 421.240 ;
        RECT 3.030 415.840 429.790 417.200 ;
        RECT 4.400 415.800 429.790 415.840 ;
        RECT 4.400 414.440 430.190 415.800 ;
        RECT 3.030 409.040 430.190 414.440 ;
        RECT 4.400 407.640 430.190 409.040 ;
        RECT 3.030 402.240 430.190 407.640 ;
        RECT 4.400 400.840 430.190 402.240 ;
        RECT 3.030 399.520 430.190 400.840 ;
        RECT 3.030 398.120 429.790 399.520 ;
        RECT 3.030 395.440 430.190 398.120 ;
        RECT 4.400 394.040 430.190 395.440 ;
        RECT 3.030 388.640 430.190 394.040 ;
        RECT 4.400 387.240 430.190 388.640 ;
        RECT 3.030 381.840 430.190 387.240 ;
        RECT 4.400 380.440 429.790 381.840 ;
        RECT 3.030 375.040 430.190 380.440 ;
        RECT 4.400 373.640 430.190 375.040 ;
        RECT 3.030 368.240 430.190 373.640 ;
        RECT 4.400 366.840 430.190 368.240 ;
        RECT 3.030 364.160 430.190 366.840 ;
        RECT 3.030 362.760 429.790 364.160 ;
        RECT 3.030 361.440 430.190 362.760 ;
        RECT 4.400 360.040 430.190 361.440 ;
        RECT 3.030 354.640 430.190 360.040 ;
        RECT 4.400 353.240 430.190 354.640 ;
        RECT 3.030 347.840 430.190 353.240 ;
        RECT 4.400 346.480 430.190 347.840 ;
        RECT 4.400 346.440 429.790 346.480 ;
        RECT 3.030 345.080 429.790 346.440 ;
        RECT 3.030 341.040 430.190 345.080 ;
        RECT 4.400 339.640 430.190 341.040 ;
        RECT 3.030 334.240 430.190 339.640 ;
        RECT 4.400 332.840 430.190 334.240 ;
        RECT 3.030 328.800 430.190 332.840 ;
        RECT 3.030 327.440 429.790 328.800 ;
        RECT 4.400 327.400 429.790 327.440 ;
        RECT 4.400 326.040 430.190 327.400 ;
        RECT 3.030 320.640 430.190 326.040 ;
        RECT 4.400 319.240 430.190 320.640 ;
        RECT 3.030 313.840 430.190 319.240 ;
        RECT 4.400 312.440 430.190 313.840 ;
        RECT 3.030 311.120 430.190 312.440 ;
        RECT 3.030 309.720 429.790 311.120 ;
        RECT 3.030 307.040 430.190 309.720 ;
        RECT 4.400 305.640 430.190 307.040 ;
        RECT 3.030 300.240 430.190 305.640 ;
        RECT 4.400 298.840 430.190 300.240 ;
        RECT 3.030 293.440 430.190 298.840 ;
        RECT 4.400 292.040 429.790 293.440 ;
        RECT 3.030 286.640 430.190 292.040 ;
        RECT 4.400 285.240 430.190 286.640 ;
        RECT 3.030 279.840 430.190 285.240 ;
        RECT 4.400 278.440 430.190 279.840 ;
        RECT 3.030 275.760 430.190 278.440 ;
        RECT 3.030 274.360 429.790 275.760 ;
        RECT 3.030 273.040 430.190 274.360 ;
        RECT 4.400 271.640 430.190 273.040 ;
        RECT 3.030 266.240 430.190 271.640 ;
        RECT 4.400 264.840 430.190 266.240 ;
        RECT 3.030 259.440 430.190 264.840 ;
        RECT 4.400 258.080 430.190 259.440 ;
        RECT 4.400 258.040 429.790 258.080 ;
        RECT 3.030 256.680 429.790 258.040 ;
        RECT 3.030 252.640 430.190 256.680 ;
        RECT 4.400 251.240 430.190 252.640 ;
        RECT 3.030 245.840 430.190 251.240 ;
        RECT 4.400 244.440 430.190 245.840 ;
        RECT 3.030 240.400 430.190 244.440 ;
        RECT 3.030 239.040 429.790 240.400 ;
        RECT 4.400 239.000 429.790 239.040 ;
        RECT 4.400 237.640 430.190 239.000 ;
        RECT 3.030 232.240 430.190 237.640 ;
        RECT 4.400 230.840 430.190 232.240 ;
        RECT 3.030 225.440 430.190 230.840 ;
        RECT 4.400 224.040 430.190 225.440 ;
        RECT 3.030 222.720 430.190 224.040 ;
        RECT 3.030 221.320 429.790 222.720 ;
        RECT 3.030 218.640 430.190 221.320 ;
        RECT 4.400 217.240 430.190 218.640 ;
        RECT 3.030 211.840 430.190 217.240 ;
        RECT 4.400 210.440 430.190 211.840 ;
        RECT 3.030 205.040 430.190 210.440 ;
        RECT 4.400 203.640 429.790 205.040 ;
        RECT 3.030 198.240 430.190 203.640 ;
        RECT 4.400 196.840 430.190 198.240 ;
        RECT 3.030 191.440 430.190 196.840 ;
        RECT 4.400 190.040 430.190 191.440 ;
        RECT 3.030 187.360 430.190 190.040 ;
        RECT 3.030 185.960 429.790 187.360 ;
        RECT 3.030 184.640 430.190 185.960 ;
        RECT 4.400 183.240 430.190 184.640 ;
        RECT 3.030 177.840 430.190 183.240 ;
        RECT 4.400 176.440 430.190 177.840 ;
        RECT 3.030 171.040 430.190 176.440 ;
        RECT 4.400 169.680 430.190 171.040 ;
        RECT 4.400 169.640 429.790 169.680 ;
        RECT 3.030 168.280 429.790 169.640 ;
        RECT 3.030 164.240 430.190 168.280 ;
        RECT 4.400 162.840 430.190 164.240 ;
        RECT 3.030 157.440 430.190 162.840 ;
        RECT 4.400 156.040 430.190 157.440 ;
        RECT 3.030 152.000 430.190 156.040 ;
        RECT 3.030 150.640 429.790 152.000 ;
        RECT 4.400 150.600 429.790 150.640 ;
        RECT 4.400 149.240 430.190 150.600 ;
        RECT 3.030 143.840 430.190 149.240 ;
        RECT 4.400 142.440 430.190 143.840 ;
        RECT 3.030 137.040 430.190 142.440 ;
        RECT 4.400 135.640 430.190 137.040 ;
        RECT 3.030 134.320 430.190 135.640 ;
        RECT 3.030 132.920 429.790 134.320 ;
        RECT 3.030 130.240 430.190 132.920 ;
        RECT 4.400 128.840 430.190 130.240 ;
        RECT 3.030 123.440 430.190 128.840 ;
        RECT 4.400 122.040 430.190 123.440 ;
        RECT 3.030 116.640 430.190 122.040 ;
        RECT 4.400 115.240 429.790 116.640 ;
        RECT 3.030 109.840 430.190 115.240 ;
        RECT 4.400 108.440 430.190 109.840 ;
        RECT 3.030 103.040 430.190 108.440 ;
        RECT 4.400 101.640 430.190 103.040 ;
        RECT 3.030 98.960 430.190 101.640 ;
        RECT 3.030 97.560 429.790 98.960 ;
        RECT 3.030 96.240 430.190 97.560 ;
        RECT 4.400 94.840 430.190 96.240 ;
        RECT 3.030 89.440 430.190 94.840 ;
        RECT 4.400 88.040 430.190 89.440 ;
        RECT 3.030 82.640 430.190 88.040 ;
        RECT 4.400 81.280 430.190 82.640 ;
        RECT 4.400 81.240 429.790 81.280 ;
        RECT 3.030 79.880 429.790 81.240 ;
        RECT 3.030 75.840 430.190 79.880 ;
        RECT 4.400 74.440 430.190 75.840 ;
        RECT 3.030 69.040 430.190 74.440 ;
        RECT 4.400 67.640 430.190 69.040 ;
        RECT 3.030 63.600 430.190 67.640 ;
        RECT 3.030 62.240 429.790 63.600 ;
        RECT 4.400 62.200 429.790 62.240 ;
        RECT 4.400 60.840 430.190 62.200 ;
        RECT 3.030 55.440 430.190 60.840 ;
        RECT 4.400 54.040 430.190 55.440 ;
        RECT 3.030 48.640 430.190 54.040 ;
        RECT 4.400 47.240 430.190 48.640 ;
        RECT 3.030 45.920 430.190 47.240 ;
        RECT 3.030 44.520 429.790 45.920 ;
        RECT 3.030 41.840 430.190 44.520 ;
        RECT 4.400 40.440 430.190 41.840 ;
        RECT 3.030 35.040 430.190 40.440 ;
        RECT 4.400 33.640 430.190 35.040 ;
        RECT 3.030 28.240 430.190 33.640 ;
        RECT 4.400 26.840 429.790 28.240 ;
        RECT 3.030 21.440 430.190 26.840 ;
        RECT 4.400 20.040 430.190 21.440 ;
        RECT 3.030 14.640 430.190 20.040 ;
        RECT 4.400 13.240 430.190 14.640 ;
        RECT 3.030 10.560 430.190 13.240 ;
        RECT 3.030 9.160 429.790 10.560 ;
        RECT 3.030 7.840 430.190 9.160 ;
        RECT 4.400 6.975 430.190 7.840 ;
      LAYER met4 ;
        RECT 2.630 10.240 11.320 428.905 ;
        RECT 13.720 10.240 88.120 428.905 ;
        RECT 90.520 10.240 164.920 428.905 ;
        RECT 167.320 10.240 241.720 428.905 ;
        RECT 244.120 10.240 318.520 428.905 ;
        RECT 320.920 10.240 395.320 428.905 ;
        RECT 397.720 10.240 415.050 428.905 ;
        RECT 2.630 9.695 415.050 10.240 ;
      LAYER met5 ;
        RECT 2.420 45.100 415.260 342.500 ;
  END
END wb_buttons_leds
END LIBRARY

