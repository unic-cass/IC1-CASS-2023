magic
tech sky130B
magscale 1 2
timestamp 1676037725
<< metal1 >>
rect 846 0 882 52140
rect 918 0 954 52140
rect 990 51429 1026 51770
rect 990 50639 1026 51271
rect 990 49849 1026 50481
rect 990 49059 1026 49691
rect 990 48269 1026 48901
rect 990 47479 1026 48111
rect 990 46689 1026 47321
rect 990 45899 1026 46531
rect 990 45109 1026 45741
rect 990 44319 1026 44951
rect 990 43529 1026 44161
rect 990 42739 1026 43371
rect 990 41949 1026 42581
rect 990 41159 1026 41791
rect 990 40369 1026 41001
rect 990 39579 1026 40211
rect 990 38789 1026 39421
rect 990 37999 1026 38631
rect 990 37209 1026 37841
rect 990 36419 1026 37051
rect 990 35629 1026 36261
rect 990 34839 1026 35471
rect 990 34049 1026 34681
rect 990 33259 1026 33891
rect 990 32469 1026 33101
rect 990 31679 1026 32311
rect 990 30889 1026 31521
rect 990 30099 1026 30731
rect 990 29309 1026 29941
rect 990 28519 1026 29151
rect 990 27729 1026 28361
rect 990 26939 1026 27571
rect 990 26149 1026 26781
rect 990 25359 1026 25991
rect 990 24569 1026 25201
rect 990 23779 1026 24411
rect 990 22989 1026 23621
rect 990 22199 1026 22831
rect 990 21409 1026 22041
rect 990 20619 1026 21251
rect 990 19829 1026 20461
rect 990 19039 1026 19671
rect 990 18249 1026 18881
rect 990 17459 1026 18091
rect 990 16669 1026 17301
rect 990 15879 1026 16511
rect 990 15089 1026 15721
rect 990 14299 1026 14931
rect 990 13509 1026 14141
rect 990 12719 1026 13351
rect 990 11929 1026 12561
rect 990 11139 1026 11771
rect 990 10349 1026 10981
rect 990 9559 1026 10191
rect 990 8769 1026 9401
rect 990 7979 1026 8611
rect 990 7189 1026 7821
rect 990 6399 1026 7031
rect 990 5609 1026 6241
rect 990 4819 1026 5451
rect 990 4029 1026 4661
rect 990 3239 1026 3871
rect 990 2449 1026 3081
rect 990 1659 1026 2291
rect 990 869 1026 1501
rect 990 370 1026 711
rect 1062 0 1098 52140
rect 1134 0 1170 52140
rect 1326 0 1362 52140
rect 1398 0 1434 52140
rect 1542 0 1578 52140
rect 1614 0 1650 52140
rect 2094 0 2130 52140
rect 2166 0 2202 52140
rect 2310 0 2346 52140
rect 2382 0 2418 52140
rect 2574 0 2610 52140
rect 2646 0 2682 52140
rect 2790 0 2826 52140
rect 2862 0 2898 52140
rect 3342 0 3378 52140
rect 3414 0 3450 52140
rect 3558 0 3594 52140
rect 3630 0 3666 52140
rect 3822 0 3858 52140
rect 3894 0 3930 52140
rect 4038 0 4074 52140
rect 4110 0 4146 52140
rect 4590 0 4626 52140
rect 4662 0 4698 52140
rect 4806 0 4842 52140
rect 4878 0 4914 52140
rect 5070 0 5106 52140
rect 5142 0 5178 52140
rect 5286 0 5322 52140
rect 5358 0 5394 52140
rect 5838 0 5874 52140
rect 5910 0 5946 52140
rect 6054 0 6090 52140
rect 6126 0 6162 52140
rect 6318 0 6354 52140
rect 6390 0 6426 52140
rect 6534 0 6570 52140
rect 6606 0 6642 52140
rect 7086 0 7122 52140
rect 7158 0 7194 52140
rect 7302 0 7338 52140
rect 7374 0 7410 52140
rect 7566 0 7602 52140
rect 7638 0 7674 52140
rect 7782 0 7818 52140
rect 7854 0 7890 52140
rect 8334 0 8370 52140
rect 8406 0 8442 52140
rect 8550 0 8586 52140
rect 8622 0 8658 52140
rect 8814 0 8850 52140
rect 8886 0 8922 52140
rect 9030 0 9066 52140
rect 9102 0 9138 52140
rect 9582 0 9618 52140
rect 9654 0 9690 52140
rect 9798 0 9834 52140
rect 9870 0 9906 52140
rect 10062 0 10098 52140
rect 10134 0 10170 52140
rect 10278 0 10314 52140
rect 10350 0 10386 52140
rect 10830 0 10866 52140
rect 10902 0 10938 52140
rect 11046 0 11082 52140
rect 11118 0 11154 52140
rect 11310 0 11346 52140
rect 11382 0 11418 52140
rect 11526 0 11562 52140
rect 11598 0 11634 52140
rect 12078 0 12114 52140
rect 12150 0 12186 52140
rect 12294 0 12330 52140
rect 12366 0 12402 52140
rect 12558 0 12594 52140
rect 12630 0 12666 52140
rect 12774 0 12810 52140
rect 12846 0 12882 52140
rect 13326 0 13362 52140
rect 13398 0 13434 52140
rect 13542 0 13578 52140
rect 13614 0 13650 52140
rect 13806 0 13842 52140
rect 13878 0 13914 52140
rect 14022 0 14058 52140
rect 14094 0 14130 52140
rect 14574 0 14610 52140
rect 14646 0 14682 52140
rect 14790 0 14826 52140
rect 14862 0 14898 52140
rect 15054 0 15090 52140
rect 15126 0 15162 52140
rect 15270 0 15306 52140
rect 15342 0 15378 52140
rect 15822 0 15858 52140
rect 15894 0 15930 52140
rect 16038 0 16074 52140
rect 16110 0 16146 52140
rect 16302 0 16338 52140
rect 16374 0 16410 52140
rect 16518 0 16554 52140
rect 16590 0 16626 52140
rect 17070 0 17106 52140
rect 17142 0 17178 52140
rect 17286 0 17322 52140
rect 17358 0 17394 52140
rect 17550 0 17586 52140
rect 17622 0 17658 52140
rect 17766 0 17802 52140
rect 17838 0 17874 52140
rect 18318 0 18354 52140
rect 18390 0 18426 52140
rect 18534 0 18570 52140
rect 18606 0 18642 52140
rect 18798 0 18834 52140
rect 18870 0 18906 52140
rect 19014 0 19050 52140
rect 19086 0 19122 52140
rect 19566 0 19602 52140
rect 19638 0 19674 52140
rect 19782 0 19818 52140
rect 19854 0 19890 52140
rect 20046 0 20082 52140
rect 20118 0 20154 52140
rect 20262 0 20298 52140
rect 20334 0 20370 52140
rect 20814 0 20850 52140
rect 20886 0 20922 52140
rect 21030 0 21066 52140
rect 21102 0 21138 52140
rect 21294 0 21330 52140
rect 21366 0 21402 52140
rect 21510 0 21546 52140
rect 21582 0 21618 52140
rect 22062 0 22098 52140
rect 22134 0 22170 52140
rect 22278 0 22314 52140
rect 22350 0 22386 52140
rect 22542 0 22578 52140
rect 22614 0 22650 52140
rect 22758 0 22794 52140
rect 22830 0 22866 52140
rect 23310 0 23346 52140
rect 23382 0 23418 52140
rect 23526 0 23562 52140
rect 23598 0 23634 52140
rect 23790 0 23826 52140
rect 23862 0 23898 52140
rect 24006 0 24042 52140
rect 24078 0 24114 52140
rect 24558 0 24594 52140
rect 24630 0 24666 52140
rect 24774 0 24810 52140
rect 24846 0 24882 52140
rect 25038 0 25074 52140
rect 25110 0 25146 52140
rect 25254 0 25290 52140
rect 25326 0 25362 52140
rect 25806 0 25842 52140
rect 25878 0 25914 52140
rect 26022 0 26058 52140
rect 26094 0 26130 52140
rect 26286 0 26322 52140
rect 26358 0 26394 52140
rect 26502 0 26538 52140
rect 26574 0 26610 52140
rect 27054 0 27090 52140
rect 27126 0 27162 52140
rect 27270 0 27306 52140
rect 27342 0 27378 52140
rect 27534 0 27570 52140
rect 27606 0 27642 52140
rect 27750 0 27786 52140
rect 27822 0 27858 52140
rect 28302 0 28338 52140
rect 28374 0 28410 52140
rect 28518 0 28554 52140
rect 28590 0 28626 52140
rect 28782 0 28818 52140
rect 28854 0 28890 52140
rect 28998 0 29034 52140
rect 29070 0 29106 52140
rect 29550 0 29586 52140
rect 29622 0 29658 52140
rect 29766 0 29802 52140
rect 29838 0 29874 52140
rect 30030 0 30066 52140
rect 30102 0 30138 52140
rect 30246 0 30282 52140
rect 30318 0 30354 52140
rect 30798 0 30834 52140
rect 30870 0 30906 52140
rect 31014 0 31050 52140
rect 31086 0 31122 52140
rect 31278 0 31314 52140
rect 31350 0 31386 52140
rect 31494 0 31530 52140
rect 31566 0 31602 52140
rect 32046 0 32082 52140
rect 32118 0 32154 52140
rect 32262 0 32298 52140
rect 32334 0 32370 52140
rect 32526 0 32562 52140
rect 32598 0 32634 52140
rect 32742 0 32778 52140
rect 32814 0 32850 52140
rect 33294 0 33330 52140
rect 33366 0 33402 52140
rect 33510 0 33546 52140
rect 33582 0 33618 52140
rect 33774 0 33810 52140
rect 33846 0 33882 52140
rect 33990 0 34026 52140
rect 34062 0 34098 52140
rect 34542 0 34578 52140
rect 34614 0 34650 52140
rect 34758 0 34794 52140
rect 34830 0 34866 52140
rect 35022 0 35058 52140
rect 35094 0 35130 52140
rect 35238 0 35274 52140
rect 35310 0 35346 52140
rect 35790 0 35826 52140
rect 35862 0 35898 52140
rect 36006 0 36042 52140
rect 36078 0 36114 52140
rect 36270 0 36306 52140
rect 36342 0 36378 52140
rect 36486 0 36522 52140
rect 36558 0 36594 52140
rect 37038 0 37074 52140
rect 37110 0 37146 52140
rect 37254 0 37290 52140
rect 37326 0 37362 52140
rect 37518 0 37554 52140
rect 37590 0 37626 52140
rect 37734 0 37770 52140
rect 37806 0 37842 52140
rect 38286 0 38322 52140
rect 38358 0 38394 52140
rect 38502 0 38538 52140
rect 38574 0 38610 52140
rect 38766 0 38802 52140
rect 38838 0 38874 52140
rect 38982 0 39018 52140
rect 39054 0 39090 52140
rect 39534 0 39570 52140
rect 39606 0 39642 52140
rect 39750 0 39786 52140
rect 39822 0 39858 52140
rect 40014 0 40050 52140
rect 40086 0 40122 52140
rect 40230 0 40266 52140
rect 40302 0 40338 52140
rect 40782 0 40818 52140
rect 40854 0 40890 52140
rect 40998 0 41034 52140
rect 41070 0 41106 52140
rect 41262 0 41298 52140
rect 41334 0 41370 52140
rect 41406 51429 41442 51770
rect 41406 50639 41442 51271
rect 41406 49849 41442 50481
rect 41406 49059 41442 49691
rect 41406 48269 41442 48901
rect 41406 47479 41442 48111
rect 41406 46689 41442 47321
rect 41406 45899 41442 46531
rect 41406 45109 41442 45741
rect 41406 44319 41442 44951
rect 41406 43529 41442 44161
rect 41406 42739 41442 43371
rect 41406 41949 41442 42581
rect 41406 41159 41442 41791
rect 41406 40369 41442 41001
rect 41406 39579 41442 40211
rect 41406 38789 41442 39421
rect 41406 37999 41442 38631
rect 41406 37209 41442 37841
rect 41406 36419 41442 37051
rect 41406 35629 41442 36261
rect 41406 34839 41442 35471
rect 41406 34049 41442 34681
rect 41406 33259 41442 33891
rect 41406 32469 41442 33101
rect 41406 31679 41442 32311
rect 41406 30889 41442 31521
rect 41406 30099 41442 30731
rect 41406 29309 41442 29941
rect 41406 28519 41442 29151
rect 41406 27729 41442 28361
rect 41406 26939 41442 27571
rect 41406 26149 41442 26781
rect 41406 25359 41442 25991
rect 41406 24569 41442 25201
rect 41406 23779 41442 24411
rect 41406 22989 41442 23621
rect 41406 22199 41442 22831
rect 41406 21409 41442 22041
rect 41406 20619 41442 21251
rect 41406 19829 41442 20461
rect 41406 19039 41442 19671
rect 41406 18249 41442 18881
rect 41406 17459 41442 18091
rect 41406 16669 41442 17301
rect 41406 15879 41442 16511
rect 41406 15089 41442 15721
rect 41406 14299 41442 14931
rect 41406 13509 41442 14141
rect 41406 12719 41442 13351
rect 41406 11929 41442 12561
rect 41406 11139 41442 11771
rect 41406 10349 41442 10981
rect 41406 9559 41442 10191
rect 41406 8769 41442 9401
rect 41406 7979 41442 8611
rect 41406 7189 41442 7821
rect 41406 6399 41442 7031
rect 41406 5609 41442 6241
rect 41406 4819 41442 5451
rect 41406 4029 41442 4661
rect 41406 3239 41442 3871
rect 41406 2449 41442 3081
rect 41406 1659 41442 2291
rect 41406 869 41442 1501
rect 41406 370 41442 711
rect 41478 0 41514 52140
rect 41550 0 41586 52140
<< metal2 >>
rect 954 51549 1062 51625
rect 41370 51549 41478 51625
rect 0 51453 42432 51501
rect 954 51295 1062 51405
rect 41370 51295 41478 51405
rect 0 51199 42432 51247
rect 954 51075 1062 51151
rect 41370 51075 41478 51151
rect 0 50979 42432 51027
rect 0 50883 42432 50931
rect 954 50759 1062 50835
rect 41370 50759 41478 50835
rect 0 50663 42432 50711
rect 954 50505 1062 50615
rect 41370 50505 41478 50615
rect 0 50409 42432 50457
rect 954 50285 1062 50361
rect 41370 50285 41478 50361
rect 0 50189 42432 50237
rect 0 50093 42432 50141
rect 954 49969 1062 50045
rect 41370 49969 41478 50045
rect 0 49873 42432 49921
rect 954 49715 1062 49825
rect 41370 49715 41478 49825
rect 0 49619 42432 49667
rect 954 49495 1062 49571
rect 41370 49495 41478 49571
rect 0 49399 42432 49447
rect 0 49303 42432 49351
rect 954 49179 1062 49255
rect 41370 49179 41478 49255
rect 0 49083 42432 49131
rect 954 48925 1062 49035
rect 41370 48925 41478 49035
rect 0 48829 42432 48877
rect 954 48705 1062 48781
rect 41370 48705 41478 48781
rect 0 48609 42432 48657
rect 0 48513 42432 48561
rect 954 48389 1062 48465
rect 41370 48389 41478 48465
rect 0 48293 42432 48341
rect 954 48135 1062 48245
rect 41370 48135 41478 48245
rect 0 48039 42432 48087
rect 954 47915 1062 47991
rect 41370 47915 41478 47991
rect 0 47819 42432 47867
rect 0 47723 42432 47771
rect 954 47599 1062 47675
rect 41370 47599 41478 47675
rect 0 47503 42432 47551
rect 954 47345 1062 47455
rect 41370 47345 41478 47455
rect 0 47249 42432 47297
rect 954 47125 1062 47201
rect 41370 47125 41478 47201
rect 0 47029 42432 47077
rect 0 46933 42432 46981
rect 954 46809 1062 46885
rect 41370 46809 41478 46885
rect 0 46713 42432 46761
rect 954 46555 1062 46665
rect 41370 46555 41478 46665
rect 0 46459 42432 46507
rect 954 46335 1062 46411
rect 41370 46335 41478 46411
rect 0 46239 42432 46287
rect 0 46143 42432 46191
rect 954 46019 1062 46095
rect 41370 46019 41478 46095
rect 0 45923 42432 45971
rect 954 45765 1062 45875
rect 41370 45765 41478 45875
rect 0 45669 42432 45717
rect 954 45545 1062 45621
rect 41370 45545 41478 45621
rect 0 45449 42432 45497
rect 0 45353 42432 45401
rect 954 45229 1062 45305
rect 41370 45229 41478 45305
rect 0 45133 42432 45181
rect 954 44975 1062 45085
rect 41370 44975 41478 45085
rect 0 44879 42432 44927
rect 954 44755 1062 44831
rect 41370 44755 41478 44831
rect 0 44659 42432 44707
rect 0 44563 42432 44611
rect 954 44439 1062 44515
rect 41370 44439 41478 44515
rect 0 44343 42432 44391
rect 954 44185 1062 44295
rect 41370 44185 41478 44295
rect 0 44089 42432 44137
rect 954 43965 1062 44041
rect 41370 43965 41478 44041
rect 0 43869 42432 43917
rect 0 43773 42432 43821
rect 954 43649 1062 43725
rect 41370 43649 41478 43725
rect 0 43553 42432 43601
rect 954 43395 1062 43505
rect 41370 43395 41478 43505
rect 0 43299 42432 43347
rect 954 43175 1062 43251
rect 41370 43175 41478 43251
rect 0 43079 42432 43127
rect 0 42983 42432 43031
rect 954 42859 1062 42935
rect 41370 42859 41478 42935
rect 0 42763 42432 42811
rect 954 42605 1062 42715
rect 41370 42605 41478 42715
rect 0 42509 42432 42557
rect 954 42385 1062 42461
rect 41370 42385 41478 42461
rect 0 42289 42432 42337
rect 0 42193 42432 42241
rect 954 42069 1062 42145
rect 41370 42069 41478 42145
rect 0 41973 42432 42021
rect 954 41815 1062 41925
rect 41370 41815 41478 41925
rect 0 41719 42432 41767
rect 954 41595 1062 41671
rect 41370 41595 41478 41671
rect 0 41499 42432 41547
rect 0 41403 42432 41451
rect 954 41279 1062 41355
rect 41370 41279 41478 41355
rect 0 41183 42432 41231
rect 954 41025 1062 41135
rect 41370 41025 41478 41135
rect 0 40929 42432 40977
rect 954 40805 1062 40881
rect 41370 40805 41478 40881
rect 0 40709 42432 40757
rect 0 40613 42432 40661
rect 954 40489 1062 40565
rect 41370 40489 41478 40565
rect 0 40393 42432 40441
rect 954 40235 1062 40345
rect 41370 40235 41478 40345
rect 0 40139 42432 40187
rect 954 40015 1062 40091
rect 41370 40015 41478 40091
rect 0 39919 42432 39967
rect 0 39823 42432 39871
rect 954 39699 1062 39775
rect 41370 39699 41478 39775
rect 0 39603 42432 39651
rect 954 39445 1062 39555
rect 41370 39445 41478 39555
rect 0 39349 42432 39397
rect 954 39225 1062 39301
rect 41370 39225 41478 39301
rect 0 39129 42432 39177
rect 0 39033 42432 39081
rect 954 38909 1062 38985
rect 41370 38909 41478 38985
rect 0 38813 42432 38861
rect 954 38655 1062 38765
rect 41370 38655 41478 38765
rect 0 38559 42432 38607
rect 954 38435 1062 38511
rect 41370 38435 41478 38511
rect 0 38339 42432 38387
rect 0 38243 42432 38291
rect 954 38119 1062 38195
rect 41370 38119 41478 38195
rect 0 38023 42432 38071
rect 954 37865 1062 37975
rect 41370 37865 41478 37975
rect 0 37769 42432 37817
rect 954 37645 1062 37721
rect 41370 37645 41478 37721
rect 0 37549 42432 37597
rect 0 37453 42432 37501
rect 954 37329 1062 37405
rect 41370 37329 41478 37405
rect 0 37233 42432 37281
rect 954 37075 1062 37185
rect 41370 37075 41478 37185
rect 0 36979 42432 37027
rect 954 36855 1062 36931
rect 41370 36855 41478 36931
rect 0 36759 42432 36807
rect 0 36663 42432 36711
rect 954 36539 1062 36615
rect 41370 36539 41478 36615
rect 0 36443 42432 36491
rect 954 36285 1062 36395
rect 41370 36285 41478 36395
rect 0 36189 42432 36237
rect 954 36065 1062 36141
rect 41370 36065 41478 36141
rect 0 35969 42432 36017
rect 0 35873 42432 35921
rect 954 35749 1062 35825
rect 41370 35749 41478 35825
rect 0 35653 42432 35701
rect 954 35495 1062 35605
rect 41370 35495 41478 35605
rect 0 35399 42432 35447
rect 954 35275 1062 35351
rect 41370 35275 41478 35351
rect 0 35179 42432 35227
rect 0 35083 42432 35131
rect 954 34959 1062 35035
rect 41370 34959 41478 35035
rect 0 34863 42432 34911
rect 954 34705 1062 34815
rect 41370 34705 41478 34815
rect 0 34609 42432 34657
rect 954 34485 1062 34561
rect 41370 34485 41478 34561
rect 0 34389 42432 34437
rect 0 34293 42432 34341
rect 954 34169 1062 34245
rect 41370 34169 41478 34245
rect 0 34073 42432 34121
rect 954 33915 1062 34025
rect 41370 33915 41478 34025
rect 0 33819 42432 33867
rect 954 33695 1062 33771
rect 41370 33695 41478 33771
rect 0 33599 42432 33647
rect 0 33503 42432 33551
rect 954 33379 1062 33455
rect 41370 33379 41478 33455
rect 0 33283 42432 33331
rect 954 33125 1062 33235
rect 41370 33125 41478 33235
rect 0 33029 42432 33077
rect 954 32905 1062 32981
rect 41370 32905 41478 32981
rect 0 32809 42432 32857
rect 0 32713 42432 32761
rect 954 32589 1062 32665
rect 41370 32589 41478 32665
rect 0 32493 42432 32541
rect 954 32335 1062 32445
rect 41370 32335 41478 32445
rect 0 32239 42432 32287
rect 954 32115 1062 32191
rect 41370 32115 41478 32191
rect 0 32019 42432 32067
rect 0 31923 42432 31971
rect 954 31799 1062 31875
rect 41370 31799 41478 31875
rect 0 31703 42432 31751
rect 954 31545 1062 31655
rect 41370 31545 41478 31655
rect 0 31449 42432 31497
rect 954 31325 1062 31401
rect 41370 31325 41478 31401
rect 0 31229 42432 31277
rect 0 31133 42432 31181
rect 954 31009 1062 31085
rect 41370 31009 41478 31085
rect 0 30913 42432 30961
rect 954 30755 1062 30865
rect 41370 30755 41478 30865
rect 0 30659 42432 30707
rect 954 30535 1062 30611
rect 41370 30535 41478 30611
rect 0 30439 42432 30487
rect 0 30343 42432 30391
rect 954 30219 1062 30295
rect 41370 30219 41478 30295
rect 0 30123 42432 30171
rect 954 29965 1062 30075
rect 41370 29965 41478 30075
rect 0 29869 42432 29917
rect 954 29745 1062 29821
rect 41370 29745 41478 29821
rect 0 29649 42432 29697
rect 0 29553 42432 29601
rect 954 29429 1062 29505
rect 41370 29429 41478 29505
rect 0 29333 42432 29381
rect 954 29175 1062 29285
rect 41370 29175 41478 29285
rect 0 29079 42432 29127
rect 954 28955 1062 29031
rect 41370 28955 41478 29031
rect 0 28859 42432 28907
rect 0 28763 42432 28811
rect 954 28639 1062 28715
rect 41370 28639 41478 28715
rect 0 28543 42432 28591
rect 954 28385 1062 28495
rect 41370 28385 41478 28495
rect 0 28289 42432 28337
rect 954 28165 1062 28241
rect 41370 28165 41478 28241
rect 0 28069 42432 28117
rect 0 27973 42432 28021
rect 954 27849 1062 27925
rect 41370 27849 41478 27925
rect 0 27753 42432 27801
rect 954 27595 1062 27705
rect 41370 27595 41478 27705
rect 0 27499 42432 27547
rect 954 27375 1062 27451
rect 41370 27375 41478 27451
rect 0 27279 42432 27327
rect 0 27183 42432 27231
rect 954 27059 1062 27135
rect 41370 27059 41478 27135
rect 0 26963 42432 27011
rect 954 26805 1062 26915
rect 41370 26805 41478 26915
rect 0 26709 42432 26757
rect 954 26585 1062 26661
rect 41370 26585 41478 26661
rect 0 26489 42432 26537
rect 0 26393 42432 26441
rect 954 26269 1062 26345
rect 41370 26269 41478 26345
rect 0 26173 42432 26221
rect 954 26015 1062 26125
rect 41370 26015 41478 26125
rect 0 25919 42432 25967
rect 954 25795 1062 25871
rect 41370 25795 41478 25871
rect 0 25699 42432 25747
rect 0 25603 42432 25651
rect 954 25479 1062 25555
rect 41370 25479 41478 25555
rect 0 25383 42432 25431
rect 954 25225 1062 25335
rect 41370 25225 41478 25335
rect 0 25129 42432 25177
rect 954 25005 1062 25081
rect 41370 25005 41478 25081
rect 0 24909 42432 24957
rect 0 24813 42432 24861
rect 954 24689 1062 24765
rect 41370 24689 41478 24765
rect 0 24593 42432 24641
rect 954 24435 1062 24545
rect 41370 24435 41478 24545
rect 0 24339 42432 24387
rect 954 24215 1062 24291
rect 41370 24215 41478 24291
rect 0 24119 42432 24167
rect 0 24023 42432 24071
rect 954 23899 1062 23975
rect 41370 23899 41478 23975
rect 0 23803 42432 23851
rect 954 23645 1062 23755
rect 41370 23645 41478 23755
rect 0 23549 42432 23597
rect 954 23425 1062 23501
rect 41370 23425 41478 23501
rect 0 23329 42432 23377
rect 0 23233 42432 23281
rect 954 23109 1062 23185
rect 41370 23109 41478 23185
rect 0 23013 42432 23061
rect 954 22855 1062 22965
rect 41370 22855 41478 22965
rect 0 22759 42432 22807
rect 954 22635 1062 22711
rect 41370 22635 41478 22711
rect 0 22539 42432 22587
rect 0 22443 42432 22491
rect 954 22319 1062 22395
rect 41370 22319 41478 22395
rect 0 22223 42432 22271
rect 954 22065 1062 22175
rect 41370 22065 41478 22175
rect 0 21969 42432 22017
rect 954 21845 1062 21921
rect 41370 21845 41478 21921
rect 0 21749 42432 21797
rect 0 21653 42432 21701
rect 954 21529 1062 21605
rect 41370 21529 41478 21605
rect 0 21433 42432 21481
rect 954 21275 1062 21385
rect 41370 21275 41478 21385
rect 0 21179 42432 21227
rect 954 21055 1062 21131
rect 41370 21055 41478 21131
rect 0 20959 42432 21007
rect 0 20863 42432 20911
rect 954 20739 1062 20815
rect 41370 20739 41478 20815
rect 0 20643 42432 20691
rect 954 20485 1062 20595
rect 41370 20485 41478 20595
rect 0 20389 42432 20437
rect 954 20265 1062 20341
rect 41370 20265 41478 20341
rect 0 20169 42432 20217
rect 0 20073 42432 20121
rect 954 19949 1062 20025
rect 41370 19949 41478 20025
rect 0 19853 42432 19901
rect 954 19695 1062 19805
rect 41370 19695 41478 19805
rect 0 19599 42432 19647
rect 954 19475 1062 19551
rect 41370 19475 41478 19551
rect 0 19379 42432 19427
rect 0 19283 42432 19331
rect 954 19159 1062 19235
rect 41370 19159 41478 19235
rect 0 19063 42432 19111
rect 954 18905 1062 19015
rect 41370 18905 41478 19015
rect 0 18809 42432 18857
rect 954 18685 1062 18761
rect 41370 18685 41478 18761
rect 0 18589 42432 18637
rect 0 18493 42432 18541
rect 954 18369 1062 18445
rect 41370 18369 41478 18445
rect 0 18273 42432 18321
rect 954 18115 1062 18225
rect 41370 18115 41478 18225
rect 0 18019 42432 18067
rect 954 17895 1062 17971
rect 41370 17895 41478 17971
rect 0 17799 42432 17847
rect 0 17703 42432 17751
rect 954 17579 1062 17655
rect 41370 17579 41478 17655
rect 0 17483 42432 17531
rect 954 17325 1062 17435
rect 41370 17325 41478 17435
rect 0 17229 42432 17277
rect 954 17105 1062 17181
rect 41370 17105 41478 17181
rect 0 17009 42432 17057
rect 0 16913 42432 16961
rect 954 16789 1062 16865
rect 41370 16789 41478 16865
rect 0 16693 42432 16741
rect 954 16535 1062 16645
rect 41370 16535 41478 16645
rect 0 16439 42432 16487
rect 954 16315 1062 16391
rect 41370 16315 41478 16391
rect 0 16219 42432 16267
rect 0 16123 42432 16171
rect 954 15999 1062 16075
rect 41370 15999 41478 16075
rect 0 15903 42432 15951
rect 954 15745 1062 15855
rect 41370 15745 41478 15855
rect 0 15649 42432 15697
rect 954 15525 1062 15601
rect 41370 15525 41478 15601
rect 0 15429 42432 15477
rect 0 15333 42432 15381
rect 954 15209 1062 15285
rect 41370 15209 41478 15285
rect 0 15113 42432 15161
rect 954 14955 1062 15065
rect 41370 14955 41478 15065
rect 0 14859 42432 14907
rect 954 14735 1062 14811
rect 41370 14735 41478 14811
rect 0 14639 42432 14687
rect 0 14543 42432 14591
rect 954 14419 1062 14495
rect 41370 14419 41478 14495
rect 0 14323 42432 14371
rect 954 14165 1062 14275
rect 41370 14165 41478 14275
rect 0 14069 42432 14117
rect 954 13945 1062 14021
rect 41370 13945 41478 14021
rect 0 13849 42432 13897
rect 0 13753 42432 13801
rect 954 13629 1062 13705
rect 41370 13629 41478 13705
rect 0 13533 42432 13581
rect 954 13375 1062 13485
rect 41370 13375 41478 13485
rect 0 13279 42432 13327
rect 954 13155 1062 13231
rect 41370 13155 41478 13231
rect 0 13059 42432 13107
rect 0 12963 42432 13011
rect 954 12839 1062 12915
rect 41370 12839 41478 12915
rect 0 12743 42432 12791
rect 954 12585 1062 12695
rect 41370 12585 41478 12695
rect 0 12489 42432 12537
rect 954 12365 1062 12441
rect 41370 12365 41478 12441
rect 0 12269 42432 12317
rect 0 12173 42432 12221
rect 954 12049 1062 12125
rect 41370 12049 41478 12125
rect 0 11953 42432 12001
rect 954 11795 1062 11905
rect 41370 11795 41478 11905
rect 0 11699 42432 11747
rect 954 11575 1062 11651
rect 41370 11575 41478 11651
rect 0 11479 42432 11527
rect 0 11383 42432 11431
rect 954 11259 1062 11335
rect 41370 11259 41478 11335
rect 0 11163 42432 11211
rect 954 11005 1062 11115
rect 41370 11005 41478 11115
rect 0 10909 42432 10957
rect 954 10785 1062 10861
rect 41370 10785 41478 10861
rect 0 10689 42432 10737
rect 0 10593 42432 10641
rect 954 10469 1062 10545
rect 41370 10469 41478 10545
rect 0 10373 42432 10421
rect 954 10215 1062 10325
rect 41370 10215 41478 10325
rect 0 10119 42432 10167
rect 954 9995 1062 10071
rect 41370 9995 41478 10071
rect 0 9899 42432 9947
rect 0 9803 42432 9851
rect 954 9679 1062 9755
rect 41370 9679 41478 9755
rect 0 9583 42432 9631
rect 954 9425 1062 9535
rect 41370 9425 41478 9535
rect 0 9329 42432 9377
rect 954 9205 1062 9281
rect 41370 9205 41478 9281
rect 0 9109 42432 9157
rect 0 9013 42432 9061
rect 954 8889 1062 8965
rect 41370 8889 41478 8965
rect 0 8793 42432 8841
rect 954 8635 1062 8745
rect 41370 8635 41478 8745
rect 0 8539 42432 8587
rect 954 8415 1062 8491
rect 41370 8415 41478 8491
rect 0 8319 42432 8367
rect 0 8223 42432 8271
rect 954 8099 1062 8175
rect 41370 8099 41478 8175
rect 0 8003 42432 8051
rect 954 7845 1062 7955
rect 41370 7845 41478 7955
rect 0 7749 42432 7797
rect 954 7625 1062 7701
rect 41370 7625 41478 7701
rect 0 7529 42432 7577
rect 0 7433 42432 7481
rect 954 7309 1062 7385
rect 41370 7309 41478 7385
rect 0 7213 42432 7261
rect 954 7055 1062 7165
rect 41370 7055 41478 7165
rect 0 6959 42432 7007
rect 954 6835 1062 6911
rect 41370 6835 41478 6911
rect 0 6739 42432 6787
rect 0 6643 42432 6691
rect 954 6519 1062 6595
rect 41370 6519 41478 6595
rect 0 6423 42432 6471
rect 954 6265 1062 6375
rect 41370 6265 41478 6375
rect 0 6169 42432 6217
rect 954 6045 1062 6121
rect 41370 6045 41478 6121
rect 0 5949 42432 5997
rect 0 5853 42432 5901
rect 954 5729 1062 5805
rect 41370 5729 41478 5805
rect 0 5633 42432 5681
rect 954 5475 1062 5585
rect 41370 5475 41478 5585
rect 0 5379 42432 5427
rect 954 5255 1062 5331
rect 41370 5255 41478 5331
rect 0 5159 42432 5207
rect 0 5063 42432 5111
rect 954 4939 1062 5015
rect 41370 4939 41478 5015
rect 0 4843 42432 4891
rect 954 4685 1062 4795
rect 41370 4685 41478 4795
rect 0 4589 42432 4637
rect 954 4465 1062 4541
rect 41370 4465 41478 4541
rect 0 4369 42432 4417
rect 0 4273 42432 4321
rect 954 4149 1062 4225
rect 41370 4149 41478 4225
rect 0 4053 42432 4101
rect 954 3895 1062 4005
rect 41370 3895 41478 4005
rect 0 3799 42432 3847
rect 954 3675 1062 3751
rect 41370 3675 41478 3751
rect 0 3579 42432 3627
rect 0 3483 42432 3531
rect 954 3359 1062 3435
rect 41370 3359 41478 3435
rect 0 3263 42432 3311
rect 954 3105 1062 3215
rect 41370 3105 41478 3215
rect 0 3009 42432 3057
rect 954 2885 1062 2961
rect 41370 2885 41478 2961
rect 0 2789 42432 2837
rect 0 2693 42432 2741
rect 954 2569 1062 2645
rect 41370 2569 41478 2645
rect 0 2473 42432 2521
rect 954 2315 1062 2425
rect 41370 2315 41478 2425
rect 0 2219 42432 2267
rect 954 2095 1062 2171
rect 41370 2095 41478 2171
rect 0 1999 42432 2047
rect 0 1903 42432 1951
rect 954 1779 1062 1855
rect 41370 1779 41478 1855
rect 0 1683 42432 1731
rect 954 1525 1062 1635
rect 41370 1525 41478 1635
rect 0 1429 42432 1477
rect 954 1305 1062 1381
rect 41370 1305 41478 1381
rect 0 1209 42432 1257
rect 0 1113 42432 1161
rect 954 989 1062 1065
rect 41370 989 41478 1065
rect 0 893 42432 941
rect 954 735 1062 845
rect 41370 735 41478 845
rect 954 515 1062 591
rect 41370 515 41478 591
rect 0 419 42432 467
<< metal3 >>
rect 887 51862 985 51960
rect 1530 51881 1590 51941
rect 2154 51881 2214 51941
rect 2778 51881 2838 51941
rect 3402 51881 3462 51941
rect 4026 51881 4086 51941
rect 4650 51881 4710 51941
rect 5274 51881 5334 51941
rect 5898 51881 5958 51941
rect 6522 51881 6582 51941
rect 7146 51881 7206 51941
rect 7770 51881 7830 51941
rect 8394 51881 8454 51941
rect 9018 51881 9078 51941
rect 9642 51881 9702 51941
rect 10266 51881 10326 51941
rect 10890 51881 10950 51941
rect 11514 51881 11574 51941
rect 12138 51881 12198 51941
rect 12762 51881 12822 51941
rect 13386 51881 13446 51941
rect 14010 51881 14070 51941
rect 14634 51881 14694 51941
rect 15258 51881 15318 51941
rect 15882 51881 15942 51941
rect 16506 51881 16566 51941
rect 17130 51881 17190 51941
rect 17754 51881 17814 51941
rect 18378 51881 18438 51941
rect 19002 51881 19062 51941
rect 19626 51881 19686 51941
rect 20250 51881 20310 51941
rect 20874 51881 20934 51941
rect 21498 51881 21558 51941
rect 22122 51881 22182 51941
rect 22746 51881 22806 51941
rect 23370 51881 23430 51941
rect 23994 51881 24054 51941
rect 24618 51881 24678 51941
rect 25242 51881 25302 51941
rect 25866 51881 25926 51941
rect 26490 51881 26550 51941
rect 27114 51881 27174 51941
rect 27738 51881 27798 51941
rect 28362 51881 28422 51941
rect 28986 51881 29046 51941
rect 29610 51881 29670 51941
rect 30234 51881 30294 51941
rect 30858 51881 30918 51941
rect 31482 51881 31542 51941
rect 32106 51881 32166 51941
rect 32730 51881 32790 51941
rect 33354 51881 33414 51941
rect 33978 51881 34038 51941
rect 34602 51881 34662 51941
rect 35226 51881 35286 51941
rect 35850 51881 35910 51941
rect 36474 51881 36534 51941
rect 37098 51881 37158 51941
rect 37722 51881 37782 51941
rect 38346 51881 38406 51941
rect 38970 51881 39030 51941
rect 39594 51881 39654 51941
rect 40218 51881 40278 51941
rect 40842 51881 40902 51941
rect 41447 51862 41545 51960
rect 210 51557 270 51617
rect 42162 51557 42222 51617
rect 210 51320 270 51380
rect 42162 51320 42222 51380
rect 210 51083 270 51143
rect 42162 51083 42222 51143
rect 210 50767 270 50827
rect 42162 50767 42222 50827
rect 210 50530 270 50590
rect 42162 50530 42222 50590
rect 210 50293 270 50353
rect 42162 50293 42222 50353
rect 210 49977 270 50037
rect 42162 49977 42222 50037
rect 210 49740 270 49800
rect 42162 49740 42222 49800
rect 210 49503 270 49563
rect 42162 49503 42222 49563
rect 210 49187 270 49247
rect 42162 49187 42222 49247
rect 210 48950 270 49010
rect 42162 48950 42222 49010
rect 210 48713 270 48773
rect 42162 48713 42222 48773
rect 210 48397 270 48457
rect 42162 48397 42222 48457
rect 210 48160 270 48220
rect 42162 48160 42222 48220
rect 210 47923 270 47983
rect 42162 47923 42222 47983
rect 210 47607 270 47667
rect 42162 47607 42222 47667
rect 210 47370 270 47430
rect 42162 47370 42222 47430
rect 210 47133 270 47193
rect 42162 47133 42222 47193
rect 210 46817 270 46877
rect 42162 46817 42222 46877
rect 210 46580 270 46640
rect 42162 46580 42222 46640
rect 210 46343 270 46403
rect 42162 46343 42222 46403
rect 210 46027 270 46087
rect 42162 46027 42222 46087
rect 210 45790 270 45850
rect 42162 45790 42222 45850
rect 210 45553 270 45613
rect 42162 45553 42222 45613
rect 210 45237 270 45297
rect 42162 45237 42222 45297
rect 210 45000 270 45060
rect 42162 45000 42222 45060
rect 210 44763 270 44823
rect 42162 44763 42222 44823
rect 210 44447 270 44507
rect 42162 44447 42222 44507
rect 210 44210 270 44270
rect 42162 44210 42222 44270
rect 210 43973 270 44033
rect 42162 43973 42222 44033
rect 210 43657 270 43717
rect 42162 43657 42222 43717
rect 210 43420 270 43480
rect 42162 43420 42222 43480
rect 210 43183 270 43243
rect 42162 43183 42222 43243
rect 210 42867 270 42927
rect 42162 42867 42222 42927
rect 210 42630 270 42690
rect 42162 42630 42222 42690
rect 210 42393 270 42453
rect 42162 42393 42222 42453
rect 210 42077 270 42137
rect 42162 42077 42222 42137
rect 210 41840 270 41900
rect 42162 41840 42222 41900
rect 210 41603 270 41663
rect 42162 41603 42222 41663
rect 210 41287 270 41347
rect 42162 41287 42222 41347
rect 210 41050 270 41110
rect 42162 41050 42222 41110
rect 210 40813 270 40873
rect 42162 40813 42222 40873
rect 210 40497 270 40557
rect 42162 40497 42222 40557
rect 210 40260 270 40320
rect 42162 40260 42222 40320
rect 210 40023 270 40083
rect 42162 40023 42222 40083
rect 210 39707 270 39767
rect 42162 39707 42222 39767
rect 210 39470 270 39530
rect 42162 39470 42222 39530
rect 210 39233 270 39293
rect 42162 39233 42222 39293
rect 210 38917 270 38977
rect 42162 38917 42222 38977
rect 210 38680 270 38740
rect 42162 38680 42222 38740
rect 210 38443 270 38503
rect 42162 38443 42222 38503
rect 210 38127 270 38187
rect 42162 38127 42222 38187
rect 210 37890 270 37950
rect 42162 37890 42222 37950
rect 210 37653 270 37713
rect 42162 37653 42222 37713
rect 210 37337 270 37397
rect 42162 37337 42222 37397
rect 210 37100 270 37160
rect 42162 37100 42222 37160
rect 210 36863 270 36923
rect 42162 36863 42222 36923
rect 210 36547 270 36607
rect 42162 36547 42222 36607
rect 210 36310 270 36370
rect 42162 36310 42222 36370
rect 210 36073 270 36133
rect 42162 36073 42222 36133
rect 210 35757 270 35817
rect 42162 35757 42222 35817
rect 210 35520 270 35580
rect 42162 35520 42222 35580
rect 210 35283 270 35343
rect 42162 35283 42222 35343
rect 210 34967 270 35027
rect 42162 34967 42222 35027
rect 210 34730 270 34790
rect 42162 34730 42222 34790
rect 210 34493 270 34553
rect 42162 34493 42222 34553
rect 210 34177 270 34237
rect 42162 34177 42222 34237
rect 210 33940 270 34000
rect 42162 33940 42222 34000
rect 210 33703 270 33763
rect 42162 33703 42222 33763
rect 210 33387 270 33447
rect 42162 33387 42222 33447
rect 210 33150 270 33210
rect 42162 33150 42222 33210
rect 210 32913 270 32973
rect 42162 32913 42222 32973
rect 210 32597 270 32657
rect 42162 32597 42222 32657
rect 210 32360 270 32420
rect 42162 32360 42222 32420
rect 210 32123 270 32183
rect 42162 32123 42222 32183
rect 210 31807 270 31867
rect 42162 31807 42222 31867
rect 210 31570 270 31630
rect 42162 31570 42222 31630
rect 210 31333 270 31393
rect 42162 31333 42222 31393
rect 210 31017 270 31077
rect 42162 31017 42222 31077
rect 210 30780 270 30840
rect 42162 30780 42222 30840
rect 210 30543 270 30603
rect 42162 30543 42222 30603
rect 210 30227 270 30287
rect 42162 30227 42222 30287
rect 210 29990 270 30050
rect 42162 29990 42222 30050
rect 210 29753 270 29813
rect 42162 29753 42222 29813
rect 210 29437 270 29497
rect 42162 29437 42222 29497
rect 210 29200 270 29260
rect 42162 29200 42222 29260
rect 210 28963 270 29023
rect 42162 28963 42222 29023
rect 210 28647 270 28707
rect 42162 28647 42222 28707
rect 210 28410 270 28470
rect 42162 28410 42222 28470
rect 210 28173 270 28233
rect 42162 28173 42222 28233
rect 210 27857 270 27917
rect 42162 27857 42222 27917
rect 210 27620 270 27680
rect 42162 27620 42222 27680
rect 210 27383 270 27443
rect 42162 27383 42222 27443
rect 210 27067 270 27127
rect 42162 27067 42222 27127
rect 210 26830 270 26890
rect 42162 26830 42222 26890
rect 210 26593 270 26653
rect 42162 26593 42222 26653
rect 210 26277 270 26337
rect 42162 26277 42222 26337
rect 210 26040 270 26100
rect 42162 26040 42222 26100
rect 210 25803 270 25863
rect 42162 25803 42222 25863
rect 210 25487 270 25547
rect 42162 25487 42222 25547
rect 210 25250 270 25310
rect 42162 25250 42222 25310
rect 210 25013 270 25073
rect 42162 25013 42222 25073
rect 210 24697 270 24757
rect 42162 24697 42222 24757
rect 210 24460 270 24520
rect 42162 24460 42222 24520
rect 210 24223 270 24283
rect 42162 24223 42222 24283
rect 210 23907 270 23967
rect 42162 23907 42222 23967
rect 210 23670 270 23730
rect 42162 23670 42222 23730
rect 210 23433 270 23493
rect 42162 23433 42222 23493
rect 210 23117 270 23177
rect 42162 23117 42222 23177
rect 210 22880 270 22940
rect 42162 22880 42222 22940
rect 210 22643 270 22703
rect 42162 22643 42222 22703
rect 210 22327 270 22387
rect 42162 22327 42222 22387
rect 210 22090 270 22150
rect 42162 22090 42222 22150
rect 210 21853 270 21913
rect 42162 21853 42222 21913
rect 210 21537 270 21597
rect 42162 21537 42222 21597
rect 210 21300 270 21360
rect 42162 21300 42222 21360
rect 210 21063 270 21123
rect 42162 21063 42222 21123
rect 210 20747 270 20807
rect 42162 20747 42222 20807
rect 210 20510 270 20570
rect 42162 20510 42222 20570
rect 210 20273 270 20333
rect 42162 20273 42222 20333
rect 210 19957 270 20017
rect 42162 19957 42222 20017
rect 210 19720 270 19780
rect 42162 19720 42222 19780
rect 210 19483 270 19543
rect 42162 19483 42222 19543
rect 210 19167 270 19227
rect 42162 19167 42222 19227
rect 210 18930 270 18990
rect 42162 18930 42222 18990
rect 210 18693 270 18753
rect 42162 18693 42222 18753
rect 210 18377 270 18437
rect 42162 18377 42222 18437
rect 210 18140 270 18200
rect 42162 18140 42222 18200
rect 210 17903 270 17963
rect 42162 17903 42222 17963
rect 210 17587 270 17647
rect 42162 17587 42222 17647
rect 210 17350 270 17410
rect 42162 17350 42222 17410
rect 210 17113 270 17173
rect 42162 17113 42222 17173
rect 210 16797 270 16857
rect 42162 16797 42222 16857
rect 210 16560 270 16620
rect 42162 16560 42222 16620
rect 210 16323 270 16383
rect 42162 16323 42222 16383
rect 210 16007 270 16067
rect 42162 16007 42222 16067
rect 210 15770 270 15830
rect 42162 15770 42222 15830
rect 210 15533 270 15593
rect 42162 15533 42222 15593
rect 210 15217 270 15277
rect 42162 15217 42222 15277
rect 210 14980 270 15040
rect 42162 14980 42222 15040
rect 210 14743 270 14803
rect 42162 14743 42222 14803
rect 210 14427 270 14487
rect 42162 14427 42222 14487
rect 210 14190 270 14250
rect 42162 14190 42222 14250
rect 210 13953 270 14013
rect 42162 13953 42222 14013
rect 210 13637 270 13697
rect 42162 13637 42222 13697
rect 210 13400 270 13460
rect 42162 13400 42222 13460
rect 210 13163 270 13223
rect 42162 13163 42222 13223
rect 210 12847 270 12907
rect 42162 12847 42222 12907
rect 210 12610 270 12670
rect 42162 12610 42222 12670
rect 210 12373 270 12433
rect 42162 12373 42222 12433
rect 210 12057 270 12117
rect 42162 12057 42222 12117
rect 210 11820 270 11880
rect 42162 11820 42222 11880
rect 210 11583 270 11643
rect 42162 11583 42222 11643
rect 210 11267 270 11327
rect 42162 11267 42222 11327
rect 210 11030 270 11090
rect 42162 11030 42222 11090
rect 210 10793 270 10853
rect 42162 10793 42222 10853
rect 210 10477 270 10537
rect 42162 10477 42222 10537
rect 210 10240 270 10300
rect 42162 10240 42222 10300
rect 210 10003 270 10063
rect 42162 10003 42222 10063
rect 210 9687 270 9747
rect 42162 9687 42222 9747
rect 210 9450 270 9510
rect 42162 9450 42222 9510
rect 210 9213 270 9273
rect 42162 9213 42222 9273
rect 210 8897 270 8957
rect 42162 8897 42222 8957
rect 210 8660 270 8720
rect 42162 8660 42222 8720
rect 210 8423 270 8483
rect 42162 8423 42222 8483
rect 210 8107 270 8167
rect 42162 8107 42222 8167
rect 210 7870 270 7930
rect 42162 7870 42222 7930
rect 210 7633 270 7693
rect 42162 7633 42222 7693
rect 210 7317 270 7377
rect 42162 7317 42222 7377
rect 210 7080 270 7140
rect 42162 7080 42222 7140
rect 210 6843 270 6903
rect 42162 6843 42222 6903
rect 210 6527 270 6587
rect 42162 6527 42222 6587
rect 210 6290 270 6350
rect 42162 6290 42222 6350
rect 210 6053 270 6113
rect 42162 6053 42222 6113
rect 210 5737 270 5797
rect 42162 5737 42222 5797
rect 210 5500 270 5560
rect 42162 5500 42222 5560
rect 210 5263 270 5323
rect 42162 5263 42222 5323
rect 210 4947 270 5007
rect 42162 4947 42222 5007
rect 210 4710 270 4770
rect 42162 4710 42222 4770
rect 210 4473 270 4533
rect 42162 4473 42222 4533
rect 210 4157 270 4217
rect 42162 4157 42222 4217
rect 210 3920 270 3980
rect 42162 3920 42222 3980
rect 210 3683 270 3743
rect 42162 3683 42222 3743
rect 210 3367 270 3427
rect 42162 3367 42222 3427
rect 210 3130 270 3190
rect 42162 3130 42222 3190
rect 210 2893 270 2953
rect 42162 2893 42222 2953
rect 210 2577 270 2637
rect 42162 2577 42222 2637
rect 210 2340 270 2400
rect 42162 2340 42222 2400
rect 210 2103 270 2163
rect 42162 2103 42222 2163
rect 210 1787 270 1847
rect 42162 1787 42222 1847
rect 210 1550 270 1610
rect 42162 1550 42222 1610
rect 210 1313 270 1373
rect 42162 1313 42222 1373
rect 210 997 270 1057
rect 42162 997 42222 1057
rect 210 760 270 820
rect 42162 760 42222 820
rect 210 523 270 583
rect 42162 523 42222 583
rect 887 180 985 278
rect 1530 199 1590 259
rect 2154 199 2214 259
rect 2778 199 2838 259
rect 3402 199 3462 259
rect 4026 199 4086 259
rect 4650 199 4710 259
rect 5274 199 5334 259
rect 5898 199 5958 259
rect 6522 199 6582 259
rect 7146 199 7206 259
rect 7770 199 7830 259
rect 8394 199 8454 259
rect 9018 199 9078 259
rect 9642 199 9702 259
rect 10266 199 10326 259
rect 10890 199 10950 259
rect 11514 199 11574 259
rect 12138 199 12198 259
rect 12762 199 12822 259
rect 13386 199 13446 259
rect 14010 199 14070 259
rect 14634 199 14694 259
rect 15258 199 15318 259
rect 15882 199 15942 259
rect 16506 199 16566 259
rect 17130 199 17190 259
rect 17754 199 17814 259
rect 18378 199 18438 259
rect 19002 199 19062 259
rect 19626 199 19686 259
rect 20250 199 20310 259
rect 20874 199 20934 259
rect 21498 199 21558 259
rect 22122 199 22182 259
rect 22746 199 22806 259
rect 23370 199 23430 259
rect 23994 199 24054 259
rect 24618 199 24678 259
rect 25242 199 25302 259
rect 25866 199 25926 259
rect 26490 199 26550 259
rect 27114 199 27174 259
rect 27738 199 27798 259
rect 28362 199 28422 259
rect 28986 199 29046 259
rect 29610 199 29670 259
rect 30234 199 30294 259
rect 30858 199 30918 259
rect 31482 199 31542 259
rect 32106 199 32166 259
rect 32730 199 32790 259
rect 33354 199 33414 259
rect 33978 199 34038 259
rect 34602 199 34662 259
rect 35226 199 35286 259
rect 35850 199 35910 259
rect 36474 199 36534 259
rect 37098 199 37158 259
rect 37722 199 37782 259
rect 38346 199 38406 259
rect 38970 199 39030 259
rect 39594 199 39654 259
rect 40218 199 40278 259
rect 40842 199 40902 259
rect 41447 180 41545 278
use bitcell_array  bitcell_array_0
timestamp 1676037725
transform 1 0 1248 0 1 790
box -42 -105 39978 50665
use col_cap_array  col_cap_array_0
timestamp 1676037725
transform 1 0 1248 0 -1 52140
box 0 0 39936 474
use col_cap_array  col_cap_array_1
timestamp 1676037725
transform 1 0 1248 0 1 0
box 0 0 39936 474
use dummy_array  dummy_array_0
timestamp 1676037725
transform 1 0 1248 0 1 51350
box -42 -105 39978 421
use dummy_array  dummy_array_1
timestamp 1676037725
transform 1 0 1248 0 -1 790
box -42 -105 39978 421
use replica_column  replica_column_0
timestamp 1676037725
transform 1 0 624 0 1 0
box -26 0 666 52140
use replica_column_0  replica_column_0_0
timestamp 1676037725
transform 1 0 41184 0 1 0
box -42 0 650 52140
use row_cap_array  row_cap_array_0
timestamp 1676037725
transform 1 0 0 0 1 0
box -42 419 624 51721
use row_cap_array_0  row_cap_array_0_0
timestamp 1676037725
transform 1 0 41808 0 1 0
box 0 419 666 51721
<< labels >>
rlabel metal1 s 41424 38959 41424 38959 4 vdd
port 1 nsew
rlabel metal1 s 41424 37379 41424 37379 4 vdd
port 1 nsew
rlabel metal1 s 41424 33720 41424 33720 4 vdd
port 1 nsew
rlabel metal1 s 41424 47150 41424 47150 4 vdd
port 1 nsew
rlabel metal1 s 41424 49229 41424 49229 4 vdd
port 1 nsew
rlabel metal1 s 41424 36589 41424 36589 4 vdd
port 1 nsew
rlabel metal1 s 41424 36880 41424 36880 4 vdd
port 1 nsew
rlabel metal1 s 41424 29770 41424 29770 4 vdd
port 1 nsew
rlabel metal1 s 41424 43990 41424 43990 4 vdd
port 1 nsew
rlabel metal1 s 41424 40040 41424 40040 4 vdd
port 1 nsew
rlabel metal1 s 41424 26319 41424 26319 4 vdd
port 1 nsew
rlabel metal1 s 41424 28190 41424 28190 4 vdd
port 1 nsew
rlabel metal1 s 41424 47649 41424 47649 4 vdd
port 1 nsew
rlabel metal1 s 41424 46859 41424 46859 4 vdd
port 1 nsew
rlabel metal1 s 41424 41620 41424 41620 4 vdd
port 1 nsew
rlabel metal1 s 41424 27400 41424 27400 4 vdd
port 1 nsew
rlabel metal1 s 41424 43200 41424 43200 4 vdd
port 1 nsew
rlabel metal1 s 41424 39250 41424 39250 4 vdd
port 1 nsew
rlabel metal1 s 41424 32639 41424 32639 4 vdd
port 1 nsew
rlabel metal1 s 41424 45570 41424 45570 4 vdd
port 1 nsew
rlabel metal1 s 41424 47940 41424 47940 4 vdd
port 1 nsew
rlabel metal1 s 41424 48439 41424 48439 4 vdd
port 1 nsew
rlabel metal1 s 41424 34510 41424 34510 4 vdd
port 1 nsew
rlabel metal1 s 41424 30269 41424 30269 4 vdd
port 1 nsew
rlabel metal1 s 41424 40539 41424 40539 4 vdd
port 1 nsew
rlabel metal1 s 41424 32930 41424 32930 4 vdd
port 1 nsew
rlabel metal1 s 41424 50019 41424 50019 4 vdd
port 1 nsew
rlabel metal1 s 41424 40830 41424 40830 4 vdd
port 1 nsew
rlabel metal1 s 41424 42410 41424 42410 4 vdd
port 1 nsew
rlabel metal1 s 41424 44780 41424 44780 4 vdd
port 1 nsew
rlabel metal1 s 41424 35799 41424 35799 4 vdd
port 1 nsew
rlabel metal1 s 41424 51599 41424 51599 4 vdd
port 1 nsew
rlabel metal1 s 41424 28689 41424 28689 4 vdd
port 1 nsew
rlabel metal1 s 41424 30560 41424 30560 4 vdd
port 1 nsew
rlabel metal1 s 41424 48730 41424 48730 4 vdd
port 1 nsew
rlabel metal1 s 41424 51100 41424 51100 4 vdd
port 1 nsew
rlabel metal1 s 41424 42119 41424 42119 4 vdd
port 1 nsew
rlabel metal1 s 41424 42909 41424 42909 4 vdd
port 1 nsew
rlabel metal1 s 41424 38169 41424 38169 4 vdd
port 1 nsew
rlabel metal1 s 41424 27899 41424 27899 4 vdd
port 1 nsew
rlabel metal1 s 41424 35300 41424 35300 4 vdd
port 1 nsew
rlabel metal1 s 41424 26610 41424 26610 4 vdd
port 1 nsew
rlabel metal1 s 41424 34219 41424 34219 4 vdd
port 1 nsew
rlabel metal1 s 41424 50310 41424 50310 4 vdd
port 1 nsew
rlabel metal1 s 41424 39749 41424 39749 4 vdd
port 1 nsew
rlabel metal1 s 41424 38460 41424 38460 4 vdd
port 1 nsew
rlabel metal1 s 41424 41329 41424 41329 4 vdd
port 1 nsew
rlabel metal1 s 41424 33429 41424 33429 4 vdd
port 1 nsew
rlabel metal1 s 41424 31350 41424 31350 4 vdd
port 1 nsew
rlabel metal1 s 41424 44489 41424 44489 4 vdd
port 1 nsew
rlabel metal1 s 41424 49520 41424 49520 4 vdd
port 1 nsew
rlabel metal1 s 41424 31059 41424 31059 4 vdd
port 1 nsew
rlabel metal1 s 41424 27109 41424 27109 4 vdd
port 1 nsew
rlabel metal1 s 41424 43699 41424 43699 4 vdd
port 1 nsew
rlabel metal1 s 41424 36090 41424 36090 4 vdd
port 1 nsew
rlabel metal1 s 41424 46069 41424 46069 4 vdd
port 1 nsew
rlabel metal1 s 41424 45279 41424 45279 4 vdd
port 1 nsew
rlabel metal1 s 41424 28980 41424 28980 4 vdd
port 1 nsew
rlabel metal1 s 41424 46360 41424 46360 4 vdd
port 1 nsew
rlabel metal1 s 41424 50809 41424 50809 4 vdd
port 1 nsew
rlabel metal1 s 41424 32140 41424 32140 4 vdd
port 1 nsew
rlabel metal1 s 41424 29479 41424 29479 4 vdd
port 1 nsew
rlabel metal1 s 41424 37670 41424 37670 4 vdd
port 1 nsew
rlabel metal1 s 41424 31849 41424 31849 4 vdd
port 1 nsew
rlabel metal1 s 41424 35009 41424 35009 4 vdd
port 1 nsew
rlabel metal1 s 1008 46360 1008 46360 4 vdd
port 1 nsew
rlabel metal1 s 1008 36880 1008 36880 4 vdd
port 1 nsew
rlabel metal1 s 1008 39749 1008 39749 4 vdd
port 1 nsew
rlabel metal1 s 1008 48439 1008 48439 4 vdd
port 1 nsew
rlabel metal1 s 1008 45570 1008 45570 4 vdd
port 1 nsew
rlabel metal1 s 1008 43990 1008 43990 4 vdd
port 1 nsew
rlabel metal1 s 1008 42410 1008 42410 4 vdd
port 1 nsew
rlabel metal1 s 1008 28689 1008 28689 4 vdd
port 1 nsew
rlabel metal1 s 1008 30560 1008 30560 4 vdd
port 1 nsew
rlabel metal1 s 1008 42909 1008 42909 4 vdd
port 1 nsew
rlabel metal1 s 1008 26610 1008 26610 4 vdd
port 1 nsew
rlabel metal1 s 1008 27400 1008 27400 4 vdd
port 1 nsew
rlabel metal1 s 1008 50310 1008 50310 4 vdd
port 1 nsew
rlabel metal1 s 1008 32930 1008 32930 4 vdd
port 1 nsew
rlabel metal1 s 1008 46859 1008 46859 4 vdd
port 1 nsew
rlabel metal1 s 1008 41620 1008 41620 4 vdd
port 1 nsew
rlabel metal1 s 1008 34510 1008 34510 4 vdd
port 1 nsew
rlabel metal1 s 1008 48730 1008 48730 4 vdd
port 1 nsew
rlabel metal1 s 1008 32639 1008 32639 4 vdd
port 1 nsew
rlabel metal1 s 1008 44780 1008 44780 4 vdd
port 1 nsew
rlabel metal1 s 1008 27109 1008 27109 4 vdd
port 1 nsew
rlabel metal1 s 1008 47940 1008 47940 4 vdd
port 1 nsew
rlabel metal1 s 1008 50019 1008 50019 4 vdd
port 1 nsew
rlabel metal1 s 1008 40040 1008 40040 4 vdd
port 1 nsew
rlabel metal1 s 1008 38460 1008 38460 4 vdd
port 1 nsew
rlabel metal1 s 1008 35300 1008 35300 4 vdd
port 1 nsew
rlabel metal1 s 1008 37379 1008 37379 4 vdd
port 1 nsew
rlabel metal1 s 1008 50809 1008 50809 4 vdd
port 1 nsew
rlabel metal1 s 1008 36589 1008 36589 4 vdd
port 1 nsew
rlabel metal1 s 1008 41329 1008 41329 4 vdd
port 1 nsew
rlabel metal1 s 1008 31350 1008 31350 4 vdd
port 1 nsew
rlabel metal1 s 1008 29770 1008 29770 4 vdd
port 1 nsew
rlabel metal1 s 1008 38169 1008 38169 4 vdd
port 1 nsew
rlabel metal1 s 1008 26319 1008 26319 4 vdd
port 1 nsew
rlabel metal1 s 1008 44489 1008 44489 4 vdd
port 1 nsew
rlabel metal1 s 1008 39250 1008 39250 4 vdd
port 1 nsew
rlabel metal1 s 1008 42119 1008 42119 4 vdd
port 1 nsew
rlabel metal1 s 1008 32140 1008 32140 4 vdd
port 1 nsew
rlabel metal1 s 1008 29479 1008 29479 4 vdd
port 1 nsew
rlabel metal1 s 1008 36090 1008 36090 4 vdd
port 1 nsew
rlabel metal1 s 1008 45279 1008 45279 4 vdd
port 1 nsew
rlabel metal1 s 1008 35799 1008 35799 4 vdd
port 1 nsew
rlabel metal1 s 1008 31059 1008 31059 4 vdd
port 1 nsew
rlabel metal1 s 1008 28980 1008 28980 4 vdd
port 1 nsew
rlabel metal1 s 1008 51599 1008 51599 4 vdd
port 1 nsew
rlabel metal1 s 1008 51100 1008 51100 4 vdd
port 1 nsew
rlabel metal1 s 1008 40539 1008 40539 4 vdd
port 1 nsew
rlabel metal1 s 1008 47150 1008 47150 4 vdd
port 1 nsew
rlabel metal1 s 1008 31849 1008 31849 4 vdd
port 1 nsew
rlabel metal1 s 1008 38959 1008 38959 4 vdd
port 1 nsew
rlabel metal1 s 1008 40830 1008 40830 4 vdd
port 1 nsew
rlabel metal1 s 1008 33720 1008 33720 4 vdd
port 1 nsew
rlabel metal1 s 1008 49520 1008 49520 4 vdd
port 1 nsew
rlabel metal1 s 1008 35009 1008 35009 4 vdd
port 1 nsew
rlabel metal1 s 1008 46069 1008 46069 4 vdd
port 1 nsew
rlabel metal1 s 1008 27899 1008 27899 4 vdd
port 1 nsew
rlabel metal1 s 1008 30269 1008 30269 4 vdd
port 1 nsew
rlabel metal1 s 1008 37670 1008 37670 4 vdd
port 1 nsew
rlabel metal1 s 1008 49229 1008 49229 4 vdd
port 1 nsew
rlabel metal1 s 1008 43699 1008 43699 4 vdd
port 1 nsew
rlabel metal1 s 1008 47649 1008 47649 4 vdd
port 1 nsew
rlabel metal1 s 1008 33429 1008 33429 4 vdd
port 1 nsew
rlabel metal1 s 1008 28190 1008 28190 4 vdd
port 1 nsew
rlabel metal1 s 1008 43200 1008 43200 4 vdd
port 1 nsew
rlabel metal1 s 1008 34219 1008 34219 4 vdd
port 1 nsew
rlabel metal1 s 11544 26070 11544 26070 4 bl1_16
port 1804 nsew
rlabel metal1 s 16608 26070 16608 26070 4 br1_24
port 1837 nsew
rlabel metal1 s 12168 26070 12168 26070 4 bl1_17
port 1808 nsew
rlabel metal1 s 17376 26070 17376 26070 4 bl0_25
port 1838 nsew
rlabel metal1 s 20904 26070 20904 26070 4 bl1_31
port 1864 nsew
rlabel metal1 s 15072 26070 15072 26070 4 bl0_22
port 1826 nsew
rlabel metal1 s 14880 26070 14880 26070 4 bl0_21
port 1822 nsew
rlabel metal1 s 19104 26070 19104 26070 4 br1_28
port 1853 nsew
rlabel metal1 s 18408 26070 18408 26070 4 bl1_27
port 1848 nsew
rlabel metal1 s 17640 26070 17640 26070 4 br0_26
port 1843 nsew
rlabel metal1 s 17304 26070 17304 26070 4 br0_25
port 1839 nsew
rlabel metal1 s 17088 26070 17088 26070 4 br1_25
port 1841 nsew
rlabel metal1 s 16392 26070 16392 26070 4 br0_24
port 1835 nsew
rlabel metal1 s 12648 26070 12648 26070 4 br0_18
port 1811 nsew
rlabel metal1 s 12312 26070 12312 26070 4 br0_17
port 1807 nsew
rlabel metal1 s 11400 26070 11400 26070 4 br0_16
port 1803 nsew
rlabel metal1 s 12096 26070 12096 26070 4 br1_17
port 1809 nsew
rlabel metal1 s 14808 26070 14808 26070 4 br0_21
port 1823 nsew
rlabel metal1 s 20280 26070 20280 26070 4 bl1_30
port 1860 nsew
rlabel metal1 s 14664 26070 14664 26070 4 bl1_21
port 1824 nsew
rlabel metal1 s 21120 26070 21120 26070 4 bl0_31
port 1862 nsew
rlabel metal1 s 17568 26070 17568 26070 4 bl0_26
port 1842 nsew
rlabel metal1 s 16128 26070 16128 26070 4 bl0_23
port 1830 nsew
rlabel metal1 s 14040 26070 14040 26070 4 bl1_20
port 1820 nsew
rlabel metal1 s 13560 26070 13560 26070 4 br0_19
port 1815 nsew
rlabel metal1 s 12864 26070 12864 26070 4 br1_18
port 1813 nsew
rlabel metal1 s 11136 26070 11136 26070 4 bl0_15
port 1798 nsew
rlabel metal1 s 20064 26070 20064 26070 4 bl0_30
port 1858 nsew
rlabel metal1 s 20832 26070 20832 26070 4 br1_31
port 1865 nsew
rlabel metal1 s 16320 26070 16320 26070 4 bl0_24
port 1834 nsew
rlabel metal1 s 19872 26070 19872 26070 4 bl0_29
port 1854 nsew
rlabel metal1 s 15288 26070 15288 26070 4 bl1_22
port 1828 nsew
rlabel metal1 s 15360 26070 15360 26070 4 br1_22
port 1829 nsew
rlabel metal1 s 15840 26070 15840 26070 4 br1_23
port 1833 nsew
rlabel metal1 s 18552 26070 18552 26070 4 br0_27
port 1847 nsew
rlabel metal1 s 21048 26070 21048 26070 4 br0_31
port 1863 nsew
rlabel metal1 s 20136 26070 20136 26070 4 br0_30
port 1859 nsew
rlabel metal1 s 11064 26070 11064 26070 4 br0_15
port 1799 nsew
rlabel metal1 s 19584 26070 19584 26070 4 br1_29
port 1857 nsew
rlabel metal1 s 16536 26070 16536 26070 4 bl1_24
port 1836 nsew
rlabel metal1 s 13632 26070 13632 26070 4 bl0_19
port 1814 nsew
rlabel metal1 s 13416 26070 13416 26070 4 bl1_19
port 1816 nsew
rlabel metal1 s 12384 26070 12384 26070 4 bl0_17
port 1806 nsew
rlabel metal1 s 18336 26070 18336 26070 4 br1_27
port 1849 nsew
rlabel metal1 s 17784 26070 17784 26070 4 bl1_26
port 1844 nsew
rlabel metal1 s 18888 26070 18888 26070 4 br0_28
port 1851 nsew
rlabel metal1 s 19656 26070 19656 26070 4 bl1_29
port 1856 nsew
rlabel metal1 s 15912 26070 15912 26070 4 bl1_23
port 1832 nsew
rlabel metal1 s 11328 26070 11328 26070 4 bl0_16
port 1802 nsew
rlabel metal1 s 11616 26070 11616 26070 4 br1_16
port 1805 nsew
rlabel metal1 s 14592 26070 14592 26070 4 br1_21
port 1825 nsew
rlabel metal1 s 12792 26070 12792 26070 4 bl1_18
port 1812 nsew
rlabel metal1 s 16056 26070 16056 26070 4 br0_23
port 1831 nsew
rlabel metal1 s 13824 26070 13824 26070 4 bl0_20
port 1818 nsew
rlabel metal1 s 19032 26070 19032 26070 4 bl1_28
port 1852 nsew
rlabel metal1 s 17856 26070 17856 26070 4 br1_26
port 1845 nsew
rlabel metal1 s 20352 26070 20352 26070 4 br1_30
port 1861 nsew
rlabel metal1 s 13896 26070 13896 26070 4 br0_20
port 1819 nsew
rlabel metal1 s 18624 26070 18624 26070 4 bl0_27
port 1846 nsew
rlabel metal1 s 19800 26070 19800 26070 4 br0_29
port 1855 nsew
rlabel metal1 s 15144 26070 15144 26070 4 br0_22
port 1827 nsew
rlabel metal1 s 12576 26070 12576 26070 4 bl0_18
port 1810 nsew
rlabel metal1 s 17160 26070 17160 26070 4 bl1_25
port 1840 nsew
rlabel metal1 s 13344 26070 13344 26070 4 br1_19
port 1817 nsew
rlabel metal1 s 14112 26070 14112 26070 4 br1_20
port 1821 nsew
rlabel metal1 s 18816 26070 18816 26070 4 bl0_28
port 1850 nsew
rlabel metal1 s 1152 26070 1152 26070 4 rbl_bl0_0
port 1994 nsew
rlabel metal1 s 3648 26070 3648 26070 4 bl0_3
port 1750 nsew
rlabel metal1 s 1008 15550 1008 15550 4 vdd
port 1 nsew
rlabel metal1 s 2664 26070 2664 26070 4 br0_2
port 1747 nsew
rlabel metal1 s 10080 26070 10080 26070 4 bl0_14
port 1794 nsew
rlabel metal1 s 9120 26070 9120 26070 4 br1_12
port 1789 nsew
rlabel metal1 s 9048 26070 9048 26070 4 bl1_12
port 1788 nsew
rlabel metal1 s 1008 25529 1008 25529 4 vdd
port 1 nsew
rlabel metal1 s 3912 26070 3912 26070 4 br0_4
port 1755 nsew
rlabel metal1 s 1008 21870 1008 21870 4 vdd
port 1 nsew
rlabel metal1 s 3840 26070 3840 26070 4 bl0_4
port 1754 nsew
rlabel metal1 s 1008 18710 1008 18710 4 vdd
port 1 nsew
rlabel metal1 s 1008 20290 1008 20290 4 vdd
port 1 nsew
rlabel metal1 s 4056 26070 4056 26070 4 bl1_4
port 1756 nsew
rlabel metal1 s 1008 16340 1008 16340 4 vdd
port 1 nsew
rlabel metal1 s 1008 22660 1008 22660 4 vdd
port 1 nsew
rlabel metal1 s 4680 26070 4680 26070 4 bl1_5
port 1760 nsew
rlabel metal1 s 8904 26070 8904 26070 4 br0_12
port 1787 nsew
rlabel metal1 s 1008 23159 1008 23159 4 vdd
port 1 nsew
rlabel metal1 s 7800 26070 7800 26070 4 bl1_10
port 1780 nsew
rlabel metal1 s 2880 26070 2880 26070 4 br1_2
port 1749 nsew
rlabel metal1 s 1008 18419 1008 18419 4 vdd
port 1 nsew
rlabel metal1 s 1008 23949 1008 23949 4 vdd
port 1 nsew
rlabel metal1 s 1008 22369 1008 22369 4 vdd
port 1 nsew
rlabel metal1 s 10920 26070 10920 26070 4 bl1_15
port 1800 nsew
rlabel metal1 s 8424 26070 8424 26070 4 bl1_11
port 1784 nsew
rlabel metal1 s 1008 15259 1008 15259 4 vdd
port 1 nsew
rlabel metal1 s 1008 13970 1008 13970 4 vdd
port 1 nsew
rlabel metal1 s 1008 19500 1008 19500 4 vdd
port 1 nsew
rlabel metal1 s 1008 17629 1008 17629 4 vdd
port 1 nsew
rlabel metal1 s 1008 21579 1008 21579 4 vdd
port 1 nsew
rlabel metal1 s 9816 26070 9816 26070 4 br0_13
port 1791 nsew
rlabel metal1 s 1008 24739 1008 24739 4 vdd
port 1 nsew
rlabel metal1 s 2592 26070 2592 26070 4 bl0_2
port 1746 nsew
rlabel metal1 s 6072 26070 6072 26070 4 br0_7
port 1767 nsew
rlabel metal1 s 7392 26070 7392 26070 4 bl0_9
port 1774 nsew
rlabel metal1 s 4608 26070 4608 26070 4 br1_5
port 1761 nsew
rlabel metal1 s 1008 14469 1008 14469 4 vdd
port 1 nsew
rlabel metal1 s 1008 17130 1008 17130 4 vdd
port 1 nsew
rlabel metal1 s 2400 26070 2400 26070 4 bl0_1
port 1742 nsew
rlabel metal1 s 1008 25030 1008 25030 4 vdd
port 1 nsew
rlabel metal1 s 5928 26070 5928 26070 4 bl1_7
port 1768 nsew
rlabel metal1 s 1008 23450 1008 23450 4 vdd
port 1 nsew
rlabel metal1 s 1008 25820 1008 25820 4 vdd
port 1 nsew
rlabel metal1 s 7656 26070 7656 26070 4 br0_10
port 1779 nsew
rlabel metal1 s 6336 26070 6336 26070 4 bl0_8
port 1770 nsew
rlabel metal1 s 1344 26070 1344 26070 4 bl0_0
port 1737 nsew
rlabel metal1 s 1008 19999 1008 19999 4 vdd
port 1 nsew
rlabel metal1 s 1008 24240 1008 24240 4 vdd
port 1 nsew
rlabel metal1 s 7104 26070 7104 26070 4 br1_9
port 1777 nsew
rlabel metal1 s 1008 16839 1008 16839 4 vdd
port 1 nsew
rlabel metal1 s 10296 26070 10296 26070 4 bl1_14
port 1796 nsew
rlabel metal1 s 1008 16049 1008 16049 4 vdd
port 1 nsew
rlabel metal1 s 7584 26070 7584 26070 4 bl0_10
port 1778 nsew
rlabel metal1 s 2808 26070 2808 26070 4 bl1_2
port 1748 nsew
rlabel metal1 s 10152 26070 10152 26070 4 br0_14
port 1795 nsew
rlabel metal1 s 7872 26070 7872 26070 4 br1_10
port 1781 nsew
rlabel metal1 s 8640 26070 8640 26070 4 bl0_11
port 1782 nsew
rlabel metal1 s 864 26070 864 26070 4 rbl_br1_0
port 2256 nsew
rlabel metal1 s 10368 26070 10368 26070 4 br1_14
port 1797 nsew
rlabel metal1 s 6144 26070 6144 26070 4 bl0_7
port 1766 nsew
rlabel metal1 s 6624 26070 6624 26070 4 br1_8
port 1773 nsew
rlabel metal1 s 936 26070 936 26070 4 rbl_bl1_0
port 2257 nsew
rlabel metal1 s 5088 26070 5088 26070 4 bl0_6
port 1762 nsew
rlabel metal1 s 8352 26070 8352 26070 4 br1_11
port 1785 nsew
rlabel metal1 s 9672 26070 9672 26070 4 bl1_13
port 1792 nsew
rlabel metal1 s 2184 26070 2184 26070 4 bl1_1
port 1744 nsew
rlabel metal1 s 10848 26070 10848 26070 4 br1_15
port 1801 nsew
rlabel metal1 s 3360 26070 3360 26070 4 br1_3
port 1753 nsew
rlabel metal1 s 2112 26070 2112 26070 4 br1_1
port 1745 nsew
rlabel metal1 s 3432 26070 3432 26070 4 bl1_3
port 1752 nsew
rlabel metal1 s 1560 26070 1560 26070 4 bl1_0
port 1740 nsew
rlabel metal1 s 1008 20789 1008 20789 4 vdd
port 1 nsew
rlabel metal1 s 1416 26070 1416 26070 4 br0_0
port 1739 nsew
rlabel metal1 s 6552 26070 6552 26070 4 bl1_8
port 1772 nsew
rlabel metal1 s 1080 26070 1080 26070 4 rbl_br0_0
port 1995 nsew
rlabel metal1 s 3576 26070 3576 26070 4 br0_3
port 1751 nsew
rlabel metal1 s 4824 26070 4824 26070 4 br0_5
port 1759 nsew
rlabel metal1 s 7320 26070 7320 26070 4 br0_9
port 1775 nsew
rlabel metal1 s 5376 26070 5376 26070 4 br1_6
port 1765 nsew
rlabel metal1 s 2328 26070 2328 26070 4 br0_1
port 1743 nsew
rlabel metal1 s 5304 26070 5304 26070 4 bl1_6
port 1764 nsew
rlabel metal1 s 1008 17920 1008 17920 4 vdd
port 1 nsew
rlabel metal1 s 5160 26070 5160 26070 4 br0_6
port 1763 nsew
rlabel metal1 s 7176 26070 7176 26070 4 bl1_9
port 1776 nsew
rlabel metal1 s 9600 26070 9600 26070 4 br1_13
port 1793 nsew
rlabel metal1 s 1008 21080 1008 21080 4 vdd
port 1 nsew
rlabel metal1 s 1632 26070 1632 26070 4 br1_0
port 1741 nsew
rlabel metal1 s 4128 26070 4128 26070 4 br1_4
port 1757 nsew
rlabel metal1 s 8568 26070 8568 26070 4 br0_11
port 1783 nsew
rlabel metal1 s 8832 26070 8832 26070 4 bl0_12
port 1786 nsew
rlabel metal1 s 4896 26070 4896 26070 4 bl0_5
port 1758 nsew
rlabel metal1 s 1008 13679 1008 13679 4 vdd
port 1 nsew
rlabel metal1 s 1008 19209 1008 19209 4 vdd
port 1 nsew
rlabel metal1 s 6408 26070 6408 26070 4 br0_8
port 1771 nsew
rlabel metal1 s 9888 26070 9888 26070 4 bl0_13
port 1790 nsew
rlabel metal1 s 5856 26070 5856 26070 4 br1_7
port 1769 nsew
rlabel metal1 s 1008 14760 1008 14760 4 vdd
port 1 nsew
rlabel metal1 s 1008 13180 1008 13180 4 vdd
port 1 nsew
rlabel metal1 s 1008 540 1008 540 4 vdd
port 1 nsew
rlabel metal1 s 1008 9729 1008 9729 4 vdd
port 1 nsew
rlabel metal1 s 1008 6860 1008 6860 4 vdd
port 1 nsew
rlabel metal1 s 1008 7650 1008 7650 4 vdd
port 1 nsew
rlabel metal1 s 1008 10020 1008 10020 4 vdd
port 1 nsew
rlabel metal1 s 1008 11309 1008 11309 4 vdd
port 1 nsew
rlabel metal1 s 1008 2910 1008 2910 4 vdd
port 1 nsew
rlabel metal1 s 1008 5280 1008 5280 4 vdd
port 1 nsew
rlabel metal1 s 1008 4989 1008 4989 4 vdd
port 1 nsew
rlabel metal1 s 1008 3700 1008 3700 4 vdd
port 1 nsew
rlabel metal1 s 1008 5779 1008 5779 4 vdd
port 1 nsew
rlabel metal1 s 1008 9230 1008 9230 4 vdd
port 1 nsew
rlabel metal1 s 1008 1039 1008 1039 4 vdd
port 1 nsew
rlabel metal1 s 1008 12889 1008 12889 4 vdd
port 1 nsew
rlabel metal1 s 1008 11600 1008 11600 4 vdd
port 1 nsew
rlabel metal1 s 1008 12390 1008 12390 4 vdd
port 1 nsew
rlabel metal1 s 1008 4199 1008 4199 4 vdd
port 1 nsew
rlabel metal1 s 1008 7359 1008 7359 4 vdd
port 1 nsew
rlabel metal1 s 1008 2120 1008 2120 4 vdd
port 1 nsew
rlabel metal1 s 1008 6569 1008 6569 4 vdd
port 1 nsew
rlabel metal1 s 1008 4490 1008 4490 4 vdd
port 1 nsew
rlabel metal1 s 1008 3409 1008 3409 4 vdd
port 1 nsew
rlabel metal1 s 1008 1829 1008 1829 4 vdd
port 1 nsew
rlabel metal1 s 1008 6070 1008 6070 4 vdd
port 1 nsew
rlabel metal1 s 1008 8149 1008 8149 4 vdd
port 1 nsew
rlabel metal1 s 1008 8440 1008 8440 4 vdd
port 1 nsew
rlabel metal1 s 1008 10810 1008 10810 4 vdd
port 1 nsew
rlabel metal1 s 1008 10519 1008 10519 4 vdd
port 1 nsew
rlabel metal1 s 1008 2619 1008 2619 4 vdd
port 1 nsew
rlabel metal1 s 1008 1330 1008 1330 4 vdd
port 1 nsew
rlabel metal1 s 1008 12099 1008 12099 4 vdd
port 1 nsew
rlabel metal1 s 1008 8939 1008 8939 4 vdd
port 1 nsew
rlabel metal1 s 37344 26070 37344 26070 4 bl0_57
port 1966 nsew
rlabel metal1 s 41424 14760 41424 14760 4 vdd
port 1 nsew
rlabel metal1 s 35808 26070 35808 26070 4 br1_55
port 1961 nsew
rlabel metal1 s 41424 21080 41424 21080 4 vdd
port 1 nsew
rlabel metal1 s 38784 26070 38784 26070 4 bl0_60
port 1978 nsew
rlabel metal1 s 41424 24739 41424 24739 4 vdd
port 1 nsew
rlabel metal1 s 39552 26070 39552 26070 4 br1_61
port 1985 nsew
rlabel metal1 s 37128 26070 37128 26070 4 bl1_57
port 1968 nsew
rlabel metal1 s 41424 19209 41424 19209 4 vdd
port 1 nsew
rlabel metal1 s 41424 25529 41424 25529 4 vdd
port 1 nsew
rlabel metal1 s 41424 21579 41424 21579 4 vdd
port 1 nsew
rlabel metal1 s 41424 24240 41424 24240 4 vdd
port 1 nsew
rlabel metal1 s 32616 26070 32616 26070 4 br0_50
port 1939 nsew
rlabel metal1 s 41424 21870 41424 21870 4 vdd
port 1 nsew
rlabel metal1 s 41424 20290 41424 20290 4 vdd
port 1 nsew
rlabel metal1 s 41424 13970 41424 13970 4 vdd
port 1 nsew
rlabel metal1 s 33792 26070 33792 26070 4 bl0_52
port 1946 nsew
rlabel metal1 s 41424 15550 41424 15550 4 vdd
port 1 nsew
rlabel metal1 s 31584 26070 31584 26070 4 br1_48
port 1933 nsew
rlabel metal1 s 41424 25820 41424 25820 4 vdd
port 1 nsew
rlabel metal1 s 41424 16340 41424 16340 4 vdd
port 1 nsew
rlabel metal1 s 34632 26070 34632 26070 4 bl1_53
port 1952 nsew
rlabel metal1 s 41424 25030 41424 25030 4 vdd
port 1 nsew
rlabel metal1 s 41424 20789 41424 20789 4 vdd
port 1 nsew
rlabel metal1 s 38304 26070 38304 26070 4 br1_59
port 1977 nsew
rlabel metal1 s 39840 26070 39840 26070 4 bl0_61
port 1982 nsew
rlabel metal1 s 37272 26070 37272 26070 4 br0_57
port 1967 nsew
rlabel metal1 s 36288 26070 36288 26070 4 bl0_56
port 1962 nsew
rlabel metal1 s 37608 26070 37608 26070 4 br0_58
port 1971 nsew
rlabel metal1 s 36360 26070 36360 26070 4 br0_56
port 1963 nsew
rlabel metal1 s 41424 18710 41424 18710 4 vdd
port 1 nsew
rlabel metal1 s 39768 26070 39768 26070 4 br0_61
port 1983 nsew
rlabel metal1 s 38376 26070 38376 26070 4 bl1_59
port 1976 nsew
rlabel metal1 s 41424 19500 41424 19500 4 vdd
port 1 nsew
rlabel metal1 s 41424 23949 41424 23949 4 vdd
port 1 nsew
rlabel metal1 s 32064 26070 32064 26070 4 br1_49
port 1937 nsew
rlabel metal1 s 35880 26070 35880 26070 4 bl1_55
port 1960 nsew
rlabel metal1 s 41424 22369 41424 22369 4 vdd
port 1 nsew
rlabel metal1 s 41424 16839 41424 16839 4 vdd
port 1 nsew
rlabel metal1 s 41424 15259 41424 15259 4 vdd
port 1 nsew
rlabel metal1 s 36096 26070 36096 26070 4 bl0_55
port 1958 nsew
rlabel metal1 s 41424 19999 41424 19999 4 vdd
port 1 nsew
rlabel metal1 s 39072 26070 39072 26070 4 br1_60
port 1981 nsew
rlabel metal1 s 38856 26070 38856 26070 4 br0_60
port 1979 nsew
rlabel metal1 s 41424 22660 41424 22660 4 vdd
port 1 nsew
rlabel metal1 s 41424 13679 41424 13679 4 vdd
port 1 nsew
rlabel metal1 s 41280 26070 41280 26070 4 rbl_bl0_1
port 1735 nsew
rlabel metal1 s 35112 26070 35112 26070 4 br0_54
port 1955 nsew
rlabel metal1 s 38592 26070 38592 26070 4 bl0_59
port 1974 nsew
rlabel metal1 s 41424 16049 41424 16049 4 vdd
port 1 nsew
rlabel metal1 s 33384 26070 33384 26070 4 bl1_51
port 1944 nsew
rlabel metal1 s 41424 18419 41424 18419 4 vdd
port 1 nsew
rlabel metal1 s 36024 26070 36024 26070 4 br0_55
port 1959 nsew
rlabel metal1 s 36576 26070 36576 26070 4 br1_56
port 1965 nsew
rlabel metal1 s 32352 26070 32352 26070 4 bl0_49
port 1934 nsew
rlabel metal1 s 35328 26070 35328 26070 4 br1_54
port 1957 nsew
rlabel metal1 s 37752 26070 37752 26070 4 bl1_58
port 1972 nsew
rlabel metal1 s 40800 26070 40800 26070 4 br1_63
port 1993 nsew
rlabel metal1 s 41016 26070 41016 26070 4 br0_63
port 1991 nsew
rlabel metal1 s 41352 26070 41352 26070 4 rbl_br0_1
port 1738 nsew
rlabel metal1 s 40104 26070 40104 26070 4 br0_62
port 1987 nsew
rlabel metal1 s 40320 26070 40320 26070 4 br1_62
port 1989 nsew
rlabel metal1 s 33528 26070 33528 26070 4 br0_51
port 1943 nsew
rlabel metal1 s 37536 26070 37536 26070 4 bl0_58
port 1970 nsew
rlabel metal1 s 35040 26070 35040 26070 4 bl0_54
port 1954 nsew
rlabel metal1 s 34008 26070 34008 26070 4 bl1_52
port 1948 nsew
rlabel metal1 s 34560 26070 34560 26070 4 br1_53
port 1953 nsew
rlabel metal1 s 32544 26070 32544 26070 4 bl0_50
port 1938 nsew
rlabel metal1 s 32280 26070 32280 26070 4 br0_49
port 1935 nsew
rlabel metal1 s 37824 26070 37824 26070 4 br1_58
port 1973 nsew
rlabel metal1 s 40872 26070 40872 26070 4 bl1_63
port 1992 nsew
rlabel metal1 s 32136 26070 32136 26070 4 bl1_49
port 1936 nsew
rlabel metal1 s 41424 17130 41424 17130 4 vdd
port 1 nsew
rlabel metal1 s 34776 26070 34776 26070 4 br0_53
port 1951 nsew
rlabel metal1 s 34080 26070 34080 26070 4 br1_52
port 1949 nsew
rlabel metal1 s 39000 26070 39000 26070 4 bl1_60
port 1980 nsew
rlabel metal1 s 32832 26070 32832 26070 4 br1_50
port 1941 nsew
rlabel metal1 s 33864 26070 33864 26070 4 br0_52
port 1947 nsew
rlabel metal1 s 41424 23159 41424 23159 4 vdd
port 1 nsew
rlabel metal1 s 40248 26070 40248 26070 4 bl1_62
port 1988 nsew
rlabel metal1 s 38520 26070 38520 26070 4 br0_59
port 1975 nsew
rlabel metal1 s 39624 26070 39624 26070 4 bl1_61
port 1984 nsew
rlabel metal1 s 41424 23450 41424 23450 4 vdd
port 1 nsew
rlabel metal1 s 41424 17629 41424 17629 4 vdd
port 1 nsew
rlabel metal1 s 41424 14469 41424 14469 4 vdd
port 1 nsew
rlabel metal1 s 41568 26070 41568 26070 4 rbl_br1_1
port 1997 nsew
rlabel metal1 s 41088 26070 41088 26070 4 bl0_63
port 1990 nsew
rlabel metal1 s 35256 26070 35256 26070 4 bl1_54
port 1956 nsew
rlabel metal1 s 33600 26070 33600 26070 4 bl0_51
port 1942 nsew
rlabel metal1 s 40032 26070 40032 26070 4 bl0_62
port 1986 nsew
rlabel metal1 s 41496 26070 41496 26070 4 rbl_bl1_1
port 1996 nsew
rlabel metal1 s 32760 26070 32760 26070 4 bl1_50
port 1940 nsew
rlabel metal1 s 34848 26070 34848 26070 4 bl0_53
port 1950 nsew
rlabel metal1 s 31512 26070 31512 26070 4 bl1_48
port 1932 nsew
rlabel metal1 s 37056 26070 37056 26070 4 br1_57
port 1969 nsew
rlabel metal1 s 36504 26070 36504 26070 4 bl1_56
port 1964 nsew
rlabel metal1 s 33312 26070 33312 26070 4 br1_51
port 1945 nsew
rlabel metal1 s 41424 17920 41424 17920 4 vdd
port 1 nsew
rlabel metal1 s 31104 26070 31104 26070 4 bl0_47
port 1926 nsew
rlabel metal1 s 22080 26070 22080 26070 4 br1_33
port 1873 nsew
rlabel metal1 s 27360 26070 27360 26070 4 bl0_41
port 1902 nsew
rlabel metal1 s 24096 26070 24096 26070 4 br1_36
port 1885 nsew
rlabel metal1 s 21312 26070 21312 26070 4 bl0_32
port 1866 nsew
rlabel metal1 s 27624 26070 27624 26070 4 br0_42
port 1907 nsew
rlabel metal1 s 22296 26070 22296 26070 4 br0_33
port 1871 nsew
rlabel metal1 s 28872 26070 28872 26070 4 br0_44
port 1915 nsew
rlabel metal1 s 24576 26070 24576 26070 4 br1_37
port 1889 nsew
rlabel metal1 s 27552 26070 27552 26070 4 bl0_42
port 1906 nsew
rlabel metal1 s 24792 26070 24792 26070 4 br0_37
port 1887 nsew
rlabel metal1 s 22152 26070 22152 26070 4 bl1_33
port 1872 nsew
rlabel metal1 s 31296 26070 31296 26070 4 bl0_48
port 1930 nsew
rlabel metal1 s 27288 26070 27288 26070 4 br0_41
port 1903 nsew
rlabel metal1 s 29640 26070 29640 26070 4 bl1_45
port 1920 nsew
rlabel metal1 s 26520 26070 26520 26070 4 bl1_40
port 1900 nsew
rlabel metal1 s 29856 26070 29856 26070 4 bl0_45
port 1918 nsew
rlabel metal1 s 28536 26070 28536 26070 4 br0_43
port 1911 nsew
rlabel metal1 s 23880 26070 23880 26070 4 br0_36
port 1883 nsew
rlabel metal1 s 29088 26070 29088 26070 4 br1_44
port 1917 nsew
rlabel metal1 s 21384 26070 21384 26070 4 br0_32
port 1867 nsew
rlabel metal1 s 25896 26070 25896 26070 4 bl1_39
port 1896 nsew
rlabel metal1 s 25056 26070 25056 26070 4 bl0_38
port 1890 nsew
rlabel metal1 s 29568 26070 29568 26070 4 br1_45
port 1921 nsew
rlabel metal1 s 31032 26070 31032 26070 4 br0_47
port 1927 nsew
rlabel metal1 s 24648 26070 24648 26070 4 bl1_37
port 1888 nsew
rlabel metal1 s 22560 26070 22560 26070 4 bl0_34
port 1874 nsew
rlabel metal1 s 27768 26070 27768 26070 4 bl1_42
port 1908 nsew
rlabel metal1 s 26112 26070 26112 26070 4 bl0_39
port 1894 nsew
rlabel metal1 s 22368 26070 22368 26070 4 bl0_33
port 1870 nsew
rlabel metal1 s 31368 26070 31368 26070 4 br0_48
port 1931 nsew
rlabel metal1 s 28320 26070 28320 26070 4 br1_43
port 1913 nsew
rlabel metal1 s 28608 26070 28608 26070 4 bl0_43
port 1910 nsew
rlabel metal1 s 24024 26070 24024 26070 4 bl1_36
port 1884 nsew
rlabel metal1 s 21600 26070 21600 26070 4 br1_32
port 1869 nsew
rlabel metal1 s 22632 26070 22632 26070 4 br0_34
port 1875 nsew
rlabel metal1 s 30336 26070 30336 26070 4 br1_46
port 1925 nsew
rlabel metal1 s 25272 26070 25272 26070 4 bl1_38
port 1892 nsew
rlabel metal1 s 30048 26070 30048 26070 4 bl0_46
port 1922 nsew
rlabel metal1 s 30264 26070 30264 26070 4 bl1_46
port 1924 nsew
rlabel metal1 s 27840 26070 27840 26070 4 br1_42
port 1909 nsew
rlabel metal1 s 23400 26070 23400 26070 4 bl1_35
port 1880 nsew
rlabel metal1 s 26304 26070 26304 26070 4 bl0_40
port 1898 nsew
rlabel metal1 s 25344 26070 25344 26070 4 br1_38
port 1893 nsew
rlabel metal1 s 23328 26070 23328 26070 4 br1_35
port 1881 nsew
rlabel metal1 s 30888 26070 30888 26070 4 bl1_47
port 1928 nsew
rlabel metal1 s 26040 26070 26040 26070 4 br0_39
port 1895 nsew
rlabel metal1 s 25128 26070 25128 26070 4 br0_38
port 1891 nsew
rlabel metal1 s 24864 26070 24864 26070 4 bl0_37
port 1886 nsew
rlabel metal1 s 30816 26070 30816 26070 4 br1_47
port 1929 nsew
rlabel metal1 s 26592 26070 26592 26070 4 br1_40
port 1901 nsew
rlabel metal1 s 27072 26070 27072 26070 4 br1_41
port 1905 nsew
rlabel metal1 s 22848 26070 22848 26070 4 br1_34
port 1877 nsew
rlabel metal1 s 28392 26070 28392 26070 4 bl1_43
port 1912 nsew
rlabel metal1 s 21528 26070 21528 26070 4 bl1_32
port 1868 nsew
rlabel metal1 s 26376 26070 26376 26070 4 br0_40
port 1899 nsew
rlabel metal1 s 29016 26070 29016 26070 4 bl1_44
port 1916 nsew
rlabel metal1 s 25824 26070 25824 26070 4 br1_39
port 1897 nsew
rlabel metal1 s 23616 26070 23616 26070 4 bl0_35
port 1878 nsew
rlabel metal1 s 23808 26070 23808 26070 4 bl0_36
port 1882 nsew
rlabel metal1 s 30120 26070 30120 26070 4 br0_46
port 1923 nsew
rlabel metal1 s 27144 26070 27144 26070 4 bl1_41
port 1904 nsew
rlabel metal1 s 29784 26070 29784 26070 4 br0_45
port 1919 nsew
rlabel metal1 s 22776 26070 22776 26070 4 bl1_34
port 1876 nsew
rlabel metal1 s 23544 26070 23544 26070 4 br0_35
port 1879 nsew
rlabel metal1 s 28800 26070 28800 26070 4 bl0_44
port 1914 nsew
rlabel metal1 s 41424 12099 41424 12099 4 vdd
port 1 nsew
rlabel metal1 s 41424 12390 41424 12390 4 vdd
port 1 nsew
rlabel metal1 s 41424 8440 41424 8440 4 vdd
port 1 nsew
rlabel metal1 s 41424 2910 41424 2910 4 vdd
port 1 nsew
rlabel metal1 s 41424 6569 41424 6569 4 vdd
port 1 nsew
rlabel metal1 s 41424 9230 41424 9230 4 vdd
port 1 nsew
rlabel metal1 s 41424 11309 41424 11309 4 vdd
port 1 nsew
rlabel metal1 s 41424 10810 41424 10810 4 vdd
port 1 nsew
rlabel metal1 s 41424 9729 41424 9729 4 vdd
port 1 nsew
rlabel metal1 s 41424 10020 41424 10020 4 vdd
port 1 nsew
rlabel metal1 s 41424 7650 41424 7650 4 vdd
port 1 nsew
rlabel metal1 s 41424 1330 41424 1330 4 vdd
port 1 nsew
rlabel metal1 s 41424 6860 41424 6860 4 vdd
port 1 nsew
rlabel metal1 s 41424 3700 41424 3700 4 vdd
port 1 nsew
rlabel metal1 s 41424 11600 41424 11600 4 vdd
port 1 nsew
rlabel metal1 s 41424 1039 41424 1039 4 vdd
port 1 nsew
rlabel metal1 s 41424 4989 41424 4989 4 vdd
port 1 nsew
rlabel metal1 s 41424 4490 41424 4490 4 vdd
port 1 nsew
rlabel metal1 s 41424 12889 41424 12889 4 vdd
port 1 nsew
rlabel metal1 s 41424 3409 41424 3409 4 vdd
port 1 nsew
rlabel metal1 s 41424 6070 41424 6070 4 vdd
port 1 nsew
rlabel metal1 s 41424 7359 41424 7359 4 vdd
port 1 nsew
rlabel metal1 s 41424 2120 41424 2120 4 vdd
port 1 nsew
rlabel metal1 s 41424 1829 41424 1829 4 vdd
port 1 nsew
rlabel metal1 s 41424 8939 41424 8939 4 vdd
port 1 nsew
rlabel metal1 s 41424 8149 41424 8149 4 vdd
port 1 nsew
rlabel metal1 s 41424 13180 41424 13180 4 vdd
port 1 nsew
rlabel metal1 s 41424 10519 41424 10519 4 vdd
port 1 nsew
rlabel metal1 s 41424 4199 41424 4199 4 vdd
port 1 nsew
rlabel metal1 s 41424 5280 41424 5280 4 vdd
port 1 nsew
rlabel metal1 s 41424 2619 41424 2619 4 vdd
port 1 nsew
rlabel metal1 s 41424 5779 41424 5779 4 vdd
port 1 nsew
rlabel metal1 s 41424 540 41424 540 4 vdd
port 1 nsew
rlabel metal2 s 41424 33970 41424 33970 4 gnd
port 2 nsew
rlabel metal2 s 41424 45267 41424 45267 4 gnd
port 2 nsew
rlabel metal2 s 41424 29467 41424 29467 4 gnd
port 2 nsew
rlabel metal2 s 41424 34760 41424 34760 4 gnd
port 2 nsew
rlabel metal2 s 41424 42660 41424 42660 4 gnd
port 2 nsew
rlabel metal2 s 41424 44793 41424 44793 4 gnd
port 2 nsew
rlabel metal2 s 41424 48980 41424 48980 4 gnd
port 2 nsew
rlabel metal2 s 41424 38947 41424 38947 4 gnd
port 2 nsew
rlabel metal2 s 41424 47163 41424 47163 4 gnd
port 2 nsew
rlabel metal2 s 41424 39737 41424 39737 4 gnd
port 2 nsew
rlabel metal2 s 41424 49770 41424 49770 4 gnd
port 2 nsew
rlabel metal2 s 41424 36340 41424 36340 4 gnd
port 2 nsew
rlabel metal2 s 41424 46847 41424 46847 4 gnd
port 2 nsew
rlabel metal2 s 41424 33417 41424 33417 4 gnd
port 2 nsew
rlabel metal2 s 41424 37920 41424 37920 4 gnd
port 2 nsew
rlabel metal2 s 41424 46057 41424 46057 4 gnd
port 2 nsew
rlabel metal2 s 41424 35313 41424 35313 4 gnd
port 2 nsew
rlabel metal2 s 41424 47953 41424 47953 4 gnd
port 2 nsew
rlabel metal2 s 41424 41633 41424 41633 4 gnd
port 2 nsew
rlabel metal2 s 41424 43213 41424 43213 4 gnd
port 2 nsew
rlabel metal2 s 41424 30257 41424 30257 4 gnd
port 2 nsew
rlabel metal2 s 41424 42897 41424 42897 4 gnd
port 2 nsew
rlabel metal2 s 41424 43687 41424 43687 4 gnd
port 2 nsew
rlabel metal2 s 41424 40053 41424 40053 4 gnd
port 2 nsew
rlabel metal2 s 41424 27887 41424 27887 4 gnd
port 2 nsew
rlabel metal2 s 41424 43450 41424 43450 4 gnd
port 2 nsew
rlabel metal2 s 41424 44240 41424 44240 4 gnd
port 2 nsew
rlabel metal2 s 41424 48743 41424 48743 4 gnd
port 2 nsew
rlabel metal2 s 41424 28677 41424 28677 4 gnd
port 2 nsew
rlabel metal2 s 41424 46610 41424 46610 4 gnd
port 2 nsew
rlabel metal2 s 41424 30020 41424 30020 4 gnd
port 2 nsew
rlabel metal2 s 41424 50797 41424 50797 4 gnd
port 2 nsew
rlabel metal2 s 41424 38710 41424 38710 4 gnd
port 2 nsew
rlabel metal2 s 41424 42423 41424 42423 4 gnd
port 2 nsew
rlabel metal2 s 41424 30573 41424 30573 4 gnd
port 2 nsew
rlabel metal2 s 41424 45030 41424 45030 4 gnd
port 2 nsew
rlabel metal2 s 41424 51113 41424 51113 4 gnd
port 2 nsew
rlabel metal2 s 41424 31363 41424 31363 4 gnd
port 2 nsew
rlabel metal2 s 41424 50007 41424 50007 4 gnd
port 2 nsew
rlabel metal2 s 41424 41080 41424 41080 4 gnd
port 2 nsew
rlabel metal2 s 41424 34207 41424 34207 4 gnd
port 2 nsew
rlabel metal2 s 41424 35550 41424 35550 4 gnd
port 2 nsew
rlabel metal2 s 41424 51587 41424 51587 4 gnd
port 2 nsew
rlabel metal2 s 41424 44003 41424 44003 4 gnd
port 2 nsew
rlabel metal2 s 41424 36577 41424 36577 4 gnd
port 2 nsew
rlabel metal2 s 41424 26307 41424 26307 4 gnd
port 2 nsew
rlabel metal2 s 41424 33180 41424 33180 4 gnd
port 2 nsew
rlabel metal2 s 41424 29230 41424 29230 4 gnd
port 2 nsew
rlabel metal2 s 41424 38473 41424 38473 4 gnd
port 2 nsew
rlabel metal2 s 41424 39263 41424 39263 4 gnd
port 2 nsew
rlabel metal2 s 41424 32943 41424 32943 4 gnd
port 2 nsew
rlabel metal2 s 41424 40527 41424 40527 4 gnd
port 2 nsew
rlabel metal2 s 41424 44477 41424 44477 4 gnd
port 2 nsew
rlabel metal2 s 41424 49217 41424 49217 4 gnd
port 2 nsew
rlabel metal2 s 41424 36103 41424 36103 4 gnd
port 2 nsew
rlabel metal2 s 41424 28993 41424 28993 4 gnd
port 2 nsew
rlabel metal2 s 41424 31047 41424 31047 4 gnd
port 2 nsew
rlabel metal2 s 41424 40290 41424 40290 4 gnd
port 2 nsew
rlabel metal2 s 41424 31837 41424 31837 4 gnd
port 2 nsew
rlabel metal2 s 41424 27650 41424 27650 4 gnd
port 2 nsew
rlabel metal2 s 41424 37683 41424 37683 4 gnd
port 2 nsew
rlabel metal2 s 41424 41870 41424 41870 4 gnd
port 2 nsew
rlabel metal2 s 41424 41317 41424 41317 4 gnd
port 2 nsew
rlabel metal2 s 41424 32627 41424 32627 4 gnd
port 2 nsew
rlabel metal2 s 41424 26623 41424 26623 4 gnd
port 2 nsew
rlabel metal2 s 41424 50323 41424 50323 4 gnd
port 2 nsew
rlabel metal2 s 41424 28440 41424 28440 4 gnd
port 2 nsew
rlabel metal2 s 41424 31600 41424 31600 4 gnd
port 2 nsew
rlabel metal2 s 41424 26860 41424 26860 4 gnd
port 2 nsew
rlabel metal2 s 41424 29783 41424 29783 4 gnd
port 2 nsew
rlabel metal2 s 41424 30810 41424 30810 4 gnd
port 2 nsew
rlabel metal2 s 41424 40843 41424 40843 4 gnd
port 2 nsew
rlabel metal2 s 41424 37367 41424 37367 4 gnd
port 2 nsew
rlabel metal2 s 41424 49533 41424 49533 4 gnd
port 2 nsew
rlabel metal2 s 41424 37130 41424 37130 4 gnd
port 2 nsew
rlabel metal2 s 41424 45583 41424 45583 4 gnd
port 2 nsew
rlabel metal2 s 41424 42107 41424 42107 4 gnd
port 2 nsew
rlabel metal2 s 41424 36893 41424 36893 4 gnd
port 2 nsew
rlabel metal2 s 41424 28203 41424 28203 4 gnd
port 2 nsew
rlabel metal2 s 41424 32153 41424 32153 4 gnd
port 2 nsew
rlabel metal2 s 41424 48190 41424 48190 4 gnd
port 2 nsew
rlabel metal2 s 41424 27413 41424 27413 4 gnd
port 2 nsew
rlabel metal2 s 41424 34997 41424 34997 4 gnd
port 2 nsew
rlabel metal2 s 41424 39500 41424 39500 4 gnd
port 2 nsew
rlabel metal2 s 41424 51350 41424 51350 4 gnd
port 2 nsew
rlabel metal2 s 41424 47637 41424 47637 4 gnd
port 2 nsew
rlabel metal2 s 41424 34523 41424 34523 4 gnd
port 2 nsew
rlabel metal2 s 41424 35787 41424 35787 4 gnd
port 2 nsew
rlabel metal2 s 41424 33733 41424 33733 4 gnd
port 2 nsew
rlabel metal2 s 41424 47400 41424 47400 4 gnd
port 2 nsew
rlabel metal2 s 41424 50560 41424 50560 4 gnd
port 2 nsew
rlabel metal2 s 41424 32390 41424 32390 4 gnd
port 2 nsew
rlabel metal2 s 41424 45820 41424 45820 4 gnd
port 2 nsew
rlabel metal2 s 41424 26070 41424 26070 4 gnd
port 2 nsew
rlabel metal2 s 41424 48427 41424 48427 4 gnd
port 2 nsew
rlabel metal2 s 41424 27097 41424 27097 4 gnd
port 2 nsew
rlabel metal2 s 41424 38157 41424 38157 4 gnd
port 2 nsew
rlabel metal2 s 41424 46373 41424 46373 4 gnd
port 2 nsew
rlabel metal2 s 21216 51223 21216 51223 4 wl1_127
port 2253 nsew
rlabel metal2 s 21216 43103 21216 43103 4 wl0_107
port 2212 nsew
rlabel metal2 s 21216 50907 21216 50907 4 wl0_126
port 2250 nsew
rlabel metal2 s 21216 48537 21216 48537 4 wl0_120
port 2238 nsew
rlabel metal2 s 21216 46483 21216 46483 4 wl1_115
port 2229 nsew
rlabel metal2 s 21216 39943 21216 39943 4 wl0_99
port 2196 nsew
rlabel metal2 s 21216 38837 21216 38837 4 wl1_96
port 2191 nsew
rlabel metal2 s 21216 50433 21216 50433 4 wl1_125
port 2249 nsew
rlabel metal2 s 21216 45693 21216 45693 4 wl1_113
port 2225 nsew
rlabel metal2 s 21216 47747 21216 47747 4 wl0_118
port 2234 nsew
rlabel metal2 s 21216 46957 21216 46957 4 wl0_116
port 2230 nsew
rlabel metal2 s 21216 40637 21216 40637 4 wl0_100
port 2198 nsew
rlabel metal2 s 21216 43323 21216 43323 4 wl1_107
port 2213 nsew
rlabel metal2 s 21216 44683 21216 44683 4 wl0_111
port 2220 nsew
rlabel metal2 s 21216 46737 21216 46737 4 wl1_116
port 2231 nsew
rlabel metal2 s 21216 39373 21216 39373 4 wl1_97
port 2193 nsew
rlabel metal2 s 21216 51003 21216 51003 4 wl0_127
port 2252 nsew
rlabel metal2 s 21216 40163 21216 40163 4 wl1_99
port 2197 nsew
rlabel metal2 s 21216 42217 21216 42217 4 wl0_104
port 2206 nsew
rlabel metal2 s 21216 47843 21216 47843 4 wl0_119
port 2236 nsew
rlabel metal2 s 21216 45473 21216 45473 4 wl0_113
port 2224 nsew
rlabel metal2 s 21216 41207 21216 41207 4 wl1_102
port 2203 nsew
rlabel metal2 s 21216 49897 21216 49897 4 wl1_124
port 2247 nsew
rlabel metal2 s 21216 45377 21216 45377 4 wl0_112
port 2222 nsew
rlabel metal2 s 21216 49423 21216 49423 4 wl0_123
port 2244 nsew
rlabel metal2 s 21216 45947 21216 45947 4 wl1_114
port 2227 nsew
rlabel metal2 s 21216 43007 21216 43007 4 wl0_106
port 2210 nsew
rlabel metal2 s 21216 47053 21216 47053 4 wl0_117
port 2232 nsew
rlabel metal2 s 21216 49327 21216 49327 4 wl0_122
port 2242 nsew
rlabel metal2 s 21216 44587 21216 44587 4 wl0_110
port 2218 nsew
rlabel metal2 s 21216 43577 21216 43577 4 wl1_108
port 2215 nsew
rlabel metal2 s 21216 43893 21216 43893 4 wl0_109
port 2216 nsew
rlabel metal2 s 21216 39057 21216 39057 4 wl0_96
port 2190 nsew
rlabel metal2 s 21216 41427 21216 41427 4 wl0_102
port 2202 nsew
rlabel metal2 s 21216 48063 21216 48063 4 wl1_119
port 2237 nsew
rlabel metal2 s 21216 40417 21216 40417 4 wl1_100
port 2199 nsew
rlabel metal2 s 21216 50687 21216 50687 4 wl1_126
port 2251 nsew
rlabel metal2 s 21216 43797 21216 43797 4 wl0_108
port 2214 nsew
rlabel metal2 s 21216 44367 21216 44367 4 wl1_110
port 2219 nsew
rlabel metal2 s 21216 40733 21216 40733 4 wl0_101
port 2200 nsew
rlabel metal2 s 21216 44903 21216 44903 4 wl1_111
port 2221 nsew
rlabel metal2 s 21216 50117 21216 50117 4 wl0_124
port 2246 nsew
rlabel metal2 s 21216 45157 21216 45157 4 wl1_112
port 2223 nsew
rlabel metal2 s 21216 39847 21216 39847 4 wl0_98
port 2194 nsew
rlabel metal2 s 21216 49643 21216 49643 4 wl1_123
port 2245 nsew
rlabel metal2 s 21216 42313 21216 42313 4 wl0_105
port 2208 nsew
rlabel metal2 s 21216 46263 21216 46263 4 wl0_115
port 2228 nsew
rlabel metal2 s 21216 49107 21216 49107 4 wl1_122
port 2243 nsew
rlabel metal2 s 21216 48853 21216 48853 4 wl1_121
port 2241 nsew
rlabel metal2 s 21216 48633 21216 48633 4 wl0_121
port 2240 nsew
rlabel metal2 s 21216 41743 21216 41743 4 wl1_103
port 2205 nsew
rlabel metal2 s 21216 39627 21216 39627 4 wl1_98
port 2195 nsew
rlabel metal2 s 21216 39153 21216 39153 4 wl0_97
port 2192 nsew
rlabel metal2 s 21216 42787 21216 42787 4 wl1_106
port 2211 nsew
rlabel metal2 s 21216 40953 21216 40953 4 wl1_101
port 2201 nsew
rlabel metal2 s 21216 47527 21216 47527 4 wl1_118
port 2235 nsew
rlabel metal2 s 21216 47273 21216 47273 4 wl1_117
port 2233 nsew
rlabel metal2 s 21216 41523 21216 41523 4 wl0_103
port 2204 nsew
rlabel metal2 s 21216 50213 21216 50213 4 wl0_125
port 2248 nsew
rlabel metal2 s 21216 42533 21216 42533 4 wl1_105
port 2209 nsew
rlabel metal2 s 21216 51477 21216 51477 4 rbl_wl1_1
port 2255 nsew
rlabel metal2 s 21216 46167 21216 46167 4 wl0_114
port 2226 nsew
rlabel metal2 s 21216 44113 21216 44113 4 wl1_109
port 2217 nsew
rlabel metal2 s 21216 41997 21216 41997 4 wl1_104
port 2207 nsew
rlabel metal2 s 21216 48317 21216 48317 4 wl1_120
port 2239 nsew
rlabel metal2 s 1008 50797 1008 50797 4 gnd
port 2 nsew
rlabel metal2 s 1008 47637 1008 47637 4 gnd
port 2 nsew
rlabel metal2 s 1008 45583 1008 45583 4 gnd
port 2 nsew
rlabel metal2 s 1008 46373 1008 46373 4 gnd
port 2 nsew
rlabel metal2 s 1008 42897 1008 42897 4 gnd
port 2 nsew
rlabel metal2 s 1008 40843 1008 40843 4 gnd
port 2 nsew
rlabel metal2 s 1008 47953 1008 47953 4 gnd
port 2 nsew
rlabel metal2 s 1008 48427 1008 48427 4 gnd
port 2 nsew
rlabel metal2 s 1008 38947 1008 38947 4 gnd
port 2 nsew
rlabel metal2 s 1008 43687 1008 43687 4 gnd
port 2 nsew
rlabel metal2 s 1008 46847 1008 46847 4 gnd
port 2 nsew
rlabel metal2 s 1008 46610 1008 46610 4 gnd
port 2 nsew
rlabel metal2 s 1008 44003 1008 44003 4 gnd
port 2 nsew
rlabel metal2 s 1008 41080 1008 41080 4 gnd
port 2 nsew
rlabel metal2 s 1008 41317 1008 41317 4 gnd
port 2 nsew
rlabel metal2 s 1008 49770 1008 49770 4 gnd
port 2 nsew
rlabel metal2 s 1008 45267 1008 45267 4 gnd
port 2 nsew
rlabel metal2 s 1008 39263 1008 39263 4 gnd
port 2 nsew
rlabel metal2 s 1008 44240 1008 44240 4 gnd
port 2 nsew
rlabel metal2 s 1008 39737 1008 39737 4 gnd
port 2 nsew
rlabel metal2 s 1008 42423 1008 42423 4 gnd
port 2 nsew
rlabel metal2 s 1008 47163 1008 47163 4 gnd
port 2 nsew
rlabel metal2 s 1008 48190 1008 48190 4 gnd
port 2 nsew
rlabel metal2 s 1008 45030 1008 45030 4 gnd
port 2 nsew
rlabel metal2 s 1008 50007 1008 50007 4 gnd
port 2 nsew
rlabel metal2 s 1008 42107 1008 42107 4 gnd
port 2 nsew
rlabel metal2 s 1008 50560 1008 50560 4 gnd
port 2 nsew
rlabel metal2 s 1008 41633 1008 41633 4 gnd
port 2 nsew
rlabel metal2 s 1008 49217 1008 49217 4 gnd
port 2 nsew
rlabel metal2 s 1008 41870 1008 41870 4 gnd
port 2 nsew
rlabel metal2 s 1008 47400 1008 47400 4 gnd
port 2 nsew
rlabel metal2 s 1008 49533 1008 49533 4 gnd
port 2 nsew
rlabel metal2 s 1008 50323 1008 50323 4 gnd
port 2 nsew
rlabel metal2 s 1008 40527 1008 40527 4 gnd
port 2 nsew
rlabel metal2 s 1008 45820 1008 45820 4 gnd
port 2 nsew
rlabel metal2 s 1008 44793 1008 44793 4 gnd
port 2 nsew
rlabel metal2 s 1008 43213 1008 43213 4 gnd
port 2 nsew
rlabel metal2 s 1008 40053 1008 40053 4 gnd
port 2 nsew
rlabel metal2 s 1008 40290 1008 40290 4 gnd
port 2 nsew
rlabel metal2 s 1008 48743 1008 48743 4 gnd
port 2 nsew
rlabel metal2 s 1008 51113 1008 51113 4 gnd
port 2 nsew
rlabel metal2 s 1008 51350 1008 51350 4 gnd
port 2 nsew
rlabel metal2 s 1008 43450 1008 43450 4 gnd
port 2 nsew
rlabel metal2 s 1008 42660 1008 42660 4 gnd
port 2 nsew
rlabel metal2 s 1008 44477 1008 44477 4 gnd
port 2 nsew
rlabel metal2 s 1008 46057 1008 46057 4 gnd
port 2 nsew
rlabel metal2 s 1008 39500 1008 39500 4 gnd
port 2 nsew
rlabel metal2 s 1008 48980 1008 48980 4 gnd
port 2 nsew
rlabel metal2 s 1008 51587 1008 51587 4 gnd
port 2 nsew
rlabel metal2 s 1008 29230 1008 29230 4 gnd
port 2 nsew
rlabel metal2 s 1008 37367 1008 37367 4 gnd
port 2 nsew
rlabel metal2 s 1008 27650 1008 27650 4 gnd
port 2 nsew
rlabel metal2 s 1008 30257 1008 30257 4 gnd
port 2 nsew
rlabel metal2 s 1008 37130 1008 37130 4 gnd
port 2 nsew
rlabel metal2 s 1008 35313 1008 35313 4 gnd
port 2 nsew
rlabel metal2 s 1008 29783 1008 29783 4 gnd
port 2 nsew
rlabel metal2 s 1008 36103 1008 36103 4 gnd
port 2 nsew
rlabel metal2 s 1008 28677 1008 28677 4 gnd
port 2 nsew
rlabel metal2 s 1008 27887 1008 27887 4 gnd
port 2 nsew
rlabel metal2 s 1008 33733 1008 33733 4 gnd
port 2 nsew
rlabel metal2 s 1008 35787 1008 35787 4 gnd
port 2 nsew
rlabel metal2 s 1008 31837 1008 31837 4 gnd
port 2 nsew
rlabel metal2 s 1008 38157 1008 38157 4 gnd
port 2 nsew
rlabel metal2 s 1008 32390 1008 32390 4 gnd
port 2 nsew
rlabel metal2 s 1008 31600 1008 31600 4 gnd
port 2 nsew
rlabel metal2 s 1008 28203 1008 28203 4 gnd
port 2 nsew
rlabel metal2 s 1008 38473 1008 38473 4 gnd
port 2 nsew
rlabel metal2 s 1008 27413 1008 27413 4 gnd
port 2 nsew
rlabel metal2 s 1008 38710 1008 38710 4 gnd
port 2 nsew
rlabel metal2 s 1008 36340 1008 36340 4 gnd
port 2 nsew
rlabel metal2 s 1008 32943 1008 32943 4 gnd
port 2 nsew
rlabel metal2 s 1008 30020 1008 30020 4 gnd
port 2 nsew
rlabel metal2 s 1008 28993 1008 28993 4 gnd
port 2 nsew
rlabel metal2 s 1008 26307 1008 26307 4 gnd
port 2 nsew
rlabel metal2 s 1008 31047 1008 31047 4 gnd
port 2 nsew
rlabel metal2 s 1008 37920 1008 37920 4 gnd
port 2 nsew
rlabel metal2 s 1008 31363 1008 31363 4 gnd
port 2 nsew
rlabel metal2 s 1008 26070 1008 26070 4 gnd
port 2 nsew
rlabel metal2 s 1008 34207 1008 34207 4 gnd
port 2 nsew
rlabel metal2 s 1008 30810 1008 30810 4 gnd
port 2 nsew
rlabel metal2 s 1008 34523 1008 34523 4 gnd
port 2 nsew
rlabel metal2 s 1008 34760 1008 34760 4 gnd
port 2 nsew
rlabel metal2 s 1008 34997 1008 34997 4 gnd
port 2 nsew
rlabel metal2 s 1008 27097 1008 27097 4 gnd
port 2 nsew
rlabel metal2 s 1008 35550 1008 35550 4 gnd
port 2 nsew
rlabel metal2 s 1008 36577 1008 36577 4 gnd
port 2 nsew
rlabel metal2 s 1008 30573 1008 30573 4 gnd
port 2 nsew
rlabel metal2 s 1008 29467 1008 29467 4 gnd
port 2 nsew
rlabel metal2 s 1008 36893 1008 36893 4 gnd
port 2 nsew
rlabel metal2 s 1008 33970 1008 33970 4 gnd
port 2 nsew
rlabel metal2 s 1008 32153 1008 32153 4 gnd
port 2 nsew
rlabel metal2 s 1008 33180 1008 33180 4 gnd
port 2 nsew
rlabel metal2 s 1008 28440 1008 28440 4 gnd
port 2 nsew
rlabel metal2 s 1008 32627 1008 32627 4 gnd
port 2 nsew
rlabel metal2 s 1008 33417 1008 33417 4 gnd
port 2 nsew
rlabel metal2 s 1008 26623 1008 26623 4 gnd
port 2 nsew
rlabel metal2 s 1008 37683 1008 37683 4 gnd
port 2 nsew
rlabel metal2 s 1008 26860 1008 26860 4 gnd
port 2 nsew
rlabel metal2 s 21216 29893 21216 29893 4 wl1_73
port 2145 nsew
rlabel metal2 s 21216 30463 21216 30463 4 wl0_75
port 2148 nsew
rlabel metal2 s 21216 33053 21216 33053 4 wl1_81
port 2161 nsew
rlabel metal2 s 21216 33843 21216 33843 4 wl1_83
port 2165 nsew
rlabel metal2 s 21216 33527 21216 33527 4 wl0_82
port 2162 nsew
rlabel metal2 s 21216 29357 21216 29357 4 wl1_72
port 2143 nsew
rlabel metal2 s 21216 30367 21216 30367 4 wl0_74
port 2146 nsew
rlabel metal2 s 21216 26197 21216 26197 4 wl1_64
port 2127 nsew
rlabel metal2 s 21216 31473 21216 31473 4 wl1_77
port 2153 nsew
rlabel metal2 s 21216 32263 21216 32263 4 wl1_79
port 2157 nsew
rlabel metal2 s 21216 27777 21216 27777 4 wl1_68
port 2135 nsew
rlabel metal2 s 21216 27523 21216 27523 4 wl1_67
port 2133 nsew
rlabel metal2 s 21216 35897 21216 35897 4 wl0_88
port 2174 nsew
rlabel metal2 s 21216 36467 21216 36467 4 wl1_90
port 2179 nsew
rlabel metal2 s 21216 30147 21216 30147 4 wl1_74
port 2147 nsew
rlabel metal2 s 21216 36783 21216 36783 4 wl0_91
port 2180 nsew
rlabel metal2 s 21216 27303 21216 27303 4 wl0_67
port 2132 nsew
rlabel metal2 s 21216 32043 21216 32043 4 wl0_79
port 2156 nsew
rlabel metal2 s 21216 38047 21216 38047 4 wl1_94
port 2187 nsew
rlabel metal2 s 21216 35203 21216 35203 4 wl0_87
port 2172 nsew
rlabel metal2 s 21216 29673 21216 29673 4 wl0_73
port 2144 nsew
rlabel metal2 s 21216 26513 21216 26513 4 wl0_65
port 2128 nsew
rlabel metal2 s 21216 38267 21216 38267 4 wl0_94
port 2186 nsew
rlabel metal2 s 21216 29577 21216 29577 4 wl0_72
port 2142 nsew
rlabel metal2 s 21216 38363 21216 38363 4 wl0_95
port 2188 nsew
rlabel metal2 s 21216 27997 21216 27997 4 wl0_68
port 2134 nsew
rlabel metal2 s 21216 37477 21216 37477 4 wl0_92
port 2182 nsew
rlabel metal2 s 21216 37573 21216 37573 4 wl0_93
port 2184 nsew
rlabel metal2 s 21216 31253 21216 31253 4 wl0_77
port 2152 nsew
rlabel metal2 s 21216 31947 21216 31947 4 wl0_78
port 2154 nsew
rlabel metal2 s 21216 28883 21216 28883 4 wl0_71
port 2140 nsew
rlabel metal2 s 21216 31727 21216 31727 4 wl1_78
port 2155 nsew
rlabel metal2 s 21216 37793 21216 37793 4 wl1_93
port 2185 nsew
rlabel metal2 s 21216 37003 21216 37003 4 wl1_91
port 2181 nsew
rlabel metal2 s 21216 32517 21216 32517 4 wl1_80
port 2159 nsew
rlabel metal2 s 21216 27207 21216 27207 4 wl0_66
port 2130 nsew
rlabel metal2 s 21216 36213 21216 36213 4 wl1_89
port 2177 nsew
rlabel metal2 s 21216 28567 21216 28567 4 wl1_70
port 2139 nsew
rlabel metal2 s 21216 33307 21216 33307 4 wl1_82
port 2163 nsew
rlabel metal2 s 21216 33623 21216 33623 4 wl0_83
port 2164 nsew
rlabel metal2 s 21216 29103 21216 29103 4 wl1_71
port 2141 nsew
rlabel metal2 s 21216 37257 21216 37257 4 wl1_92
port 2183 nsew
rlabel metal2 s 21216 26733 21216 26733 4 wl1_65
port 2129 nsew
rlabel metal2 s 21216 34097 21216 34097 4 wl1_84
port 2167 nsew
rlabel metal2 s 21216 34633 21216 34633 4 wl1_85
port 2169 nsew
rlabel metal2 s 21216 32737 21216 32737 4 wl0_80
port 2158 nsew
rlabel metal2 s 21216 31157 21216 31157 4 wl0_76
port 2150 nsew
rlabel metal2 s 21216 30937 21216 30937 4 wl1_76
port 2151 nsew
rlabel metal2 s 21216 35107 21216 35107 4 wl0_86
port 2170 nsew
rlabel metal2 s 21216 38583 21216 38583 4 wl1_95
port 2189 nsew
rlabel metal2 s 21216 35993 21216 35993 4 wl0_89
port 2176 nsew
rlabel metal2 s 21216 35677 21216 35677 4 wl1_88
port 2175 nsew
rlabel metal2 s 21216 34887 21216 34887 4 wl1_86
port 2171 nsew
rlabel metal2 s 21216 30683 21216 30683 4 wl1_75
port 2149 nsew
rlabel metal2 s 21216 26987 21216 26987 4 wl1_66
port 2131 nsew
rlabel metal2 s 21216 28313 21216 28313 4 wl1_69
port 2137 nsew
rlabel metal2 s 21216 36687 21216 36687 4 wl0_90
port 2178 nsew
rlabel metal2 s 21216 28787 21216 28787 4 wl0_70
port 2138 nsew
rlabel metal2 s 21216 26417 21216 26417 4 wl0_64
port 2126 nsew
rlabel metal2 s 21216 28093 21216 28093 4 wl0_69
port 2136 nsew
rlabel metal2 s 21216 34317 21216 34317 4 wl0_84
port 2166 nsew
rlabel metal2 s 21216 35423 21216 35423 4 wl1_87
port 2173 nsew
rlabel metal2 s 21216 34413 21216 34413 4 wl0_85
port 2168 nsew
rlabel metal2 s 21216 32833 21216 32833 4 wl0_81
port 2160 nsew
rlabel metal2 s 21216 24837 21216 24837 4 wl0_60
port 2118 nsew
rlabel metal2 s 21216 16147 21216 16147 4 wl0_38
port 2074 nsew
rlabel metal2 s 21216 13557 21216 13557 4 wl1_32
port 2063 nsew
rlabel metal2 s 21216 16463 21216 16463 4 wl1_39
port 2077 nsew
rlabel metal2 s 21216 20667 21216 20667 4 wl1_50
port 2099 nsew
rlabel metal2 s 21216 21203 21216 21203 4 wl1_51
port 2101 nsew
rlabel metal2 s 21216 19307 21216 19307 4 wl0_46
port 2090 nsew
rlabel metal2 s 21216 20983 21216 20983 4 wl0_51
port 2100 nsew
rlabel metal2 s 21216 23353 21216 23353 4 wl0_57
port 2112 nsew
rlabel metal2 s 21216 23257 21216 23257 4 wl0_56
port 2110 nsew
rlabel metal2 s 21216 21457 21216 21457 4 wl1_52
port 2103 nsew
rlabel metal2 s 21216 16717 21216 16717 4 wl1_40
port 2079 nsew
rlabel metal2 s 21216 22563 21216 22563 4 wl0_55
port 2108 nsew
rlabel metal2 s 21216 24617 21216 24617 4 wl1_60
port 2119 nsew
rlabel metal2 s 21216 13777 21216 13777 4 wl0_32
port 2062 nsew
rlabel metal2 s 21216 14093 21216 14093 4 wl1_33
port 2065 nsew
rlabel metal2 s 21216 18043 21216 18043 4 wl1_43
port 2085 nsew
rlabel metal2 s 21216 21677 21216 21677 4 wl0_52
port 2102 nsew
rlabel metal2 s 21216 19403 21216 19403 4 wl0_47
port 2092 nsew
rlabel metal2 s 21216 17253 21216 17253 4 wl1_41
port 2081 nsew
rlabel metal2 s 21216 16243 21216 16243 4 wl0_39
port 2076 nsew
rlabel metal2 s 21216 19877 21216 19877 4 wl1_48
port 2095 nsew
rlabel metal2 s 21216 18613 21216 18613 4 wl0_45
port 2088 nsew
rlabel metal2 s 21216 22247 21216 22247 4 wl1_54
port 2107 nsew
rlabel metal2 s 21216 19087 21216 19087 4 wl1_46
port 2091 nsew
rlabel metal2 s 21216 25153 21216 25153 4 wl1_61
port 2121 nsew
rlabel metal2 s 21216 17727 21216 17727 4 wl0_42
port 2082 nsew
rlabel metal2 s 21216 15357 21216 15357 4 wl0_36
port 2070 nsew
rlabel metal2 s 21216 18833 21216 18833 4 wl1_45
port 2089 nsew
rlabel metal2 s 21216 25723 21216 25723 4 wl0_63
port 2124 nsew
rlabel metal2 s 21216 25943 21216 25943 4 wl1_63
port 2125 nsew
rlabel metal2 s 21216 15673 21216 15673 4 wl1_37
port 2073 nsew
rlabel metal2 s 21216 14663 21216 14663 4 wl0_35
port 2068 nsew
rlabel metal2 s 21216 15927 21216 15927 4 wl1_38
port 2075 nsew
rlabel metal2 s 21216 20887 21216 20887 4 wl0_50
port 2098 nsew
rlabel metal2 s 21216 25407 21216 25407 4 wl1_62
port 2123 nsew
rlabel metal2 s 21216 15137 21216 15137 4 wl1_36
port 2071 nsew
rlabel metal2 s 21216 20097 21216 20097 4 wl0_48
port 2094 nsew
rlabel metal2 s 21216 24047 21216 24047 4 wl0_58
port 2114 nsew
rlabel metal2 s 21216 21993 21216 21993 4 wl1_53
port 2105 nsew
rlabel metal2 s 21216 18517 21216 18517 4 wl0_44
port 2086 nsew
rlabel metal2 s 21216 22467 21216 22467 4 wl0_54
port 2106 nsew
rlabel metal2 s 21216 17507 21216 17507 4 wl1_42
port 2083 nsew
rlabel metal2 s 21216 19623 21216 19623 4 wl1_47
port 2093 nsew
rlabel metal2 s 21216 14347 21216 14347 4 wl1_34
port 2067 nsew
rlabel metal2 s 21216 22783 21216 22783 4 wl1_55
port 2109 nsew
rlabel metal2 s 21216 13303 21216 13303 4 wl1_31
port 2061 nsew
rlabel metal2 s 21216 20193 21216 20193 4 wl0_49
port 2096 nsew
rlabel metal2 s 21216 13873 21216 13873 4 wl0_33
port 2064 nsew
rlabel metal2 s 21216 17823 21216 17823 4 wl0_43
port 2084 nsew
rlabel metal2 s 21216 23573 21216 23573 4 wl1_57
port 2113 nsew
rlabel metal2 s 21216 15453 21216 15453 4 wl0_37
port 2072 nsew
rlabel metal2 s 21216 23037 21216 23037 4 wl1_56
port 2111 nsew
rlabel metal2 s 21216 24933 21216 24933 4 wl0_61
port 2120 nsew
rlabel metal2 s 21216 24363 21216 24363 4 wl1_59
port 2117 nsew
rlabel metal2 s 21216 16937 21216 16937 4 wl0_40
port 2078 nsew
rlabel metal2 s 21216 17033 21216 17033 4 wl0_41
port 2080 nsew
rlabel metal2 s 21216 18297 21216 18297 4 wl1_44
port 2087 nsew
rlabel metal2 s 21216 25627 21216 25627 4 wl0_62
port 2122 nsew
rlabel metal2 s 21216 23827 21216 23827 4 wl1_58
port 2115 nsew
rlabel metal2 s 21216 14567 21216 14567 4 wl0_34
port 2066 nsew
rlabel metal2 s 21216 20413 21216 20413 4 wl1_49
port 2097 nsew
rlabel metal2 s 21216 24143 21216 24143 4 wl0_59
port 2116 nsew
rlabel metal2 s 21216 14883 21216 14883 4 wl1_35
port 2069 nsew
rlabel metal2 s 21216 21773 21216 21773 4 wl0_53
port 2104 nsew
rlabel metal2 s 1008 16590 1008 16590 4 gnd
port 2 nsew
rlabel metal2 s 1008 18170 1008 18170 4 gnd
port 2 nsew
rlabel metal2 s 1008 24490 1008 24490 4 gnd
port 2 nsew
rlabel metal2 s 1008 19197 1008 19197 4 gnd
port 2 nsew
rlabel metal2 s 1008 21330 1008 21330 4 gnd
port 2 nsew
rlabel metal2 s 1008 20777 1008 20777 4 gnd
port 2 nsew
rlabel metal2 s 1008 20540 1008 20540 4 gnd
port 2 nsew
rlabel metal2 s 1008 19513 1008 19513 4 gnd
port 2 nsew
rlabel metal2 s 1008 15563 1008 15563 4 gnd
port 2 nsew
rlabel metal2 s 1008 23700 1008 23700 4 gnd
port 2 nsew
rlabel metal2 s 1008 25517 1008 25517 4 gnd
port 2 nsew
rlabel metal2 s 1008 16827 1008 16827 4 gnd
port 2 nsew
rlabel metal2 s 1008 22910 1008 22910 4 gnd
port 2 nsew
rlabel metal2 s 1008 14220 1008 14220 4 gnd
port 2 nsew
rlabel metal2 s 1008 16037 1008 16037 4 gnd
port 2 nsew
rlabel metal2 s 1008 18723 1008 18723 4 gnd
port 2 nsew
rlabel metal2 s 1008 23463 1008 23463 4 gnd
port 2 nsew
rlabel metal2 s 1008 21883 1008 21883 4 gnd
port 2 nsew
rlabel metal2 s 1008 18407 1008 18407 4 gnd
port 2 nsew
rlabel metal2 s 1008 17380 1008 17380 4 gnd
port 2 nsew
rlabel metal2 s 1008 14773 1008 14773 4 gnd
port 2 nsew
rlabel metal2 s 1008 22120 1008 22120 4 gnd
port 2 nsew
rlabel metal2 s 1008 24253 1008 24253 4 gnd
port 2 nsew
rlabel metal2 s 1008 22357 1008 22357 4 gnd
port 2 nsew
rlabel metal2 s 1008 16353 1008 16353 4 gnd
port 2 nsew
rlabel metal2 s 1008 13430 1008 13430 4 gnd
port 2 nsew
rlabel metal2 s 1008 23937 1008 23937 4 gnd
port 2 nsew
rlabel metal2 s 1008 22673 1008 22673 4 gnd
port 2 nsew
rlabel metal2 s 1008 25280 1008 25280 4 gnd
port 2 nsew
rlabel metal2 s 1008 17617 1008 17617 4 gnd
port 2 nsew
rlabel metal2 s 1008 15010 1008 15010 4 gnd
port 2 nsew
rlabel metal2 s 1008 25043 1008 25043 4 gnd
port 2 nsew
rlabel metal2 s 1008 24727 1008 24727 4 gnd
port 2 nsew
rlabel metal2 s 1008 13983 1008 13983 4 gnd
port 2 nsew
rlabel metal2 s 1008 21093 1008 21093 4 gnd
port 2 nsew
rlabel metal2 s 1008 18960 1008 18960 4 gnd
port 2 nsew
rlabel metal2 s 1008 15800 1008 15800 4 gnd
port 2 nsew
rlabel metal2 s 1008 17933 1008 17933 4 gnd
port 2 nsew
rlabel metal2 s 1008 23147 1008 23147 4 gnd
port 2 nsew
rlabel metal2 s 1008 25833 1008 25833 4 gnd
port 2 nsew
rlabel metal2 s 1008 20303 1008 20303 4 gnd
port 2 nsew
rlabel metal2 s 1008 19750 1008 19750 4 gnd
port 2 nsew
rlabel metal2 s 1008 17143 1008 17143 4 gnd
port 2 nsew
rlabel metal2 s 1008 21567 1008 21567 4 gnd
port 2 nsew
rlabel metal2 s 1008 15247 1008 15247 4 gnd
port 2 nsew
rlabel metal2 s 1008 19987 1008 19987 4 gnd
port 2 nsew
rlabel metal2 s 1008 13667 1008 13667 4 gnd
port 2 nsew
rlabel metal2 s 1008 14457 1008 14457 4 gnd
port 2 nsew
rlabel metal2 s 1008 9243 1008 9243 4 gnd
port 2 nsew
rlabel metal2 s 1008 10270 1008 10270 4 gnd
port 2 nsew
rlabel metal2 s 1008 7110 1008 7110 4 gnd
port 2 nsew
rlabel metal2 s 1008 3160 1008 3160 4 gnd
port 2 nsew
rlabel metal2 s 1008 6557 1008 6557 4 gnd
port 2 nsew
rlabel metal2 s 1008 6320 1008 6320 4 gnd
port 2 nsew
rlabel metal2 s 1008 790 1008 790 4 gnd
port 2 nsew
rlabel metal2 s 1008 5293 1008 5293 4 gnd
port 2 nsew
rlabel metal2 s 1008 10823 1008 10823 4 gnd
port 2 nsew
rlabel metal2 s 1008 5767 1008 5767 4 gnd
port 2 nsew
rlabel metal2 s 1008 12087 1008 12087 4 gnd
port 2 nsew
rlabel metal2 s 1008 3713 1008 3713 4 gnd
port 2 nsew
rlabel metal2 s 1008 8453 1008 8453 4 gnd
port 2 nsew
rlabel metal2 s 1008 6083 1008 6083 4 gnd
port 2 nsew
rlabel metal2 s 1008 10033 1008 10033 4 gnd
port 2 nsew
rlabel metal2 s 1008 4740 1008 4740 4 gnd
port 2 nsew
rlabel metal2 s 1008 3950 1008 3950 4 gnd
port 2 nsew
rlabel metal2 s 1008 11850 1008 11850 4 gnd
port 2 nsew
rlabel metal2 s 1008 8137 1008 8137 4 gnd
port 2 nsew
rlabel metal2 s 1008 7663 1008 7663 4 gnd
port 2 nsew
rlabel metal2 s 1008 12640 1008 12640 4 gnd
port 2 nsew
rlabel metal2 s 1008 1027 1008 1027 4 gnd
port 2 nsew
rlabel metal2 s 1008 11297 1008 11297 4 gnd
port 2 nsew
rlabel metal2 s 1008 8690 1008 8690 4 gnd
port 2 nsew
rlabel metal2 s 1008 11060 1008 11060 4 gnd
port 2 nsew
rlabel metal2 s 1008 12877 1008 12877 4 gnd
port 2 nsew
rlabel metal2 s 1008 7347 1008 7347 4 gnd
port 2 nsew
rlabel metal2 s 1008 8927 1008 8927 4 gnd
port 2 nsew
rlabel metal2 s 1008 6873 1008 6873 4 gnd
port 2 nsew
rlabel metal2 s 1008 12403 1008 12403 4 gnd
port 2 nsew
rlabel metal2 s 1008 5530 1008 5530 4 gnd
port 2 nsew
rlabel metal2 s 1008 1343 1008 1343 4 gnd
port 2 nsew
rlabel metal2 s 1008 2133 1008 2133 4 gnd
port 2 nsew
rlabel metal2 s 1008 7900 1008 7900 4 gnd
port 2 nsew
rlabel metal2 s 1008 13193 1008 13193 4 gnd
port 2 nsew
rlabel metal2 s 1008 2370 1008 2370 4 gnd
port 2 nsew
rlabel metal2 s 1008 2923 1008 2923 4 gnd
port 2 nsew
rlabel metal2 s 1008 2607 1008 2607 4 gnd
port 2 nsew
rlabel metal2 s 1008 4187 1008 4187 4 gnd
port 2 nsew
rlabel metal2 s 1008 1580 1008 1580 4 gnd
port 2 nsew
rlabel metal2 s 1008 1817 1008 1817 4 gnd
port 2 nsew
rlabel metal2 s 1008 3397 1008 3397 4 gnd
port 2 nsew
rlabel metal2 s 1008 9480 1008 9480 4 gnd
port 2 nsew
rlabel metal2 s 1008 11613 1008 11613 4 gnd
port 2 nsew
rlabel metal2 s 1008 4503 1008 4503 4 gnd
port 2 nsew
rlabel metal2 s 1008 4977 1008 4977 4 gnd
port 2 nsew
rlabel metal2 s 1008 9717 1008 9717 4 gnd
port 2 nsew
rlabel metal2 s 1008 10507 1008 10507 4 gnd
port 2 nsew
rlabel metal2 s 1008 553 1008 553 4 gnd
port 2 nsew
rlabel metal2 s 21216 11723 21216 11723 4 wl1_27
port 2053 nsew
rlabel metal2 s 21216 1707 21216 1707 4 wl1_2
port 2003 nsew
rlabel metal2 s 21216 10713 21216 10713 4 wl0_25
port 2048 nsew
rlabel metal2 s 21216 5973 21216 5973 4 wl0_13
port 2024 nsew
rlabel metal2 s 21216 5403 21216 5403 4 wl1_11
port 2021 nsew
rlabel metal2 s 21216 6983 21216 6983 4 wl1_15
port 2029 nsew
rlabel metal2 s 21216 10617 21216 10617 4 wl0_24
port 2046 nsew
rlabel metal2 s 21216 11407 21216 11407 4 wl0_26
port 2050 nsew
rlabel metal2 s 21216 3603 21216 3603 4 wl0_7
port 2012 nsew
rlabel metal2 s 21216 6193 21216 6193 4 wl1_13
port 2025 nsew
rlabel metal2 s 21216 9353 21216 9353 4 wl1_21
port 2041 nsew
rlabel metal2 s 21216 9037 21216 9037 4 wl0_20
port 2038 nsew
rlabel metal2 s 21216 1453 21216 1453 4 wl1_1
port 2001 nsew
rlabel metal2 s 21216 11977 21216 11977 4 wl1_28
port 2055 nsew
rlabel metal2 s 21216 2717 21216 2717 4 wl0_4
port 2006 nsew
rlabel metal2 s 21216 11503 21216 11503 4 wl0_27
port 2052 nsew
rlabel metal2 s 21216 3287 21216 3287 4 wl1_6
port 2011 nsew
rlabel metal2 s 21216 12987 21216 12987 4 wl0_30
port 2058 nsew
rlabel metal2 s 21216 12293 21216 12293 4 wl0_29
port 2056 nsew
rlabel metal2 s 21216 5877 21216 5877 4 wl0_12
port 2022 nsew
rlabel metal2 s 21216 11187 21216 11187 4 wl1_26
port 2051 nsew
rlabel metal2 s 21216 13083 21216 13083 4 wl0_31
port 2060 nsew
rlabel metal2 s 21216 2243 21216 2243 4 wl1_3
port 2005 nsew
rlabel metal2 s 21216 443 21216 443 4 rbl_wl0_0
port 2254 nsew
rlabel metal2 s 21216 8343 21216 8343 4 wl0_19
port 2036 nsew
rlabel metal2 s 21216 12197 21216 12197 4 wl0_28
port 2054 nsew
rlabel metal2 s 21216 12513 21216 12513 4 wl1_29
port 2057 nsew
rlabel metal2 s 21216 2813 21216 2813 4 wl0_5
port 2008 nsew
rlabel metal2 s 21216 1137 21216 1137 4 wl0_0
port 1998 nsew
rlabel metal2 s 21216 3033 21216 3033 4 wl1_5
port 2009 nsew
rlabel metal2 s 21216 10397 21216 10397 4 wl1_24
port 2047 nsew
rlabel metal2 s 21216 9923 21216 9923 4 wl0_23
port 2044 nsew
rlabel metal2 s 21216 7237 21216 7237 4 wl1_16
port 2031 nsew
rlabel metal2 s 21216 2497 21216 2497 4 wl1_4
port 2007 nsew
rlabel metal2 s 21216 5183 21216 5183 4 wl0_11
port 2020 nsew
rlabel metal2 s 21216 1927 21216 1927 4 wl0_2
port 2002 nsew
rlabel metal2 s 21216 4393 21216 4393 4 wl0_9
port 2016 nsew
rlabel metal2 s 21216 917 21216 917 4 wl1_0
port 1999 nsew
rlabel metal2 s 21216 7773 21216 7773 4 wl1_17
port 2033 nsew
rlabel metal2 s 21216 12767 21216 12767 4 wl1_30
port 2059 nsew
rlabel metal2 s 21216 1233 21216 1233 4 wl0_1
port 2000 nsew
rlabel metal2 s 21216 8563 21216 8563 4 wl1_19
port 2037 nsew
rlabel metal2 s 21216 2023 21216 2023 4 wl0_3
port 2004 nsew
rlabel metal2 s 21216 10933 21216 10933 4 wl1_25
port 2049 nsew
rlabel metal2 s 21216 3823 21216 3823 4 wl1_7
port 2013 nsew
rlabel metal2 s 21216 8027 21216 8027 4 wl1_18
port 2035 nsew
rlabel metal2 s 21216 6667 21216 6667 4 wl0_14
port 2026 nsew
rlabel metal2 s 21216 6447 21216 6447 4 wl1_14
port 2027 nsew
rlabel metal2 s 21216 4297 21216 4297 4 wl0_8
port 2014 nsew
rlabel metal2 s 21216 5087 21216 5087 4 wl0_10
port 2018 nsew
rlabel metal2 s 21216 7553 21216 7553 4 wl0_17
port 2032 nsew
rlabel metal2 s 21216 10143 21216 10143 4 wl1_23
port 2045 nsew
rlabel metal2 s 21216 3507 21216 3507 4 wl0_6
port 2010 nsew
rlabel metal2 s 21216 8247 21216 8247 4 wl0_18
port 2034 nsew
rlabel metal2 s 21216 8817 21216 8817 4 wl1_20
port 2039 nsew
rlabel metal2 s 21216 7457 21216 7457 4 wl0_16
port 2030 nsew
rlabel metal2 s 21216 5657 21216 5657 4 wl1_12
port 2023 nsew
rlabel metal2 s 21216 4867 21216 4867 4 wl1_10
port 2019 nsew
rlabel metal2 s 21216 9827 21216 9827 4 wl0_22
port 2042 nsew
rlabel metal2 s 21216 4613 21216 4613 4 wl1_9
port 2017 nsew
rlabel metal2 s 21216 6763 21216 6763 4 wl0_15
port 2028 nsew
rlabel metal2 s 21216 9607 21216 9607 4 wl1_22
port 2043 nsew
rlabel metal2 s 21216 9133 21216 9133 4 wl0_21
port 2040 nsew
rlabel metal2 s 21216 4077 21216 4077 4 wl1_8
port 2015 nsew
rlabel metal2 s 41424 23937 41424 23937 4 gnd
port 2 nsew
rlabel metal2 s 41424 21330 41424 21330 4 gnd
port 2 nsew
rlabel metal2 s 41424 15247 41424 15247 4 gnd
port 2 nsew
rlabel metal2 s 41424 13193 41424 13193 4 gnd
port 2 nsew
rlabel metal2 s 41424 5530 41424 5530 4 gnd
port 2 nsew
rlabel metal2 s 41424 24490 41424 24490 4 gnd
port 2 nsew
rlabel metal2 s 41424 5293 41424 5293 4 gnd
port 2 nsew
rlabel metal2 s 41424 20540 41424 20540 4 gnd
port 2 nsew
rlabel metal2 s 41424 23147 41424 23147 4 gnd
port 2 nsew
rlabel metal2 s 41424 553 41424 553 4 gnd
port 2 nsew
rlabel metal2 s 41424 3397 41424 3397 4 gnd
port 2 nsew
rlabel metal2 s 41424 17143 41424 17143 4 gnd
port 2 nsew
rlabel metal2 s 41424 14220 41424 14220 4 gnd
port 2 nsew
rlabel metal2 s 41424 24253 41424 24253 4 gnd
port 2 nsew
rlabel metal2 s 41424 7110 41424 7110 4 gnd
port 2 nsew
rlabel metal2 s 41424 14773 41424 14773 4 gnd
port 2 nsew
rlabel metal2 s 41424 4977 41424 4977 4 gnd
port 2 nsew
rlabel metal2 s 41424 11060 41424 11060 4 gnd
port 2 nsew
rlabel metal2 s 41424 1027 41424 1027 4 gnd
port 2 nsew
rlabel metal2 s 41424 8453 41424 8453 4 gnd
port 2 nsew
rlabel metal2 s 41424 17617 41424 17617 4 gnd
port 2 nsew
rlabel metal2 s 41424 16827 41424 16827 4 gnd
port 2 nsew
rlabel metal2 s 41424 19513 41424 19513 4 gnd
port 2 nsew
rlabel metal2 s 41424 1817 41424 1817 4 gnd
port 2 nsew
rlabel metal2 s 41424 5767 41424 5767 4 gnd
port 2 nsew
rlabel metal2 s 41424 18960 41424 18960 4 gnd
port 2 nsew
rlabel metal2 s 41424 10823 41424 10823 4 gnd
port 2 nsew
rlabel metal2 s 41424 7347 41424 7347 4 gnd
port 2 nsew
rlabel metal2 s 41424 15010 41424 15010 4 gnd
port 2 nsew
rlabel metal2 s 41424 10507 41424 10507 4 gnd
port 2 nsew
rlabel metal2 s 41424 2923 41424 2923 4 gnd
port 2 nsew
rlabel metal2 s 41424 12403 41424 12403 4 gnd
port 2 nsew
rlabel metal2 s 41424 20777 41424 20777 4 gnd
port 2 nsew
rlabel metal2 s 41424 21567 41424 21567 4 gnd
port 2 nsew
rlabel metal2 s 41424 13667 41424 13667 4 gnd
port 2 nsew
rlabel metal2 s 41424 18407 41424 18407 4 gnd
port 2 nsew
rlabel metal2 s 41424 3713 41424 3713 4 gnd
port 2 nsew
rlabel metal2 s 41424 1580 41424 1580 4 gnd
port 2 nsew
rlabel metal2 s 41424 18723 41424 18723 4 gnd
port 2 nsew
rlabel metal2 s 41424 25280 41424 25280 4 gnd
port 2 nsew
rlabel metal2 s 41424 22120 41424 22120 4 gnd
port 2 nsew
rlabel metal2 s 41424 8927 41424 8927 4 gnd
port 2 nsew
rlabel metal2 s 41424 12877 41424 12877 4 gnd
port 2 nsew
rlabel metal2 s 41424 9717 41424 9717 4 gnd
port 2 nsew
rlabel metal2 s 41424 23463 41424 23463 4 gnd
port 2 nsew
rlabel metal2 s 41424 20303 41424 20303 4 gnd
port 2 nsew
rlabel metal2 s 41424 17933 41424 17933 4 gnd
port 2 nsew
rlabel metal2 s 41424 11850 41424 11850 4 gnd
port 2 nsew
rlabel metal2 s 41424 22673 41424 22673 4 gnd
port 2 nsew
rlabel metal2 s 41424 15800 41424 15800 4 gnd
port 2 nsew
rlabel metal2 s 41424 22910 41424 22910 4 gnd
port 2 nsew
rlabel metal2 s 41424 16037 41424 16037 4 gnd
port 2 nsew
rlabel metal2 s 41424 6320 41424 6320 4 gnd
port 2 nsew
rlabel metal2 s 41424 19987 41424 19987 4 gnd
port 2 nsew
rlabel metal2 s 41424 6557 41424 6557 4 gnd
port 2 nsew
rlabel metal2 s 41424 3160 41424 3160 4 gnd
port 2 nsew
rlabel metal2 s 41424 22357 41424 22357 4 gnd
port 2 nsew
rlabel metal2 s 41424 19197 41424 19197 4 gnd
port 2 nsew
rlabel metal2 s 41424 25043 41424 25043 4 gnd
port 2 nsew
rlabel metal2 s 41424 12087 41424 12087 4 gnd
port 2 nsew
rlabel metal2 s 41424 16353 41424 16353 4 gnd
port 2 nsew
rlabel metal2 s 41424 23700 41424 23700 4 gnd
port 2 nsew
rlabel metal2 s 41424 6873 41424 6873 4 gnd
port 2 nsew
rlabel metal2 s 41424 4740 41424 4740 4 gnd
port 2 nsew
rlabel metal2 s 41424 18170 41424 18170 4 gnd
port 2 nsew
rlabel metal2 s 41424 14457 41424 14457 4 gnd
port 2 nsew
rlabel metal2 s 41424 13983 41424 13983 4 gnd
port 2 nsew
rlabel metal2 s 41424 6083 41424 6083 4 gnd
port 2 nsew
rlabel metal2 s 41424 16590 41424 16590 4 gnd
port 2 nsew
rlabel metal2 s 41424 15563 41424 15563 4 gnd
port 2 nsew
rlabel metal2 s 41424 21093 41424 21093 4 gnd
port 2 nsew
rlabel metal2 s 41424 17380 41424 17380 4 gnd
port 2 nsew
rlabel metal2 s 41424 8690 41424 8690 4 gnd
port 2 nsew
rlabel metal2 s 41424 10033 41424 10033 4 gnd
port 2 nsew
rlabel metal2 s 41424 10270 41424 10270 4 gnd
port 2 nsew
rlabel metal2 s 41424 3950 41424 3950 4 gnd
port 2 nsew
rlabel metal2 s 41424 21883 41424 21883 4 gnd
port 2 nsew
rlabel metal2 s 41424 2370 41424 2370 4 gnd
port 2 nsew
rlabel metal2 s 41424 2133 41424 2133 4 gnd
port 2 nsew
rlabel metal2 s 41424 7663 41424 7663 4 gnd
port 2 nsew
rlabel metal2 s 41424 4187 41424 4187 4 gnd
port 2 nsew
rlabel metal2 s 41424 11613 41424 11613 4 gnd
port 2 nsew
rlabel metal2 s 41424 7900 41424 7900 4 gnd
port 2 nsew
rlabel metal2 s 41424 2607 41424 2607 4 gnd
port 2 nsew
rlabel metal2 s 41424 19750 41424 19750 4 gnd
port 2 nsew
rlabel metal2 s 41424 13430 41424 13430 4 gnd
port 2 nsew
rlabel metal2 s 41424 25517 41424 25517 4 gnd
port 2 nsew
rlabel metal2 s 41424 9480 41424 9480 4 gnd
port 2 nsew
rlabel metal2 s 41424 790 41424 790 4 gnd
port 2 nsew
rlabel metal2 s 41424 12640 41424 12640 4 gnd
port 2 nsew
rlabel metal2 s 41424 24727 41424 24727 4 gnd
port 2 nsew
rlabel metal2 s 41424 25833 41424 25833 4 gnd
port 2 nsew
rlabel metal2 s 41424 9243 41424 9243 4 gnd
port 2 nsew
rlabel metal2 s 41424 1343 41424 1343 4 gnd
port 2 nsew
rlabel metal2 s 41424 8137 41424 8137 4 gnd
port 2 nsew
rlabel metal2 s 41424 4503 41424 4503 4 gnd
port 2 nsew
rlabel metal2 s 41424 11297 41424 11297 4 gnd
port 2 nsew
rlabel metal3 s 42192 44793 42192 44793 4 gnd
port 2 nsew
rlabel metal3 s 42192 44477 42192 44477 4 gnd
port 2 nsew
rlabel metal3 s 42192 40527 42192 40527 4 gnd
port 2 nsew
rlabel metal3 s 42192 47400 42192 47400 4 gnd
port 2 nsew
rlabel metal3 s 42192 42897 42192 42897 4 gnd
port 2 nsew
rlabel metal3 s 42192 44240 42192 44240 4 gnd
port 2 nsew
rlabel metal3 s 42192 41080 42192 41080 4 gnd
port 2 nsew
rlabel metal3 s 42192 44003 42192 44003 4 gnd
port 2 nsew
rlabel metal3 s 42192 45820 42192 45820 4 gnd
port 2 nsew
rlabel metal3 s 42192 39737 42192 39737 4 gnd
port 2 nsew
rlabel metal3 s 42192 46610 42192 46610 4 gnd
port 2 nsew
rlabel metal3 s 42192 47953 42192 47953 4 gnd
port 2 nsew
rlabel metal3 s 42192 48427 42192 48427 4 gnd
port 2 nsew
rlabel metal3 s 42192 43450 42192 43450 4 gnd
port 2 nsew
rlabel metal3 s 42192 51587 42192 51587 4 gnd
port 2 nsew
rlabel metal3 s 42192 48190 42192 48190 4 gnd
port 2 nsew
rlabel metal3 s 42192 41633 42192 41633 4 gnd
port 2 nsew
rlabel metal3 s 42192 47637 42192 47637 4 gnd
port 2 nsew
rlabel metal3 s 42192 39500 42192 39500 4 gnd
port 2 nsew
rlabel metal3 s 42192 49770 42192 49770 4 gnd
port 2 nsew
rlabel metal3 s 42192 40843 42192 40843 4 gnd
port 2 nsew
rlabel metal3 s 42192 51350 42192 51350 4 gnd
port 2 nsew
rlabel metal3 s 42192 48743 42192 48743 4 gnd
port 2 nsew
rlabel metal3 s 42192 41870 42192 41870 4 gnd
port 2 nsew
rlabel metal3 s 42192 40053 42192 40053 4 gnd
port 2 nsew
rlabel metal3 s 42192 50797 42192 50797 4 gnd
port 2 nsew
rlabel metal3 s 42192 50007 42192 50007 4 gnd
port 2 nsew
rlabel metal3 s 42192 42660 42192 42660 4 gnd
port 2 nsew
rlabel metal3 s 42192 48980 42192 48980 4 gnd
port 2 nsew
rlabel metal3 s 42192 45030 42192 45030 4 gnd
port 2 nsew
rlabel metal3 s 42192 49217 42192 49217 4 gnd
port 2 nsew
rlabel metal3 s 42192 42423 42192 42423 4 gnd
port 2 nsew
rlabel metal3 s 42192 45267 42192 45267 4 gnd
port 2 nsew
rlabel metal3 s 42192 41317 42192 41317 4 gnd
port 2 nsew
rlabel metal3 s 42192 42107 42192 42107 4 gnd
port 2 nsew
rlabel metal3 s 42192 47163 42192 47163 4 gnd
port 2 nsew
rlabel metal3 s 42192 46373 42192 46373 4 gnd
port 2 nsew
rlabel metal3 s 42192 39263 42192 39263 4 gnd
port 2 nsew
rlabel metal3 s 42192 40290 42192 40290 4 gnd
port 2 nsew
rlabel metal3 s 42192 51113 42192 51113 4 gnd
port 2 nsew
rlabel metal3 s 42192 46847 42192 46847 4 gnd
port 2 nsew
rlabel metal3 s 42192 43213 42192 43213 4 gnd
port 2 nsew
rlabel metal3 s 42192 45583 42192 45583 4 gnd
port 2 nsew
rlabel metal3 s 42192 43687 42192 43687 4 gnd
port 2 nsew
rlabel metal3 s 42192 49533 42192 49533 4 gnd
port 2 nsew
rlabel metal3 s 42192 46057 42192 46057 4 gnd
port 2 nsew
rlabel metal3 s 42192 50560 42192 50560 4 gnd
port 2 nsew
rlabel metal3 s 42192 50323 42192 50323 4 gnd
port 2 nsew
rlabel metal3 s 34632 51911 34632 51911 4 vdd
port 1 nsew
rlabel metal3 s 39000 51911 39000 51911 4 vdd
port 1 nsew
rlabel metal3 s 41496 51911 41496 51911 4 vdd
port 1 nsew
rlabel metal3 s 37752 51911 37752 51911 4 vdd
port 1 nsew
rlabel metal3 s 37128 51911 37128 51911 4 vdd
port 1 nsew
rlabel metal3 s 36504 51911 36504 51911 4 vdd
port 1 nsew
rlabel metal3 s 35256 51911 35256 51911 4 vdd
port 1 nsew
rlabel metal3 s 32136 51911 32136 51911 4 vdd
port 1 nsew
rlabel metal3 s 35880 51911 35880 51911 4 vdd
port 1 nsew
rlabel metal3 s 39624 51911 39624 51911 4 vdd
port 1 nsew
rlabel metal3 s 40248 51911 40248 51911 4 vdd
port 1 nsew
rlabel metal3 s 32760 51911 32760 51911 4 vdd
port 1 nsew
rlabel metal3 s 38376 51911 38376 51911 4 vdd
port 1 nsew
rlabel metal3 s 33384 51911 33384 51911 4 vdd
port 1 nsew
rlabel metal3 s 34008 51911 34008 51911 4 vdd
port 1 nsew
rlabel metal3 s 40872 51911 40872 51911 4 vdd
port 1 nsew
rlabel metal3 s 30264 51911 30264 51911 4 vdd
port 1 nsew
rlabel metal3 s 24648 51911 24648 51911 4 vdd
port 1 nsew
rlabel metal3 s 25896 51911 25896 51911 4 vdd
port 1 nsew
rlabel metal3 s 23400 51911 23400 51911 4 vdd
port 1 nsew
rlabel metal3 s 30888 51911 30888 51911 4 vdd
port 1 nsew
rlabel metal3 s 25272 51911 25272 51911 4 vdd
port 1 nsew
rlabel metal3 s 28392 51911 28392 51911 4 vdd
port 1 nsew
rlabel metal3 s 29640 51911 29640 51911 4 vdd
port 1 nsew
rlabel metal3 s 22152 51911 22152 51911 4 vdd
port 1 nsew
rlabel metal3 s 27768 51911 27768 51911 4 vdd
port 1 nsew
rlabel metal3 s 29016 51911 29016 51911 4 vdd
port 1 nsew
rlabel metal3 s 26520 51911 26520 51911 4 vdd
port 1 nsew
rlabel metal3 s 24024 51911 24024 51911 4 vdd
port 1 nsew
rlabel metal3 s 21528 51911 21528 51911 4 vdd
port 1 nsew
rlabel metal3 s 27144 51911 27144 51911 4 vdd
port 1 nsew
rlabel metal3 s 22776 51911 22776 51911 4 vdd
port 1 nsew
rlabel metal3 s 31512 51911 31512 51911 4 vdd
port 1 nsew
rlabel metal3 s 42192 29783 42192 29783 4 gnd
port 2 nsew
rlabel metal3 s 42192 30020 42192 30020 4 gnd
port 2 nsew
rlabel metal3 s 42192 30257 42192 30257 4 gnd
port 2 nsew
rlabel metal3 s 42192 37683 42192 37683 4 gnd
port 2 nsew
rlabel metal3 s 42192 32627 42192 32627 4 gnd
port 2 nsew
rlabel metal3 s 42192 30573 42192 30573 4 gnd
port 2 nsew
rlabel metal3 s 42192 36103 42192 36103 4 gnd
port 2 nsew
rlabel metal3 s 42192 37367 42192 37367 4 gnd
port 2 nsew
rlabel metal3 s 42192 28993 42192 28993 4 gnd
port 2 nsew
rlabel metal3 s 42192 36340 42192 36340 4 gnd
port 2 nsew
rlabel metal3 s 42192 38710 42192 38710 4 gnd
port 2 nsew
rlabel metal3 s 42192 29230 42192 29230 4 gnd
port 2 nsew
rlabel metal3 s 42192 34997 42192 34997 4 gnd
port 2 nsew
rlabel metal3 s 42192 32153 42192 32153 4 gnd
port 2 nsew
rlabel metal3 s 42192 26623 42192 26623 4 gnd
port 2 nsew
rlabel metal3 s 42192 38157 42192 38157 4 gnd
port 2 nsew
rlabel metal3 s 42192 29467 42192 29467 4 gnd
port 2 nsew
rlabel metal3 s 42192 33733 42192 33733 4 gnd
port 2 nsew
rlabel metal3 s 42192 32390 42192 32390 4 gnd
port 2 nsew
rlabel metal3 s 42192 38473 42192 38473 4 gnd
port 2 nsew
rlabel metal3 s 42192 27097 42192 27097 4 gnd
port 2 nsew
rlabel metal3 s 42192 31363 42192 31363 4 gnd
port 2 nsew
rlabel metal3 s 42192 34523 42192 34523 4 gnd
port 2 nsew
rlabel metal3 s 42192 34760 42192 34760 4 gnd
port 2 nsew
rlabel metal3 s 42192 31047 42192 31047 4 gnd
port 2 nsew
rlabel metal3 s 42192 34207 42192 34207 4 gnd
port 2 nsew
rlabel metal3 s 42192 37920 42192 37920 4 gnd
port 2 nsew
rlabel metal3 s 42192 37130 42192 37130 4 gnd
port 2 nsew
rlabel metal3 s 42192 35313 42192 35313 4 gnd
port 2 nsew
rlabel metal3 s 42192 35787 42192 35787 4 gnd
port 2 nsew
rlabel metal3 s 42192 30810 42192 30810 4 gnd
port 2 nsew
rlabel metal3 s 42192 32943 42192 32943 4 gnd
port 2 nsew
rlabel metal3 s 42192 27413 42192 27413 4 gnd
port 2 nsew
rlabel metal3 s 42192 33180 42192 33180 4 gnd
port 2 nsew
rlabel metal3 s 42192 28677 42192 28677 4 gnd
port 2 nsew
rlabel metal3 s 42192 27650 42192 27650 4 gnd
port 2 nsew
rlabel metal3 s 42192 35550 42192 35550 4 gnd
port 2 nsew
rlabel metal3 s 42192 36577 42192 36577 4 gnd
port 2 nsew
rlabel metal3 s 42192 38947 42192 38947 4 gnd
port 2 nsew
rlabel metal3 s 42192 28203 42192 28203 4 gnd
port 2 nsew
rlabel metal3 s 42192 31600 42192 31600 4 gnd
port 2 nsew
rlabel metal3 s 42192 26307 42192 26307 4 gnd
port 2 nsew
rlabel metal3 s 42192 27887 42192 27887 4 gnd
port 2 nsew
rlabel metal3 s 42192 26860 42192 26860 4 gnd
port 2 nsew
rlabel metal3 s 42192 28440 42192 28440 4 gnd
port 2 nsew
rlabel metal3 s 42192 36893 42192 36893 4 gnd
port 2 nsew
rlabel metal3 s 42192 31837 42192 31837 4 gnd
port 2 nsew
rlabel metal3 s 42192 33970 42192 33970 4 gnd
port 2 nsew
rlabel metal3 s 42192 33417 42192 33417 4 gnd
port 2 nsew
rlabel metal3 s 17784 51911 17784 51911 4 vdd
port 1 nsew
rlabel metal3 s 13416 51911 13416 51911 4 vdd
port 1 nsew
rlabel metal3 s 19032 51911 19032 51911 4 vdd
port 1 nsew
rlabel metal3 s 20904 51911 20904 51911 4 vdd
port 1 nsew
rlabel metal3 s 20280 51911 20280 51911 4 vdd
port 1 nsew
rlabel metal3 s 18408 51911 18408 51911 4 vdd
port 1 nsew
rlabel metal3 s 15912 51911 15912 51911 4 vdd
port 1 nsew
rlabel metal3 s 16536 51911 16536 51911 4 vdd
port 1 nsew
rlabel metal3 s 14040 51911 14040 51911 4 vdd
port 1 nsew
rlabel metal3 s 14664 51911 14664 51911 4 vdd
port 1 nsew
rlabel metal3 s 12792 51911 12792 51911 4 vdd
port 1 nsew
rlabel metal3 s 15288 51911 15288 51911 4 vdd
port 1 nsew
rlabel metal3 s 19656 51911 19656 51911 4 vdd
port 1 nsew
rlabel metal3 s 11544 51911 11544 51911 4 vdd
port 1 nsew
rlabel metal3 s 17160 51911 17160 51911 4 vdd
port 1 nsew
rlabel metal3 s 12168 51911 12168 51911 4 vdd
port 1 nsew
rlabel metal3 s 10920 51911 10920 51911 4 vdd
port 1 nsew
rlabel metal3 s 240 40290 240 40290 4 gnd
port 2 nsew
rlabel metal3 s 240 44003 240 44003 4 gnd
port 2 nsew
rlabel metal3 s 240 49533 240 49533 4 gnd
port 2 nsew
rlabel metal3 s 240 47953 240 47953 4 gnd
port 2 nsew
rlabel metal3 s 240 46847 240 46847 4 gnd
port 2 nsew
rlabel metal3 s 240 43213 240 43213 4 gnd
port 2 nsew
rlabel metal3 s 240 46373 240 46373 4 gnd
port 2 nsew
rlabel metal3 s 240 45030 240 45030 4 gnd
port 2 nsew
rlabel metal3 s 240 39737 240 39737 4 gnd
port 2 nsew
rlabel metal3 s 240 44793 240 44793 4 gnd
port 2 nsew
rlabel metal3 s 240 50797 240 50797 4 gnd
port 2 nsew
rlabel metal3 s 240 49217 240 49217 4 gnd
port 2 nsew
rlabel metal3 s 240 46057 240 46057 4 gnd
port 2 nsew
rlabel metal3 s 240 51350 240 51350 4 gnd
port 2 nsew
rlabel metal3 s 240 51113 240 51113 4 gnd
port 2 nsew
rlabel metal3 s 240 50323 240 50323 4 gnd
port 2 nsew
rlabel metal3 s 240 39500 240 39500 4 gnd
port 2 nsew
rlabel metal3 s 240 47163 240 47163 4 gnd
port 2 nsew
rlabel metal3 s 240 44477 240 44477 4 gnd
port 2 nsew
rlabel metal3 s 240 41080 240 41080 4 gnd
port 2 nsew
rlabel metal3 s 240 42897 240 42897 4 gnd
port 2 nsew
rlabel metal3 s 240 41317 240 41317 4 gnd
port 2 nsew
rlabel metal3 s 2808 51911 2808 51911 4 vdd
port 1 nsew
rlabel metal3 s 240 45267 240 45267 4 gnd
port 2 nsew
rlabel metal3 s 2184 51911 2184 51911 4 vdd
port 1 nsew
rlabel metal3 s 936 51911 936 51911 4 vdd
port 1 nsew
rlabel metal3 s 240 44240 240 44240 4 gnd
port 2 nsew
rlabel metal3 s 240 47637 240 47637 4 gnd
port 2 nsew
rlabel metal3 s 240 41870 240 41870 4 gnd
port 2 nsew
rlabel metal3 s 240 51587 240 51587 4 gnd
port 2 nsew
rlabel metal3 s 240 50007 240 50007 4 gnd
port 2 nsew
rlabel metal3 s 240 40843 240 40843 4 gnd
port 2 nsew
rlabel metal3 s 8424 51911 8424 51911 4 vdd
port 1 nsew
rlabel metal3 s 240 48190 240 48190 4 gnd
port 2 nsew
rlabel metal3 s 240 48427 240 48427 4 gnd
port 2 nsew
rlabel metal3 s 6552 51911 6552 51911 4 vdd
port 1 nsew
rlabel metal3 s 5928 51911 5928 51911 4 vdd
port 1 nsew
rlabel metal3 s 240 43687 240 43687 4 gnd
port 2 nsew
rlabel metal3 s 240 42660 240 42660 4 gnd
port 2 nsew
rlabel metal3 s 240 48980 240 48980 4 gnd
port 2 nsew
rlabel metal3 s 240 42107 240 42107 4 gnd
port 2 nsew
rlabel metal3 s 3432 51911 3432 51911 4 vdd
port 1 nsew
rlabel metal3 s 4056 51911 4056 51911 4 vdd
port 1 nsew
rlabel metal3 s 7800 51911 7800 51911 4 vdd
port 1 nsew
rlabel metal3 s 240 45820 240 45820 4 gnd
port 2 nsew
rlabel metal3 s 240 47400 240 47400 4 gnd
port 2 nsew
rlabel metal3 s 240 48743 240 48743 4 gnd
port 2 nsew
rlabel metal3 s 10296 51911 10296 51911 4 vdd
port 1 nsew
rlabel metal3 s 4680 51911 4680 51911 4 vdd
port 1 nsew
rlabel metal3 s 240 41633 240 41633 4 gnd
port 2 nsew
rlabel metal3 s 240 45583 240 45583 4 gnd
port 2 nsew
rlabel metal3 s 9048 51911 9048 51911 4 vdd
port 1 nsew
rlabel metal3 s 240 49770 240 49770 4 gnd
port 2 nsew
rlabel metal3 s 240 43450 240 43450 4 gnd
port 2 nsew
rlabel metal3 s 240 42423 240 42423 4 gnd
port 2 nsew
rlabel metal3 s 240 46610 240 46610 4 gnd
port 2 nsew
rlabel metal3 s 5304 51911 5304 51911 4 vdd
port 1 nsew
rlabel metal3 s 7176 51911 7176 51911 4 vdd
port 1 nsew
rlabel metal3 s 240 39263 240 39263 4 gnd
port 2 nsew
rlabel metal3 s 240 50560 240 50560 4 gnd
port 2 nsew
rlabel metal3 s 1560 51911 1560 51911 4 vdd
port 1 nsew
rlabel metal3 s 9672 51911 9672 51911 4 vdd
port 1 nsew
rlabel metal3 s 240 40053 240 40053 4 gnd
port 2 nsew
rlabel metal3 s 240 40527 240 40527 4 gnd
port 2 nsew
rlabel metal3 s 240 33970 240 33970 4 gnd
port 2 nsew
rlabel metal3 s 240 26860 240 26860 4 gnd
port 2 nsew
rlabel metal3 s 240 34997 240 34997 4 gnd
port 2 nsew
rlabel metal3 s 240 27887 240 27887 4 gnd
port 2 nsew
rlabel metal3 s 240 28440 240 28440 4 gnd
port 2 nsew
rlabel metal3 s 240 38947 240 38947 4 gnd
port 2 nsew
rlabel metal3 s 240 34760 240 34760 4 gnd
port 2 nsew
rlabel metal3 s 240 38473 240 38473 4 gnd
port 2 nsew
rlabel metal3 s 240 28677 240 28677 4 gnd
port 2 nsew
rlabel metal3 s 240 30810 240 30810 4 gnd
port 2 nsew
rlabel metal3 s 240 32390 240 32390 4 gnd
port 2 nsew
rlabel metal3 s 240 33417 240 33417 4 gnd
port 2 nsew
rlabel metal3 s 240 27413 240 27413 4 gnd
port 2 nsew
rlabel metal3 s 240 33180 240 33180 4 gnd
port 2 nsew
rlabel metal3 s 240 30257 240 30257 4 gnd
port 2 nsew
rlabel metal3 s 240 31047 240 31047 4 gnd
port 2 nsew
rlabel metal3 s 240 27650 240 27650 4 gnd
port 2 nsew
rlabel metal3 s 240 37367 240 37367 4 gnd
port 2 nsew
rlabel metal3 s 240 31837 240 31837 4 gnd
port 2 nsew
rlabel metal3 s 240 28993 240 28993 4 gnd
port 2 nsew
rlabel metal3 s 240 33733 240 33733 4 gnd
port 2 nsew
rlabel metal3 s 240 38157 240 38157 4 gnd
port 2 nsew
rlabel metal3 s 240 32943 240 32943 4 gnd
port 2 nsew
rlabel metal3 s 240 32627 240 32627 4 gnd
port 2 nsew
rlabel metal3 s 240 32153 240 32153 4 gnd
port 2 nsew
rlabel metal3 s 240 36893 240 36893 4 gnd
port 2 nsew
rlabel metal3 s 240 35550 240 35550 4 gnd
port 2 nsew
rlabel metal3 s 240 30020 240 30020 4 gnd
port 2 nsew
rlabel metal3 s 240 37920 240 37920 4 gnd
port 2 nsew
rlabel metal3 s 240 34523 240 34523 4 gnd
port 2 nsew
rlabel metal3 s 240 31363 240 31363 4 gnd
port 2 nsew
rlabel metal3 s 240 31600 240 31600 4 gnd
port 2 nsew
rlabel metal3 s 240 28203 240 28203 4 gnd
port 2 nsew
rlabel metal3 s 240 29783 240 29783 4 gnd
port 2 nsew
rlabel metal3 s 240 35787 240 35787 4 gnd
port 2 nsew
rlabel metal3 s 240 29467 240 29467 4 gnd
port 2 nsew
rlabel metal3 s 240 36340 240 36340 4 gnd
port 2 nsew
rlabel metal3 s 240 27097 240 27097 4 gnd
port 2 nsew
rlabel metal3 s 240 38710 240 38710 4 gnd
port 2 nsew
rlabel metal3 s 240 37130 240 37130 4 gnd
port 2 nsew
rlabel metal3 s 240 35313 240 35313 4 gnd
port 2 nsew
rlabel metal3 s 240 30573 240 30573 4 gnd
port 2 nsew
rlabel metal3 s 240 29230 240 29230 4 gnd
port 2 nsew
rlabel metal3 s 240 26307 240 26307 4 gnd
port 2 nsew
rlabel metal3 s 240 36577 240 36577 4 gnd
port 2 nsew
rlabel metal3 s 240 26623 240 26623 4 gnd
port 2 nsew
rlabel metal3 s 240 37683 240 37683 4 gnd
port 2 nsew
rlabel metal3 s 240 36103 240 36103 4 gnd
port 2 nsew
rlabel metal3 s 240 34207 240 34207 4 gnd
port 2 nsew
rlabel metal3 s 240 24253 240 24253 4 gnd
port 2 nsew
rlabel metal3 s 240 24490 240 24490 4 gnd
port 2 nsew
rlabel metal3 s 240 19197 240 19197 4 gnd
port 2 nsew
rlabel metal3 s 240 13193 240 13193 4 gnd
port 2 nsew
rlabel metal3 s 240 23937 240 23937 4 gnd
port 2 nsew
rlabel metal3 s 240 13430 240 13430 4 gnd
port 2 nsew
rlabel metal3 s 240 22120 240 22120 4 gnd
port 2 nsew
rlabel metal3 s 240 16037 240 16037 4 gnd
port 2 nsew
rlabel metal3 s 240 15247 240 15247 4 gnd
port 2 nsew
rlabel metal3 s 240 25833 240 25833 4 gnd
port 2 nsew
rlabel metal3 s 240 16590 240 16590 4 gnd
port 2 nsew
rlabel metal3 s 240 25043 240 25043 4 gnd
port 2 nsew
rlabel metal3 s 240 21330 240 21330 4 gnd
port 2 nsew
rlabel metal3 s 240 16353 240 16353 4 gnd
port 2 nsew
rlabel metal3 s 240 16827 240 16827 4 gnd
port 2 nsew
rlabel metal3 s 240 15010 240 15010 4 gnd
port 2 nsew
rlabel metal3 s 240 23463 240 23463 4 gnd
port 2 nsew
rlabel metal3 s 240 23147 240 23147 4 gnd
port 2 nsew
rlabel metal3 s 240 17933 240 17933 4 gnd
port 2 nsew
rlabel metal3 s 240 21883 240 21883 4 gnd
port 2 nsew
rlabel metal3 s 240 20777 240 20777 4 gnd
port 2 nsew
rlabel metal3 s 240 14457 240 14457 4 gnd
port 2 nsew
rlabel metal3 s 240 20303 240 20303 4 gnd
port 2 nsew
rlabel metal3 s 240 14773 240 14773 4 gnd
port 2 nsew
rlabel metal3 s 240 18407 240 18407 4 gnd
port 2 nsew
rlabel metal3 s 240 15563 240 15563 4 gnd
port 2 nsew
rlabel metal3 s 240 19987 240 19987 4 gnd
port 2 nsew
rlabel metal3 s 240 20540 240 20540 4 gnd
port 2 nsew
rlabel metal3 s 240 23700 240 23700 4 gnd
port 2 nsew
rlabel metal3 s 240 13983 240 13983 4 gnd
port 2 nsew
rlabel metal3 s 240 21093 240 21093 4 gnd
port 2 nsew
rlabel metal3 s 240 17617 240 17617 4 gnd
port 2 nsew
rlabel metal3 s 240 21567 240 21567 4 gnd
port 2 nsew
rlabel metal3 s 240 19513 240 19513 4 gnd
port 2 nsew
rlabel metal3 s 240 18170 240 18170 4 gnd
port 2 nsew
rlabel metal3 s 240 24727 240 24727 4 gnd
port 2 nsew
rlabel metal3 s 240 17380 240 17380 4 gnd
port 2 nsew
rlabel metal3 s 240 25280 240 25280 4 gnd
port 2 nsew
rlabel metal3 s 240 22673 240 22673 4 gnd
port 2 nsew
rlabel metal3 s 240 15800 240 15800 4 gnd
port 2 nsew
rlabel metal3 s 240 17143 240 17143 4 gnd
port 2 nsew
rlabel metal3 s 240 14220 240 14220 4 gnd
port 2 nsew
rlabel metal3 s 240 26070 240 26070 4 gnd
port 2 nsew
rlabel metal3 s 240 19750 240 19750 4 gnd
port 2 nsew
rlabel metal3 s 240 22357 240 22357 4 gnd
port 2 nsew
rlabel metal3 s 240 13667 240 13667 4 gnd
port 2 nsew
rlabel metal3 s 240 22910 240 22910 4 gnd
port 2 nsew
rlabel metal3 s 240 18960 240 18960 4 gnd
port 2 nsew
rlabel metal3 s 240 18723 240 18723 4 gnd
port 2 nsew
rlabel metal3 s 240 25517 240 25517 4 gnd
port 2 nsew
rlabel metal3 s 240 3397 240 3397 4 gnd
port 2 nsew
rlabel metal3 s 240 10270 240 10270 4 gnd
port 2 nsew
rlabel metal3 s 4680 229 4680 229 4 vdd
port 1 nsew
rlabel metal3 s 240 7347 240 7347 4 gnd
port 2 nsew
rlabel metal3 s 240 1343 240 1343 4 gnd
port 2 nsew
rlabel metal3 s 240 6557 240 6557 4 gnd
port 2 nsew
rlabel metal3 s 7176 229 7176 229 4 vdd
port 1 nsew
rlabel metal3 s 7800 229 7800 229 4 vdd
port 1 nsew
rlabel metal3 s 240 9243 240 9243 4 gnd
port 2 nsew
rlabel metal3 s 240 8137 240 8137 4 gnd
port 2 nsew
rlabel metal3 s 240 2370 240 2370 4 gnd
port 2 nsew
rlabel metal3 s 240 4503 240 4503 4 gnd
port 2 nsew
rlabel metal3 s 240 4977 240 4977 4 gnd
port 2 nsew
rlabel metal3 s 9048 229 9048 229 4 vdd
port 1 nsew
rlabel metal3 s 240 790 240 790 4 gnd
port 2 nsew
rlabel metal3 s 240 8690 240 8690 4 gnd
port 2 nsew
rlabel metal3 s 240 4740 240 4740 4 gnd
port 2 nsew
rlabel metal3 s 3432 229 3432 229 4 vdd
port 1 nsew
rlabel metal3 s 2184 229 2184 229 4 vdd
port 1 nsew
rlabel metal3 s 240 1817 240 1817 4 gnd
port 2 nsew
rlabel metal3 s 240 12087 240 12087 4 gnd
port 2 nsew
rlabel metal3 s 240 5530 240 5530 4 gnd
port 2 nsew
rlabel metal3 s 240 5767 240 5767 4 gnd
port 2 nsew
rlabel metal3 s 240 10823 240 10823 4 gnd
port 2 nsew
rlabel metal3 s 240 553 240 553 4 gnd
port 2 nsew
rlabel metal3 s 240 8927 240 8927 4 gnd
port 2 nsew
rlabel metal3 s 6552 229 6552 229 4 vdd
port 1 nsew
rlabel metal3 s 240 7110 240 7110 4 gnd
port 2 nsew
rlabel metal3 s 240 2923 240 2923 4 gnd
port 2 nsew
rlabel metal3 s 240 1027 240 1027 4 gnd
port 2 nsew
rlabel metal3 s 240 8453 240 8453 4 gnd
port 2 nsew
rlabel metal3 s 240 6083 240 6083 4 gnd
port 2 nsew
rlabel metal3 s 240 2133 240 2133 4 gnd
port 2 nsew
rlabel metal3 s 240 3713 240 3713 4 gnd
port 2 nsew
rlabel metal3 s 2808 229 2808 229 4 vdd
port 1 nsew
rlabel metal3 s 9672 229 9672 229 4 vdd
port 1 nsew
rlabel metal3 s 240 3160 240 3160 4 gnd
port 2 nsew
rlabel metal3 s 240 2607 240 2607 4 gnd
port 2 nsew
rlabel metal3 s 240 7900 240 7900 4 gnd
port 2 nsew
rlabel metal3 s 240 5293 240 5293 4 gnd
port 2 nsew
rlabel metal3 s 240 12640 240 12640 4 gnd
port 2 nsew
rlabel metal3 s 240 11850 240 11850 4 gnd
port 2 nsew
rlabel metal3 s 240 12403 240 12403 4 gnd
port 2 nsew
rlabel metal3 s 240 10033 240 10033 4 gnd
port 2 nsew
rlabel metal3 s 1560 229 1560 229 4 vdd
port 1 nsew
rlabel metal3 s 240 11297 240 11297 4 gnd
port 2 nsew
rlabel metal3 s 240 11613 240 11613 4 gnd
port 2 nsew
rlabel metal3 s 240 6873 240 6873 4 gnd
port 2 nsew
rlabel metal3 s 240 9717 240 9717 4 gnd
port 2 nsew
rlabel metal3 s 240 10507 240 10507 4 gnd
port 2 nsew
rlabel metal3 s 240 6320 240 6320 4 gnd
port 2 nsew
rlabel metal3 s 240 12877 240 12877 4 gnd
port 2 nsew
rlabel metal3 s 936 229 936 229 4 vdd
port 1 nsew
rlabel metal3 s 10296 229 10296 229 4 vdd
port 1 nsew
rlabel metal3 s 5928 229 5928 229 4 vdd
port 1 nsew
rlabel metal3 s 240 9480 240 9480 4 gnd
port 2 nsew
rlabel metal3 s 4056 229 4056 229 4 vdd
port 1 nsew
rlabel metal3 s 240 7663 240 7663 4 gnd
port 2 nsew
rlabel metal3 s 240 3950 240 3950 4 gnd
port 2 nsew
rlabel metal3 s 240 1580 240 1580 4 gnd
port 2 nsew
rlabel metal3 s 240 11060 240 11060 4 gnd
port 2 nsew
rlabel metal3 s 5304 229 5304 229 4 vdd
port 1 nsew
rlabel metal3 s 240 4187 240 4187 4 gnd
port 2 nsew
rlabel metal3 s 8424 229 8424 229 4 vdd
port 1 nsew
rlabel metal3 s 20280 229 20280 229 4 vdd
port 1 nsew
rlabel metal3 s 15912 229 15912 229 4 vdd
port 1 nsew
rlabel metal3 s 16536 229 16536 229 4 vdd
port 1 nsew
rlabel metal3 s 11544 229 11544 229 4 vdd
port 1 nsew
rlabel metal3 s 18408 229 18408 229 4 vdd
port 1 nsew
rlabel metal3 s 20904 229 20904 229 4 vdd
port 1 nsew
rlabel metal3 s 19032 229 19032 229 4 vdd
port 1 nsew
rlabel metal3 s 13416 229 13416 229 4 vdd
port 1 nsew
rlabel metal3 s 19656 229 19656 229 4 vdd
port 1 nsew
rlabel metal3 s 14664 229 14664 229 4 vdd
port 1 nsew
rlabel metal3 s 12168 229 12168 229 4 vdd
port 1 nsew
rlabel metal3 s 17160 229 17160 229 4 vdd
port 1 nsew
rlabel metal3 s 15288 229 15288 229 4 vdd
port 1 nsew
rlabel metal3 s 12792 229 12792 229 4 vdd
port 1 nsew
rlabel metal3 s 17784 229 17784 229 4 vdd
port 1 nsew
rlabel metal3 s 10920 229 10920 229 4 vdd
port 1 nsew
rlabel metal3 s 14040 229 14040 229 4 vdd
port 1 nsew
rlabel metal3 s 42192 15800 42192 15800 4 gnd
port 2 nsew
rlabel metal3 s 42192 20540 42192 20540 4 gnd
port 2 nsew
rlabel metal3 s 42192 17143 42192 17143 4 gnd
port 2 nsew
rlabel metal3 s 42192 26070 42192 26070 4 gnd
port 2 nsew
rlabel metal3 s 42192 19513 42192 19513 4 gnd
port 2 nsew
rlabel metal3 s 42192 21567 42192 21567 4 gnd
port 2 nsew
rlabel metal3 s 42192 25043 42192 25043 4 gnd
port 2 nsew
rlabel metal3 s 42192 21330 42192 21330 4 gnd
port 2 nsew
rlabel metal3 s 42192 24490 42192 24490 4 gnd
port 2 nsew
rlabel metal3 s 42192 21883 42192 21883 4 gnd
port 2 nsew
rlabel metal3 s 42192 14220 42192 14220 4 gnd
port 2 nsew
rlabel metal3 s 42192 22673 42192 22673 4 gnd
port 2 nsew
rlabel metal3 s 42192 20777 42192 20777 4 gnd
port 2 nsew
rlabel metal3 s 42192 23700 42192 23700 4 gnd
port 2 nsew
rlabel metal3 s 42192 16827 42192 16827 4 gnd
port 2 nsew
rlabel metal3 s 42192 13430 42192 13430 4 gnd
port 2 nsew
rlabel metal3 s 42192 16353 42192 16353 4 gnd
port 2 nsew
rlabel metal3 s 42192 16590 42192 16590 4 gnd
port 2 nsew
rlabel metal3 s 42192 20303 42192 20303 4 gnd
port 2 nsew
rlabel metal3 s 42192 17933 42192 17933 4 gnd
port 2 nsew
rlabel metal3 s 42192 13983 42192 13983 4 gnd
port 2 nsew
rlabel metal3 s 42192 19750 42192 19750 4 gnd
port 2 nsew
rlabel metal3 s 42192 25280 42192 25280 4 gnd
port 2 nsew
rlabel metal3 s 42192 15010 42192 15010 4 gnd
port 2 nsew
rlabel metal3 s 42192 18407 42192 18407 4 gnd
port 2 nsew
rlabel metal3 s 42192 19197 42192 19197 4 gnd
port 2 nsew
rlabel metal3 s 42192 25517 42192 25517 4 gnd
port 2 nsew
rlabel metal3 s 42192 17617 42192 17617 4 gnd
port 2 nsew
rlabel metal3 s 42192 24727 42192 24727 4 gnd
port 2 nsew
rlabel metal3 s 42192 22357 42192 22357 4 gnd
port 2 nsew
rlabel metal3 s 42192 15247 42192 15247 4 gnd
port 2 nsew
rlabel metal3 s 42192 14773 42192 14773 4 gnd
port 2 nsew
rlabel metal3 s 42192 18170 42192 18170 4 gnd
port 2 nsew
rlabel metal3 s 42192 16037 42192 16037 4 gnd
port 2 nsew
rlabel metal3 s 42192 13193 42192 13193 4 gnd
port 2 nsew
rlabel metal3 s 42192 15563 42192 15563 4 gnd
port 2 nsew
rlabel metal3 s 42192 19987 42192 19987 4 gnd
port 2 nsew
rlabel metal3 s 42192 17380 42192 17380 4 gnd
port 2 nsew
rlabel metal3 s 42192 18723 42192 18723 4 gnd
port 2 nsew
rlabel metal3 s 42192 23463 42192 23463 4 gnd
port 2 nsew
rlabel metal3 s 42192 23937 42192 23937 4 gnd
port 2 nsew
rlabel metal3 s 42192 21093 42192 21093 4 gnd
port 2 nsew
rlabel metal3 s 42192 25833 42192 25833 4 gnd
port 2 nsew
rlabel metal3 s 42192 22910 42192 22910 4 gnd
port 2 nsew
rlabel metal3 s 42192 14457 42192 14457 4 gnd
port 2 nsew
rlabel metal3 s 42192 18960 42192 18960 4 gnd
port 2 nsew
rlabel metal3 s 42192 24253 42192 24253 4 gnd
port 2 nsew
rlabel metal3 s 42192 23147 42192 23147 4 gnd
port 2 nsew
rlabel metal3 s 42192 13667 42192 13667 4 gnd
port 2 nsew
rlabel metal3 s 42192 22120 42192 22120 4 gnd
port 2 nsew
rlabel metal3 s 27144 229 27144 229 4 vdd
port 1 nsew
rlabel metal3 s 30888 229 30888 229 4 vdd
port 1 nsew
rlabel metal3 s 24648 229 24648 229 4 vdd
port 1 nsew
rlabel metal3 s 22776 229 22776 229 4 vdd
port 1 nsew
rlabel metal3 s 21528 229 21528 229 4 vdd
port 1 nsew
rlabel metal3 s 28392 229 28392 229 4 vdd
port 1 nsew
rlabel metal3 s 23400 229 23400 229 4 vdd
port 1 nsew
rlabel metal3 s 26520 229 26520 229 4 vdd
port 1 nsew
rlabel metal3 s 25896 229 25896 229 4 vdd
port 1 nsew
rlabel metal3 s 25272 229 25272 229 4 vdd
port 1 nsew
rlabel metal3 s 27768 229 27768 229 4 vdd
port 1 nsew
rlabel metal3 s 30264 229 30264 229 4 vdd
port 1 nsew
rlabel metal3 s 29640 229 29640 229 4 vdd
port 1 nsew
rlabel metal3 s 31512 229 31512 229 4 vdd
port 1 nsew
rlabel metal3 s 29016 229 29016 229 4 vdd
port 1 nsew
rlabel metal3 s 22152 229 22152 229 4 vdd
port 1 nsew
rlabel metal3 s 24024 229 24024 229 4 vdd
port 1 nsew
rlabel metal3 s 42192 3397 42192 3397 4 gnd
port 2 nsew
rlabel metal3 s 32136 229 32136 229 4 vdd
port 1 nsew
rlabel metal3 s 34632 229 34632 229 4 vdd
port 1 nsew
rlabel metal3 s 42192 2923 42192 2923 4 gnd
port 2 nsew
rlabel metal3 s 37752 229 37752 229 4 vdd
port 1 nsew
rlabel metal3 s 42192 10270 42192 10270 4 gnd
port 2 nsew
rlabel metal3 s 42192 3950 42192 3950 4 gnd
port 2 nsew
rlabel metal3 s 42192 4503 42192 4503 4 gnd
port 2 nsew
rlabel metal3 s 42192 6873 42192 6873 4 gnd
port 2 nsew
rlabel metal3 s 42192 8690 42192 8690 4 gnd
port 2 nsew
rlabel metal3 s 42192 9717 42192 9717 4 gnd
port 2 nsew
rlabel metal3 s 42192 4187 42192 4187 4 gnd
port 2 nsew
rlabel metal3 s 35880 229 35880 229 4 vdd
port 1 nsew
rlabel metal3 s 42192 7900 42192 7900 4 gnd
port 2 nsew
rlabel metal3 s 38376 229 38376 229 4 vdd
port 1 nsew
rlabel metal3 s 41496 229 41496 229 4 vdd
port 1 nsew
rlabel metal3 s 42192 6083 42192 6083 4 gnd
port 2 nsew
rlabel metal3 s 42192 12087 42192 12087 4 gnd
port 2 nsew
rlabel metal3 s 42192 8137 42192 8137 4 gnd
port 2 nsew
rlabel metal3 s 35256 229 35256 229 4 vdd
port 1 nsew
rlabel metal3 s 42192 2370 42192 2370 4 gnd
port 2 nsew
rlabel metal3 s 42192 6320 42192 6320 4 gnd
port 2 nsew
rlabel metal3 s 37128 229 37128 229 4 vdd
port 1 nsew
rlabel metal3 s 42192 10033 42192 10033 4 gnd
port 2 nsew
rlabel metal3 s 42192 11613 42192 11613 4 gnd
port 2 nsew
rlabel metal3 s 42192 12877 42192 12877 4 gnd
port 2 nsew
rlabel metal3 s 42192 12403 42192 12403 4 gnd
port 2 nsew
rlabel metal3 s 42192 1580 42192 1580 4 gnd
port 2 nsew
rlabel metal3 s 42192 2607 42192 2607 4 gnd
port 2 nsew
rlabel metal3 s 42192 553 42192 553 4 gnd
port 2 nsew
rlabel metal3 s 42192 5767 42192 5767 4 gnd
port 2 nsew
rlabel metal3 s 39000 229 39000 229 4 vdd
port 1 nsew
rlabel metal3 s 42192 3713 42192 3713 4 gnd
port 2 nsew
rlabel metal3 s 36504 229 36504 229 4 vdd
port 1 nsew
rlabel metal3 s 42192 5530 42192 5530 4 gnd
port 2 nsew
rlabel metal3 s 42192 7110 42192 7110 4 gnd
port 2 nsew
rlabel metal3 s 39624 229 39624 229 4 vdd
port 1 nsew
rlabel metal3 s 42192 4977 42192 4977 4 gnd
port 2 nsew
rlabel metal3 s 42192 2133 42192 2133 4 gnd
port 2 nsew
rlabel metal3 s 42192 1027 42192 1027 4 gnd
port 2 nsew
rlabel metal3 s 42192 12640 42192 12640 4 gnd
port 2 nsew
rlabel metal3 s 42192 11850 42192 11850 4 gnd
port 2 nsew
rlabel metal3 s 42192 10507 42192 10507 4 gnd
port 2 nsew
rlabel metal3 s 42192 1343 42192 1343 4 gnd
port 2 nsew
rlabel metal3 s 33384 229 33384 229 4 vdd
port 1 nsew
rlabel metal3 s 42192 11060 42192 11060 4 gnd
port 2 nsew
rlabel metal3 s 42192 9243 42192 9243 4 gnd
port 2 nsew
rlabel metal3 s 40248 229 40248 229 4 vdd
port 1 nsew
rlabel metal3 s 42192 3160 42192 3160 4 gnd
port 2 nsew
rlabel metal3 s 42192 5293 42192 5293 4 gnd
port 2 nsew
rlabel metal3 s 42192 7663 42192 7663 4 gnd
port 2 nsew
rlabel metal3 s 40872 229 40872 229 4 vdd
port 1 nsew
rlabel metal3 s 32760 229 32760 229 4 vdd
port 1 nsew
rlabel metal3 s 42192 10823 42192 10823 4 gnd
port 2 nsew
rlabel metal3 s 42192 4740 42192 4740 4 gnd
port 2 nsew
rlabel metal3 s 34008 229 34008 229 4 vdd
port 1 nsew
rlabel metal3 s 42192 11297 42192 11297 4 gnd
port 2 nsew
rlabel metal3 s 42192 6557 42192 6557 4 gnd
port 2 nsew
rlabel metal3 s 42192 790 42192 790 4 gnd
port 2 nsew
rlabel metal3 s 42192 9480 42192 9480 4 gnd
port 2 nsew
rlabel metal3 s 42192 8453 42192 8453 4 gnd
port 2 nsew
rlabel metal3 s 42192 7347 42192 7347 4 gnd
port 2 nsew
rlabel metal3 s 42192 8927 42192 8927 4 gnd
port 2 nsew
rlabel metal3 s 42192 1817 42192 1817 4 gnd
port 2 nsew
<< properties >>
string FIXED_BBOX 0 0 42432 52140
string GDS_END 5096578
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sram_1rw1r_32_256_8_sky130.gds
string GDS_START 4888228
<< end >>
