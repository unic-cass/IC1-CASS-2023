magic
tech sky130B
magscale 1 2
timestamp 1676037725
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_0
timestamp 1676037725
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd__example_5595914180851  sky130_fd_pr__hvdfl1sd__example_5595914180851_0
timestamp 1676037725
transform 1 0 100 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 31960798
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 31959870
<< end >>
