magic
tech sky130B
magscale 1 2
timestamp 1676037725
<< nwell >>
rect -38 261 774 582
<< pwell >>
rect 1 21 735 203
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 177
rect 165 47 195 177
rect 318 47 348 177
rect 430 47 460 177
rect 531 47 561 177
rect 627 47 657 177
<< scpmoshvt >>
rect 79 297 109 497
rect 163 297 193 497
rect 351 297 381 497
rect 459 297 489 497
rect 555 297 585 497
rect 627 297 657 497
<< ndiff >>
rect 27 165 79 177
rect 27 131 35 165
rect 69 131 79 165
rect 27 93 79 131
rect 27 59 35 93
rect 69 59 79 93
rect 27 47 79 59
rect 109 169 165 177
rect 109 135 120 169
rect 154 135 165 169
rect 109 101 165 135
rect 109 67 119 101
rect 153 67 165 101
rect 109 47 165 67
rect 195 89 318 177
rect 195 55 205 89
rect 239 55 274 89
rect 308 55 318 89
rect 195 47 318 55
rect 348 47 430 177
rect 460 157 531 177
rect 460 123 471 157
rect 505 123 531 157
rect 460 89 531 123
rect 460 55 471 89
rect 505 55 531 89
rect 460 47 531 55
rect 561 89 627 177
rect 561 55 577 89
rect 611 55 627 89
rect 561 47 627 55
rect 657 165 709 177
rect 657 131 667 165
rect 701 131 709 165
rect 657 97 709 131
rect 657 63 667 97
rect 701 63 709 97
rect 657 47 709 63
<< pdiff >>
rect 27 484 79 497
rect 27 450 35 484
rect 69 450 79 484
rect 27 416 79 450
rect 27 382 35 416
rect 69 382 79 416
rect 27 348 79 382
rect 27 314 35 348
rect 69 314 79 348
rect 27 297 79 314
rect 109 430 163 497
rect 109 396 119 430
rect 153 396 163 430
rect 109 342 163 396
rect 109 308 119 342
rect 153 308 163 342
rect 109 297 163 308
rect 193 485 245 497
rect 193 451 203 485
rect 237 451 245 485
rect 193 417 245 451
rect 193 383 203 417
rect 237 383 245 417
rect 193 297 245 383
rect 299 485 351 497
rect 299 451 307 485
rect 341 451 351 485
rect 299 417 351 451
rect 299 383 307 417
rect 341 383 351 417
rect 299 297 351 383
rect 381 488 459 497
rect 381 454 404 488
rect 438 454 459 488
rect 381 297 459 454
rect 489 485 555 497
rect 489 451 509 485
rect 543 451 555 485
rect 489 417 555 451
rect 489 383 509 417
rect 543 383 555 417
rect 489 297 555 383
rect 585 297 627 497
rect 657 436 709 497
rect 657 402 667 436
rect 701 402 709 436
rect 657 368 709 402
rect 657 334 667 368
rect 701 334 709 368
rect 657 297 709 334
<< ndiffc >>
rect 35 131 69 165
rect 35 59 69 93
rect 120 135 154 169
rect 119 67 153 101
rect 205 55 239 89
rect 274 55 308 89
rect 471 123 505 157
rect 471 55 505 89
rect 577 55 611 89
rect 667 131 701 165
rect 667 63 701 97
<< pdiffc >>
rect 35 450 69 484
rect 35 382 69 416
rect 35 314 69 348
rect 119 396 153 430
rect 119 308 153 342
rect 203 451 237 485
rect 203 383 237 417
rect 307 451 341 485
rect 307 383 341 417
rect 404 454 438 488
rect 509 451 543 485
rect 509 383 543 417
rect 667 402 701 436
rect 667 334 701 368
<< poly >>
rect 79 497 109 523
rect 163 497 193 523
rect 351 497 381 523
rect 459 497 489 523
rect 555 497 585 523
rect 627 497 657 523
rect 79 265 109 297
rect 163 265 193 297
rect 351 265 381 297
rect 459 265 489 297
rect 555 265 585 297
rect 79 249 244 265
rect 79 215 200 249
rect 234 215 244 249
rect 79 200 244 215
rect 79 177 109 200
rect 165 199 244 200
rect 302 249 381 265
rect 302 215 312 249
rect 346 215 381 249
rect 302 199 381 215
rect 165 177 195 199
rect 318 198 381 199
rect 430 249 489 265
rect 430 215 440 249
rect 474 215 489 249
rect 430 199 489 215
rect 531 249 585 265
rect 531 215 541 249
rect 575 215 585 249
rect 531 199 585 215
rect 627 265 657 297
rect 627 249 715 265
rect 627 215 669 249
rect 703 215 715 249
rect 627 199 715 215
rect 318 177 348 198
rect 430 177 460 199
rect 531 177 561 199
rect 627 177 657 199
rect 79 21 109 47
rect 165 21 195 47
rect 318 21 348 47
rect 430 21 460 47
rect 531 21 561 47
rect 627 21 657 47
<< polycont >>
rect 200 215 234 249
rect 312 215 346 249
rect 440 215 474 249
rect 541 215 575 249
rect 669 215 703 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 18 484 77 527
rect 18 450 35 484
rect 69 450 77 484
rect 200 485 251 527
rect 18 416 77 450
rect 18 382 35 416
rect 69 382 77 416
rect 18 348 77 382
rect 18 314 35 348
rect 69 314 77 348
rect 18 298 77 314
rect 111 430 157 467
rect 111 396 119 430
rect 153 396 157 430
rect 111 342 157 396
rect 200 451 203 485
rect 237 451 251 485
rect 200 417 251 451
rect 200 383 203 417
rect 237 383 251 417
rect 200 366 251 383
rect 291 485 357 493
rect 291 451 307 485
rect 341 451 357 485
rect 291 417 357 451
rect 391 488 446 527
rect 391 454 404 488
rect 438 454 446 488
rect 391 438 446 454
rect 493 485 559 493
rect 493 451 509 485
rect 543 451 559 485
rect 291 383 307 417
rect 341 404 357 417
rect 493 417 559 451
rect 493 404 509 417
rect 341 383 509 404
rect 543 383 559 417
rect 291 368 559 383
rect 651 436 717 465
rect 651 402 667 436
rect 701 402 717 436
rect 651 368 717 402
rect 111 308 119 342
rect 153 308 157 342
rect 651 334 667 368
rect 701 334 717 368
rect 651 332 717 334
rect 18 165 77 181
rect 18 131 35 165
rect 69 131 77 165
rect 18 93 77 131
rect 18 59 35 93
rect 69 59 77 93
rect 18 17 77 59
rect 111 169 157 308
rect 111 135 120 169
rect 154 135 157 169
rect 200 298 717 332
rect 200 249 262 298
rect 234 215 262 249
rect 200 175 262 215
rect 296 249 362 255
rect 296 215 312 249
rect 346 215 362 249
rect 296 209 362 215
rect 396 249 490 255
rect 396 215 440 249
rect 474 215 490 249
rect 396 209 490 215
rect 524 249 614 255
rect 524 215 541 249
rect 575 215 614 249
rect 524 209 614 215
rect 652 249 719 255
rect 652 215 669 249
rect 703 215 719 249
rect 652 209 719 215
rect 200 165 717 175
rect 200 157 667 165
rect 200 139 471 157
rect 111 127 157 135
rect 111 101 155 127
rect 111 67 119 101
rect 153 67 155 101
rect 455 123 471 139
rect 505 139 667 157
rect 505 123 521 139
rect 455 89 521 123
rect 651 131 667 139
rect 701 131 717 165
rect 111 51 155 67
rect 189 55 205 89
rect 239 55 274 89
rect 308 55 359 89
rect 455 55 471 89
rect 505 55 521 89
rect 562 89 617 105
rect 562 55 577 89
rect 611 55 617 89
rect 651 97 717 131
rect 651 63 667 97
rect 701 63 717 97
rect 651 55 717 63
rect 189 17 359 55
rect 562 17 617 55
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
flabel locali s 122 425 156 459 0 FreeSans 400 0 0 0 X
port 9 nsew signal output
flabel locali s 304 221 338 255 0 FreeSans 400 0 0 0 A2
port 2 nsew signal input
flabel locali s 396 221 430 255 0 FreeSans 400 0 0 0 A1
port 1 nsew signal input
flabel locali s 580 221 614 255 0 FreeSans 400 0 0 0 B1
port 3 nsew signal input
flabel locali s 672 221 706 255 0 FreeSans 400 0 0 0 C1
port 4 nsew signal input
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 a211o_2
rlabel metal1 s 0 -48 736 48 1 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 496 736 592 1 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 736 544
string GDS_END 3635572
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3629008
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 18.400 0.000 
<< end >>
