magic
tech sky130A
magscale 1 2
timestamp 1676037725
<< nwell >>
rect -66 377 3138 897
<< pwell >>
rect 454 217 1974 283
rect 2623 217 3068 317
rect 4 43 3068 217
rect -26 -43 3098 43
<< mvnmos >>
rect 87 107 187 191
rect 243 107 343 191
rect 537 173 637 257
rect 679 173 779 257
rect 835 173 935 257
rect 991 173 1091 257
rect 1133 173 1233 257
rect 1280 173 1380 257
rect 1633 107 1733 257
rect 1789 107 1889 257
rect 2706 207 2806 291
rect 1989 107 2089 191
rect 2131 107 2231 191
rect 2287 107 2387 191
rect 2429 107 2529 191
rect 2885 141 2985 291
<< mvpmos >>
rect 83 537 183 687
rect 239 537 339 687
rect 509 632 609 716
rect 665 632 765 716
rect 821 632 921 716
rect 977 632 1077 716
rect 1119 632 1219 716
rect 1291 632 1391 716
rect 1619 543 1719 743
rect 1775 543 1875 743
rect 1954 543 2054 627
rect 2096 543 2196 627
rect 2273 543 2373 627
rect 2429 543 2529 627
rect 2714 443 2814 593
rect 2889 443 2989 743
<< mvndiff >>
rect 480 232 537 257
rect 480 198 492 232
rect 526 198 537 232
rect 30 166 87 191
rect 30 132 42 166
rect 76 132 87 166
rect 30 107 87 132
rect 187 166 243 191
rect 187 132 198 166
rect 232 132 243 166
rect 187 107 243 132
rect 343 166 400 191
rect 480 173 537 198
rect 637 173 679 257
rect 779 232 835 257
rect 779 198 790 232
rect 824 198 835 232
rect 779 173 835 198
rect 935 232 991 257
rect 935 198 946 232
rect 980 198 991 232
rect 935 173 991 198
rect 1091 173 1133 257
rect 1233 173 1280 257
rect 1380 173 1633 257
rect 343 132 354 166
rect 388 132 400 166
rect 1560 169 1633 173
rect 343 107 400 132
rect 1560 135 1572 169
rect 1606 135 1633 169
rect 1560 107 1633 135
rect 1733 249 1789 257
rect 1733 215 1744 249
rect 1778 215 1789 249
rect 1733 157 1789 215
rect 1733 123 1744 157
rect 1778 123 1789 157
rect 1733 107 1789 123
rect 1889 249 1948 257
rect 1889 215 1902 249
rect 1936 215 1948 249
rect 1889 191 1948 215
rect 2649 266 2706 291
rect 2649 232 2661 266
rect 2695 232 2706 266
rect 2649 207 2706 232
rect 2806 283 2885 291
rect 2806 249 2840 283
rect 2874 249 2885 283
rect 2806 207 2885 249
rect 1889 157 1989 191
rect 1889 123 1902 157
rect 1936 123 1989 157
rect 1889 107 1989 123
rect 2089 107 2131 191
rect 2231 166 2287 191
rect 2231 132 2242 166
rect 2276 132 2287 166
rect 2231 107 2287 132
rect 2387 107 2429 191
rect 2529 166 2586 191
rect 2828 183 2885 207
rect 2529 132 2540 166
rect 2574 132 2586 166
rect 2828 149 2840 183
rect 2874 149 2885 183
rect 2828 141 2885 149
rect 2985 283 3042 291
rect 2985 249 2996 283
rect 3030 249 3042 283
rect 2985 183 3042 249
rect 2985 149 2996 183
rect 3030 149 3042 183
rect 2985 141 3042 149
rect 2529 107 2586 132
<< mvpdiff >>
rect 1562 730 1619 743
rect 30 675 83 687
rect 30 641 38 675
rect 72 641 83 675
rect 30 583 83 641
rect 30 549 38 583
rect 72 549 83 583
rect 30 537 83 549
rect 183 679 239 687
rect 183 645 194 679
rect 228 645 239 679
rect 183 579 239 645
rect 183 545 194 579
rect 228 545 239 579
rect 183 537 239 545
rect 339 675 392 687
rect 339 641 350 675
rect 384 641 392 675
rect 339 583 392 641
rect 452 674 509 716
rect 452 640 464 674
rect 498 640 509 674
rect 452 632 509 640
rect 609 708 665 716
rect 609 674 620 708
rect 654 674 665 708
rect 609 632 665 674
rect 765 674 821 716
rect 765 640 776 674
rect 810 640 821 674
rect 765 632 821 640
rect 921 682 977 716
rect 921 648 932 682
rect 966 648 977 682
rect 921 632 977 648
rect 1077 632 1119 716
rect 1219 693 1291 716
rect 1219 659 1230 693
rect 1264 659 1291 693
rect 1219 632 1291 659
rect 1391 682 1448 716
rect 1391 648 1402 682
rect 1436 648 1448 682
rect 1391 632 1448 648
rect 1562 696 1574 730
rect 1608 696 1619 730
rect 339 549 350 583
rect 384 549 392 583
rect 339 537 392 549
rect 1562 543 1619 696
rect 1719 585 1775 743
rect 1719 551 1730 585
rect 1764 551 1775 585
rect 1719 543 1775 551
rect 1875 735 1932 743
rect 1875 701 1886 735
rect 1920 701 1932 735
rect 1875 660 1932 701
rect 1875 626 1886 660
rect 1920 627 1932 660
rect 2836 731 2889 743
rect 2836 697 2844 731
rect 2878 697 2889 731
rect 2836 651 2889 697
rect 1920 626 1954 627
rect 1875 585 1954 626
rect 1875 551 1886 585
rect 1920 551 1954 585
rect 1875 543 1954 551
rect 2054 543 2096 627
rect 2196 602 2273 627
rect 2196 568 2207 602
rect 2241 568 2273 602
rect 2196 543 2273 568
rect 2373 602 2429 627
rect 2373 568 2384 602
rect 2418 568 2429 602
rect 2373 543 2429 568
rect 2529 615 2586 627
rect 2529 581 2540 615
rect 2574 581 2586 615
rect 2836 617 2844 651
rect 2878 617 2889 651
rect 2836 593 2889 617
rect 2529 543 2586 581
rect 2657 585 2714 593
rect 2657 551 2669 585
rect 2703 551 2714 585
rect 2657 485 2714 551
rect 2657 451 2669 485
rect 2703 451 2714 485
rect 2657 443 2714 451
rect 2814 569 2889 593
rect 2814 535 2844 569
rect 2878 535 2889 569
rect 2814 489 2889 535
rect 2814 455 2844 489
rect 2878 455 2889 489
rect 2814 443 2889 455
rect 2989 731 3042 743
rect 2989 697 3000 731
rect 3034 697 3042 731
rect 2989 651 3042 697
rect 2989 617 3000 651
rect 3034 617 3042 651
rect 2989 569 3042 617
rect 2989 535 3000 569
rect 3034 535 3042 569
rect 2989 489 3042 535
rect 2989 455 3000 489
rect 3034 455 3042 489
rect 2989 443 3042 455
<< mvndiffc >>
rect 492 198 526 232
rect 42 132 76 166
rect 198 132 232 166
rect 790 198 824 232
rect 946 198 980 232
rect 354 132 388 166
rect 1572 135 1606 169
rect 1744 215 1778 249
rect 1744 123 1778 157
rect 1902 215 1936 249
rect 2661 232 2695 266
rect 2840 249 2874 283
rect 1902 123 1936 157
rect 2242 132 2276 166
rect 2540 132 2574 166
rect 2840 149 2874 183
rect 2996 249 3030 283
rect 2996 149 3030 183
<< mvpdiffc >>
rect 38 641 72 675
rect 38 549 72 583
rect 194 645 228 679
rect 194 545 228 579
rect 350 641 384 675
rect 464 640 498 674
rect 620 674 654 708
rect 776 640 810 674
rect 932 648 966 682
rect 1230 659 1264 693
rect 1402 648 1436 682
rect 1574 696 1608 730
rect 350 549 384 583
rect 1730 551 1764 585
rect 1886 701 1920 735
rect 1886 626 1920 660
rect 2844 697 2878 731
rect 1886 551 1920 585
rect 2207 568 2241 602
rect 2384 568 2418 602
rect 2540 581 2574 615
rect 2844 617 2878 651
rect 2669 551 2703 585
rect 2669 451 2703 485
rect 2844 535 2878 569
rect 2844 455 2878 489
rect 3000 697 3034 731
rect 3000 617 3034 651
rect 3000 535 3034 569
rect 3000 455 3034 489
<< mvpsubdiff >>
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3072 17
<< mvnsubdiff >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2239 831
rect 2273 797 2335 831
rect 2369 797 2431 831
rect 2465 797 2527 831
rect 2561 797 2623 831
rect 2657 797 2719 831
rect 2753 797 2815 831
rect 2849 797 2911 831
rect 2945 797 3007 831
rect 3041 797 3072 831
<< mvpsubdiffcont >>
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
rect 3007 -17 3041 17
<< mvnsubdiffcont >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 895 797 929 831
rect 991 797 1025 831
rect 1087 797 1121 831
rect 1183 797 1217 831
rect 1279 797 1313 831
rect 1375 797 1409 831
rect 1471 797 1505 831
rect 1567 797 1601 831
rect 1663 797 1697 831
rect 1759 797 1793 831
rect 1855 797 1889 831
rect 1951 797 1985 831
rect 2047 797 2081 831
rect 2143 797 2177 831
rect 2239 797 2273 831
rect 2335 797 2369 831
rect 2431 797 2465 831
rect 2527 797 2561 831
rect 2623 797 2657 831
rect 2719 797 2753 831
rect 2815 797 2849 831
rect 2911 797 2945 831
rect 3007 797 3041 831
<< poly >>
rect 1619 743 1719 769
rect 1775 743 1875 769
rect 2889 743 2989 769
rect 509 716 609 742
rect 665 716 765 742
rect 821 716 921 742
rect 977 716 1077 742
rect 1119 716 1219 742
rect 1291 716 1391 742
rect 83 687 183 713
rect 239 687 339 713
rect 83 373 183 537
rect 239 511 339 537
rect 239 489 343 511
rect 239 455 264 489
rect 298 455 343 489
rect 239 421 343 455
rect 239 387 264 421
rect 298 387 343 421
rect 83 353 187 373
rect 239 367 343 387
rect 83 319 128 353
rect 162 319 187 353
rect 83 285 187 319
rect 83 251 128 285
rect 162 251 187 285
rect 83 217 187 251
rect 87 191 187 217
rect 243 191 343 367
rect 509 462 609 632
rect 665 610 765 632
rect 665 510 779 610
rect 821 584 921 632
rect 821 550 851 584
rect 885 550 921 584
rect 821 534 921 550
rect 977 584 1077 632
rect 977 550 1012 584
rect 1046 550 1077 584
rect 977 534 1077 550
rect 509 442 637 462
rect 509 408 555 442
rect 589 408 637 442
rect 509 374 637 408
rect 509 340 555 374
rect 589 340 637 374
rect 509 279 637 340
rect 537 257 637 279
rect 679 405 779 510
rect 963 492 1077 534
rect 1119 606 1219 632
rect 1291 606 1391 632
rect 1119 506 1238 606
rect 679 371 699 405
rect 733 371 779 405
rect 679 337 779 371
rect 679 303 699 337
rect 733 303 779 337
rect 679 257 779 303
rect 835 457 1077 492
rect 1133 468 1238 506
rect 835 415 949 457
rect 1133 434 1184 468
rect 1218 434 1238 468
rect 835 257 935 415
rect 991 399 1091 415
rect 991 365 1011 399
rect 1045 365 1091 399
rect 991 331 1091 365
rect 991 297 1011 331
rect 1045 297 1091 331
rect 991 257 1091 297
rect 1133 400 1238 434
rect 1133 366 1184 400
rect 1218 366 1238 400
rect 1133 279 1238 366
rect 1280 399 1391 606
rect 1954 627 2054 653
rect 2096 627 2196 653
rect 2273 627 2373 653
rect 2429 627 2529 653
rect 2714 593 2814 619
rect 1280 365 1337 399
rect 1371 365 1391 399
rect 1619 379 1719 543
rect 1775 517 1875 543
rect 1775 495 1866 517
rect 1775 461 1816 495
rect 1850 461 1866 495
rect 1954 487 2054 543
rect 1775 427 1866 461
rect 1775 393 1816 427
rect 1850 393 1866 427
rect 1280 345 1391 365
rect 1133 257 1233 279
rect 1280 257 1380 345
rect 1552 329 1733 379
rect 1775 373 1866 393
rect 1908 471 2054 487
rect 1908 437 1941 471
rect 1975 437 2054 471
rect 1908 417 2054 437
rect 2096 517 2196 543
rect 2096 417 2231 517
rect 1908 331 1951 417
rect 2131 396 2231 417
rect 2131 362 2177 396
rect 2211 362 2231 396
rect 1552 295 1572 329
rect 1606 295 1733 329
rect 1552 279 1733 295
rect 1633 257 1733 279
rect 1789 279 1951 331
rect 1993 335 2089 355
rect 1993 301 2009 335
rect 2043 301 2089 335
rect 1789 257 1889 279
rect 1993 267 2089 301
rect 537 147 637 173
rect 679 147 779 173
rect 835 147 935 173
rect 991 147 1091 173
rect 1133 147 1233 173
rect 1280 147 1380 173
rect 1993 237 2009 267
rect 1989 233 2009 237
rect 2043 233 2089 267
rect 1989 191 2089 233
rect 2131 328 2231 362
rect 2131 294 2177 328
rect 2211 294 2231 328
rect 2131 191 2231 294
rect 2273 351 2373 543
rect 2429 471 2529 543
rect 2429 437 2449 471
rect 2483 437 2529 471
rect 2429 417 2529 437
rect 2714 417 2814 443
rect 2889 417 2989 443
rect 2273 331 2387 351
rect 2273 297 2307 331
rect 2341 297 2387 331
rect 2273 263 2387 297
rect 2273 229 2307 263
rect 2341 229 2387 263
rect 2273 213 2387 229
rect 2287 191 2387 213
rect 2429 317 2814 417
rect 2874 385 2989 417
rect 2874 351 2894 385
rect 2928 351 2989 385
rect 2874 317 2989 351
rect 2429 191 2529 317
rect 2706 291 2806 317
rect 2885 291 2985 317
rect 2706 181 2806 207
rect 2885 115 2985 141
rect 87 81 187 107
rect 243 81 343 107
rect 1633 81 1733 107
rect 1789 81 1889 107
rect 1989 81 2089 107
rect 2131 81 2231 107
rect 2287 81 2387 107
rect 2429 81 2529 107
<< polycont >>
rect 264 455 298 489
rect 264 387 298 421
rect 128 319 162 353
rect 128 251 162 285
rect 851 550 885 584
rect 1012 550 1046 584
rect 555 408 589 442
rect 555 340 589 374
rect 699 371 733 405
rect 699 303 733 337
rect 1184 434 1218 468
rect 1011 365 1045 399
rect 1011 297 1045 331
rect 1184 366 1218 400
rect 1337 365 1371 399
rect 1816 461 1850 495
rect 1816 393 1850 427
rect 1941 437 1975 471
rect 2177 362 2211 396
rect 1572 295 1606 329
rect 2009 301 2043 335
rect 2009 233 2043 267
rect 2177 294 2211 328
rect 2449 437 2483 471
rect 2307 297 2341 331
rect 2307 229 2341 263
rect 2894 351 2928 385
<< locali >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2239 831
rect 2273 797 2335 831
rect 2369 797 2431 831
rect 2465 797 2527 831
rect 2561 797 2623 831
rect 2657 797 2719 831
rect 2753 797 2815 831
rect 2849 797 2911 831
rect 2945 797 3007 831
rect 3041 797 3072 831
rect 126 735 244 741
rect 126 701 132 735
rect 166 701 204 735
rect 238 701 244 735
rect 22 675 88 691
rect 22 641 38 675
rect 72 641 88 675
rect 22 583 88 641
rect 22 549 38 583
rect 72 549 88 583
rect 22 505 88 549
rect 126 679 244 701
rect 126 645 194 679
rect 228 645 244 679
rect 126 579 244 645
rect 126 545 194 579
rect 228 545 244 579
rect 280 727 568 761
rect 280 505 314 727
rect 22 489 314 505
rect 22 471 264 489
rect 22 166 76 471
rect 248 455 264 471
rect 298 455 314 489
rect 112 353 178 430
rect 248 421 314 455
rect 248 387 264 421
rect 298 387 314 421
rect 248 371 314 387
rect 350 675 400 691
rect 384 641 400 675
rect 350 583 400 641
rect 384 549 400 583
rect 350 430 400 549
rect 448 674 498 691
rect 448 640 464 674
rect 448 568 498 640
rect 534 638 568 727
rect 604 735 670 741
rect 604 701 610 735
rect 644 708 670 735
rect 604 674 620 701
rect 654 674 670 708
rect 706 727 1054 761
rect 706 638 740 727
rect 534 604 740 638
rect 776 674 810 691
rect 916 682 982 691
rect 916 648 932 682
rect 966 648 982 682
rect 916 640 982 648
rect 776 568 810 640
rect 448 534 810 568
rect 846 584 890 600
rect 846 550 851 584
rect 885 550 890 584
rect 846 534 890 550
rect 776 498 810 534
rect 539 442 647 498
rect 776 464 820 498
rect 350 424 455 430
rect 350 390 415 424
rect 449 390 455 424
rect 350 384 455 390
rect 539 408 555 442
rect 589 408 647 442
rect 112 319 128 353
rect 162 319 178 353
rect 112 285 178 319
rect 112 251 128 285
rect 162 251 178 285
rect 112 235 178 251
rect 350 199 404 384
rect 539 374 647 408
rect 539 340 555 374
rect 589 340 647 374
rect 539 324 647 340
rect 22 132 42 166
rect 22 99 76 132
rect 112 166 302 199
rect 112 132 198 166
rect 232 132 302 166
rect 112 113 302 132
rect 112 79 118 113
rect 152 79 190 113
rect 224 79 262 113
rect 296 79 302 113
rect 338 166 404 199
rect 338 132 354 166
rect 388 132 404 166
rect 338 99 404 132
rect 440 232 558 249
rect 440 198 492 232
rect 526 198 558 232
rect 440 113 558 198
rect 112 73 302 79
rect 440 79 446 113
rect 480 79 518 113
rect 552 79 558 113
rect 613 126 647 324
rect 683 405 749 421
rect 683 371 699 405
rect 733 371 749 405
rect 683 337 749 371
rect 683 303 699 337
rect 733 303 749 337
rect 683 162 749 303
rect 786 265 820 464
rect 856 430 890 534
rect 926 500 960 640
rect 1020 609 1054 727
rect 1090 735 1280 741
rect 1090 701 1096 735
rect 1130 701 1168 735
rect 1202 701 1240 735
rect 1274 701 1280 735
rect 1090 693 1280 701
rect 1090 659 1230 693
rect 1264 659 1280 693
rect 1090 645 1280 659
rect 1316 727 1522 761
rect 1316 609 1350 727
rect 1020 600 1350 609
rect 996 584 1350 600
rect 996 550 1012 584
rect 1046 575 1350 584
rect 1386 682 1452 691
rect 1386 648 1402 682
rect 1436 648 1452 682
rect 1046 550 1062 575
rect 996 536 1062 550
rect 1386 539 1452 648
rect 1488 655 1522 727
rect 1558 735 1748 751
rect 1558 701 1564 735
rect 1598 730 1636 735
rect 1608 701 1636 730
rect 1670 701 1708 735
rect 1742 701 1748 735
rect 1558 696 1574 701
rect 1608 696 1748 701
rect 1558 691 1748 696
rect 1886 735 1936 751
rect 1920 701 1936 735
rect 1886 660 1936 701
rect 1488 621 1850 655
rect 1098 505 1452 539
rect 1714 551 1730 585
rect 1764 551 1780 585
rect 1098 500 1132 505
rect 926 466 1132 500
rect 1714 469 1780 551
rect 856 424 1061 430
rect 856 390 895 424
rect 929 399 1061 424
rect 929 390 1011 399
rect 856 384 1011 390
rect 995 365 1011 384
rect 1045 365 1061 399
rect 995 331 1061 365
rect 995 297 1011 331
rect 1045 297 1061 331
rect 995 285 1061 297
rect 1098 329 1132 466
rect 1168 468 1780 469
rect 1168 434 1184 468
rect 1218 435 1780 468
rect 1218 434 1234 435
rect 1168 400 1234 434
rect 1168 366 1184 400
rect 1218 366 1234 400
rect 1168 365 1234 366
rect 1321 365 1337 399
rect 1371 365 1692 399
rect 1098 295 1572 329
rect 1606 295 1622 329
rect 786 232 840 265
rect 1098 249 1132 295
rect 1658 259 1692 365
rect 786 198 790 232
rect 824 198 840 232
rect 786 165 840 198
rect 930 232 1132 249
rect 930 198 946 232
rect 980 215 1132 232
rect 1168 225 1692 259
rect 980 198 996 215
rect 930 165 996 198
rect 1168 126 1202 225
rect 613 92 1202 126
rect 1432 169 1622 189
rect 1432 135 1572 169
rect 1606 135 1622 169
rect 1432 113 1622 135
rect 440 73 558 79
rect 1432 79 1438 113
rect 1472 79 1510 113
rect 1544 79 1582 113
rect 1616 79 1622 113
rect 1432 73 1622 79
rect 1658 87 1692 225
rect 1728 265 1780 435
rect 1816 495 1850 621
rect 1920 626 1936 660
rect 1886 585 1936 626
rect 1920 569 1936 585
rect 2097 735 2287 741
rect 2097 701 2103 735
rect 2137 701 2175 735
rect 2209 701 2247 735
rect 2281 701 2287 735
rect 2097 602 2287 701
rect 2454 735 2633 741
rect 2488 701 2526 735
rect 2560 701 2598 735
rect 2632 701 2633 735
rect 1920 551 2061 569
rect 1886 535 2061 551
rect 2097 568 2207 602
rect 2241 568 2287 602
rect 2097 535 2287 568
rect 2368 602 2418 635
rect 2368 568 2384 602
rect 2454 615 2633 701
rect 2454 581 2540 615
rect 2574 581 2633 615
rect 2755 735 2944 747
rect 2755 701 2760 735
rect 2794 701 2832 735
rect 2866 731 2904 735
rect 2878 701 2904 731
rect 2938 701 2944 735
rect 2755 697 2844 701
rect 2878 697 2944 701
rect 2755 651 2944 697
rect 2755 617 2844 651
rect 2878 617 2944 651
rect 2454 577 2633 581
rect 2669 585 2719 601
rect 2368 541 2418 568
rect 2703 551 2719 585
rect 1816 427 1850 461
rect 1816 351 1850 393
rect 1925 471 1991 487
rect 1925 437 1941 471
rect 1975 437 1991 471
rect 2027 471 2061 535
rect 2368 507 2569 541
rect 2027 437 2449 471
rect 2483 437 2499 471
rect 1925 424 1991 437
rect 1925 390 1951 424
rect 1985 390 1991 424
rect 1925 387 1991 390
rect 1816 335 2050 351
rect 1816 317 2009 335
rect 1993 301 2009 317
rect 2043 301 2050 335
rect 1993 267 2050 301
rect 1728 249 1794 265
rect 1728 215 1744 249
rect 1778 215 1794 249
rect 1728 157 1794 215
rect 1728 123 1744 157
rect 1778 123 1794 157
rect 1886 249 1952 265
rect 1886 215 1902 249
rect 1936 215 1952 249
rect 1993 233 2009 267
rect 2043 233 2050 267
rect 1993 217 2050 233
rect 1886 157 1952 215
rect 2086 157 2120 437
rect 2535 401 2569 507
rect 2161 396 2569 401
rect 2161 362 2177 396
rect 2211 367 2569 396
rect 2211 362 2227 367
rect 2161 328 2227 362
rect 2161 294 2177 328
rect 2211 294 2227 328
rect 2161 289 2227 294
rect 2291 297 2307 331
rect 2341 297 2357 331
rect 2291 263 2357 297
rect 2291 253 2307 263
rect 1886 123 1902 157
rect 1936 123 2120 157
rect 2156 229 2307 253
rect 2341 229 2357 263
rect 2156 219 2357 229
rect 2156 87 2190 219
rect 2524 199 2569 367
rect 2669 485 2719 551
rect 2703 451 2719 485
rect 2669 401 2719 451
rect 2755 569 2944 617
rect 2755 535 2844 569
rect 2878 535 2944 569
rect 2755 489 2944 535
rect 2755 455 2844 489
rect 2878 455 2944 489
rect 2755 439 2944 455
rect 2980 731 3047 747
rect 2980 697 3000 731
rect 3034 697 3047 731
rect 2980 651 3047 697
rect 2980 617 3000 651
rect 3034 617 3047 651
rect 2980 569 3047 617
rect 2980 535 3000 569
rect 3034 535 3047 569
rect 2980 489 3047 535
rect 2980 455 3000 489
rect 3034 455 3047 489
rect 2669 385 2944 401
rect 2669 351 2894 385
rect 2928 351 2944 385
rect 2669 335 2944 351
rect 2669 299 2711 335
rect 2645 266 2711 299
rect 2645 232 2661 266
rect 2695 232 2711 266
rect 2645 199 2711 232
rect 2747 283 2937 299
rect 2747 249 2840 283
rect 2874 249 2937 283
rect 1658 53 2190 87
rect 2226 166 2416 183
rect 2226 132 2242 166
rect 2276 132 2416 166
rect 2226 113 2416 132
rect 2226 79 2232 113
rect 2266 79 2304 113
rect 2338 79 2376 113
rect 2410 79 2416 113
rect 2524 166 2590 199
rect 2524 132 2540 166
rect 2574 132 2590 166
rect 2524 99 2590 132
rect 2747 183 2937 249
rect 2747 149 2840 183
rect 2874 149 2937 183
rect 2747 113 2937 149
rect 2980 283 3047 455
rect 2980 249 2996 283
rect 3030 249 3047 283
rect 2980 183 3047 249
rect 2980 149 2996 183
rect 3030 149 3047 183
rect 2980 133 3047 149
rect 2226 73 2416 79
rect 2747 79 2753 113
rect 2787 79 2825 113
rect 2859 79 2897 113
rect 2931 79 2937 113
rect 2747 73 2937 79
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3072 17
<< viali >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 895 797 929 831
rect 991 797 1025 831
rect 1087 797 1121 831
rect 1183 797 1217 831
rect 1279 797 1313 831
rect 1375 797 1409 831
rect 1471 797 1505 831
rect 1567 797 1601 831
rect 1663 797 1697 831
rect 1759 797 1793 831
rect 1855 797 1889 831
rect 1951 797 1985 831
rect 2047 797 2081 831
rect 2143 797 2177 831
rect 2239 797 2273 831
rect 2335 797 2369 831
rect 2431 797 2465 831
rect 2527 797 2561 831
rect 2623 797 2657 831
rect 2719 797 2753 831
rect 2815 797 2849 831
rect 2911 797 2945 831
rect 3007 797 3041 831
rect 132 701 166 735
rect 204 701 238 735
rect 610 708 644 735
rect 610 701 620 708
rect 620 701 644 708
rect 415 390 449 424
rect 118 79 152 113
rect 190 79 224 113
rect 262 79 296 113
rect 446 79 480 113
rect 518 79 552 113
rect 1096 701 1130 735
rect 1168 701 1202 735
rect 1240 701 1274 735
rect 1564 730 1598 735
rect 1564 701 1574 730
rect 1574 701 1598 730
rect 1636 701 1670 735
rect 1708 701 1742 735
rect 895 390 929 424
rect 1438 79 1472 113
rect 1510 79 1544 113
rect 1582 79 1616 113
rect 2103 701 2137 735
rect 2175 701 2209 735
rect 2247 701 2281 735
rect 2454 701 2488 735
rect 2526 701 2560 735
rect 2598 701 2632 735
rect 2760 701 2794 735
rect 2832 731 2866 735
rect 2832 701 2844 731
rect 2844 701 2866 731
rect 2904 701 2938 735
rect 1951 390 1985 424
rect 2232 79 2266 113
rect 2304 79 2338 113
rect 2376 79 2410 113
rect 2753 79 2787 113
rect 2825 79 2859 113
rect 2897 79 2931 113
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
rect 3007 -17 3041 17
<< metal1 >>
rect 0 831 3072 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2239 831
rect 2273 797 2335 831
rect 2369 797 2431 831
rect 2465 797 2527 831
rect 2561 797 2623 831
rect 2657 797 2719 831
rect 2753 797 2815 831
rect 2849 797 2911 831
rect 2945 797 3007 831
rect 3041 797 3072 831
rect 0 791 3072 797
rect 0 735 3072 763
rect 0 701 132 735
rect 166 701 204 735
rect 238 701 610 735
rect 644 701 1096 735
rect 1130 701 1168 735
rect 1202 701 1240 735
rect 1274 701 1564 735
rect 1598 701 1636 735
rect 1670 701 1708 735
rect 1742 701 2103 735
rect 2137 701 2175 735
rect 2209 701 2247 735
rect 2281 701 2454 735
rect 2488 701 2526 735
rect 2560 701 2598 735
rect 2632 701 2760 735
rect 2794 701 2832 735
rect 2866 701 2904 735
rect 2938 701 3072 735
rect 0 689 3072 701
rect 403 424 461 430
rect 403 390 415 424
rect 449 421 461 424
rect 883 424 941 430
rect 883 421 895 424
rect 449 393 895 421
rect 449 390 461 393
rect 403 384 461 390
rect 883 390 895 393
rect 929 421 941 424
rect 1939 424 1997 430
rect 1939 421 1951 424
rect 929 393 1951 421
rect 929 390 941 393
rect 883 384 941 390
rect 1939 390 1951 393
rect 1985 390 1997 424
rect 1939 384 1997 390
rect 0 113 3072 125
rect 0 79 118 113
rect 152 79 190 113
rect 224 79 262 113
rect 296 79 446 113
rect 480 79 518 113
rect 552 79 1438 113
rect 1472 79 1510 113
rect 1544 79 1582 113
rect 1616 79 2232 113
rect 2266 79 2304 113
rect 2338 79 2376 113
rect 2410 79 2753 113
rect 2787 79 2825 113
rect 2859 79 2897 113
rect 2931 79 3072 113
rect 0 51 3072 79
rect 0 17 3072 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3072 17
rect 0 -23 3072 -17
<< labels >>
rlabel comment s 0 0 0 0 4 dfrtp_1
flabel metal1 s 0 51 3072 125 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel metal1 s 0 0 3072 23 0 FreeSans 340 0 0 0 VNB
port 5 nsew ground bidirectional
flabel metal1 s 0 689 3072 763 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 791 3072 814 0 FreeSans 340 0 0 0 VPB
port 6 nsew power bidirectional
flabel locali s 703 168 737 202 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 607 464 641 498 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 3007 168 3041 202 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 3007 242 3041 276 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 3007 316 3041 350 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 3007 390 3041 424 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 3007 464 3041 498 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 3007 538 3041 572 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 3007 612 3041 646 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 3072 814
string GDS_END 948166
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string GDS_START 919000
string LEFclass CORE
string LEFsite unithv
string LEFsymmetry X Y
<< end >>
