magic
tech sky130A
magscale 1 2
timestamp 1676037725
<< nwell >>
rect -38 261 1142 582
<< pwell >>
rect 28 21 1078 203
rect 29 -17 63 21
<< locali >>
rect 474 332 524 425
rect 17 289 406 323
rect 17 215 142 289
rect 188 215 296 255
rect 340 215 406 289
rect 474 181 532 332
rect 662 215 841 255
rect 891 215 1087 255
rect 214 145 532 181
rect 214 129 280 145
rect 466 51 532 145
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 54 391 104 493
rect 138 427 188 527
rect 222 391 272 493
rect 306 427 356 527
rect 390 459 608 493
rect 390 391 440 459
rect 54 357 440 391
rect 558 359 608 459
rect 662 393 712 493
rect 746 427 796 527
rect 830 459 1048 493
rect 830 393 880 459
rect 662 357 880 393
rect 914 323 964 425
rect 590 289 964 323
rect 998 291 1048 459
rect 590 265 624 289
rect 566 199 624 265
rect 62 17 96 179
rect 130 95 180 179
rect 590 181 624 199
rect 590 145 972 181
rect 130 51 364 95
rect 398 17 432 111
rect 566 17 704 111
rect 738 51 804 145
rect 838 17 872 111
rect 906 51 972 145
rect 1006 17 1040 181
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
<< metal1 >>
rect 0 561 1104 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 0 496 1104 527
rect 0 17 1104 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
rect 0 -48 1104 -17
<< labels >>
rlabel locali s 662 215 841 255 6 A1_N
port 1 nsew signal input
rlabel locali s 891 215 1087 255 6 A2_N
port 2 nsew signal input
rlabel locali s 340 215 406 289 6 B1
port 3 nsew signal input
rlabel locali s 17 215 142 289 6 B1
port 3 nsew signal input
rlabel locali s 17 289 406 323 6 B1
port 3 nsew signal input
rlabel locali s 188 215 296 255 6 B2
port 4 nsew signal input
rlabel metal1 s 0 -48 1104 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 28 21 1078 203 6 VNB
port 6 nsew ground bidirectional
rlabel nwell s -38 261 1142 582 6 VPB
port 7 nsew power bidirectional
rlabel metal1 s 0 496 1104 592 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 466 51 532 145 6 Y
port 9 nsew signal output
rlabel locali s 214 129 280 145 6 Y
port 9 nsew signal output
rlabel locali s 214 145 532 181 6 Y
port 9 nsew signal output
rlabel locali s 474 181 532 332 6 Y
port 9 nsew signal output
rlabel locali s 474 332 524 425 6 Y
port 9 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1104 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 3950532
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3941734
<< end >>
