magic
tech sky130A
magscale 1 2
timestamp 1676037725
<< nwell >>
rect -38 261 774 582
<< pwell >>
rect 98 163 368 203
rect 1 27 729 163
rect 30 21 368 27
rect 30 -17 64 21
<< scnmos >>
rect 79 53 109 137
rect 176 47 206 177
rect 260 47 290 177
rect 357 53 387 137
rect 453 53 483 137
rect 537 53 567 137
rect 621 53 651 137
<< scpmoshvt >>
rect 79 297 109 381
rect 176 297 206 497
rect 260 297 290 497
rect 357 297 387 381
rect 453 297 483 381
rect 525 297 555 381
rect 621 297 651 381
<< ndiff >>
rect 124 137 176 177
rect 27 117 79 137
rect 27 83 35 117
rect 69 83 79 117
rect 27 53 79 83
rect 109 97 176 137
rect 109 63 126 97
rect 160 63 176 97
rect 109 53 176 63
rect 124 47 176 53
rect 206 120 260 177
rect 206 86 216 120
rect 250 86 260 120
rect 206 47 260 86
rect 290 137 342 177
rect 290 97 357 137
rect 290 63 303 97
rect 337 63 357 97
rect 290 53 357 63
rect 387 111 453 137
rect 387 77 397 111
rect 431 77 453 111
rect 387 53 453 77
rect 483 97 537 137
rect 483 63 493 97
rect 527 63 537 97
rect 483 53 537 63
rect 567 111 621 137
rect 567 77 577 111
rect 611 77 621 111
rect 567 53 621 77
rect 651 117 703 137
rect 651 83 661 117
rect 695 83 703 117
rect 651 53 703 83
rect 290 47 342 53
<< pdiff >>
rect 107 501 161 513
rect 107 467 119 501
rect 153 497 161 501
rect 305 501 358 513
rect 305 497 313 501
rect 153 467 176 497
rect 107 437 176 467
rect 124 381 176 437
rect 27 361 79 381
rect 27 327 35 361
rect 69 327 79 361
rect 27 297 79 327
rect 109 297 176 381
rect 206 349 260 497
rect 206 315 216 349
rect 250 315 260 349
rect 206 297 260 315
rect 290 467 313 497
rect 347 467 358 501
rect 290 437 358 467
rect 290 381 342 437
rect 290 297 357 381
rect 387 297 453 381
rect 483 297 525 381
rect 555 297 621 381
rect 651 348 703 381
rect 651 314 661 348
rect 695 314 703 348
rect 651 297 703 314
<< ndiffc >>
rect 35 83 69 117
rect 126 63 160 97
rect 216 86 250 120
rect 303 63 337 97
rect 397 77 431 111
rect 493 63 527 97
rect 577 77 611 111
rect 661 83 695 117
<< pdiffc >>
rect 119 467 153 501
rect 35 327 69 361
rect 216 315 250 349
rect 313 467 347 501
rect 661 314 695 348
<< poly >>
rect 176 497 206 523
rect 260 497 290 523
rect 79 381 109 407
rect 423 477 489 487
rect 423 443 439 477
rect 473 443 489 477
rect 423 433 489 443
rect 588 477 654 487
rect 588 443 604 477
rect 638 443 654 477
rect 588 433 654 443
rect 357 381 387 407
rect 453 381 483 433
rect 525 381 555 407
rect 621 381 651 433
rect 79 265 109 297
rect 25 249 109 265
rect 25 215 35 249
rect 69 215 109 249
rect 25 199 109 215
rect 79 137 109 199
rect 176 265 206 297
rect 260 265 290 297
rect 357 265 387 297
rect 176 249 302 265
rect 176 215 258 249
rect 292 215 302 249
rect 176 199 302 215
rect 357 249 411 265
rect 357 215 367 249
rect 401 215 411 249
rect 357 199 411 215
rect 176 177 206 199
rect 260 177 290 199
rect 79 27 109 53
rect 357 137 387 199
rect 453 137 483 297
rect 525 265 555 297
rect 525 249 579 265
rect 525 215 535 249
rect 569 215 579 249
rect 525 199 579 215
rect 537 137 567 199
rect 621 137 651 297
rect 176 21 206 47
rect 260 21 290 47
rect 357 27 387 53
rect 453 27 483 53
rect 537 27 567 53
rect 621 27 651 53
<< polycont >>
rect 439 443 473 477
rect 604 443 638 477
rect 35 215 69 249
rect 258 215 292 249
rect 367 215 401 249
rect 535 215 569 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 103 501 169 527
rect 103 467 119 501
rect 153 467 169 501
rect 296 501 363 527
rect 296 467 313 501
rect 347 467 363 501
rect 397 477 534 483
rect 397 443 439 477
rect 473 443 534 477
rect 102 399 343 433
rect 397 425 534 443
rect 572 443 604 477
rect 638 443 669 477
rect 102 378 153 399
rect 17 361 153 378
rect 288 391 343 399
rect 572 391 606 443
rect 17 327 35 361
rect 69 327 153 361
rect 17 321 153 327
rect 17 249 85 287
rect 17 215 35 249
rect 69 215 85 249
rect 119 181 153 321
rect 17 147 153 181
rect 187 349 250 365
rect 288 357 606 391
rect 187 315 216 349
rect 645 348 712 363
rect 645 323 661 348
rect 187 299 250 315
rect 284 314 661 323
rect 695 314 712 348
rect 187 158 221 299
rect 284 290 712 314
rect 283 289 712 290
rect 283 285 333 289
rect 283 284 331 285
rect 283 282 329 284
rect 283 280 326 282
rect 283 278 325 280
rect 283 276 324 278
rect 283 274 322 276
rect 283 271 320 274
rect 283 265 317 271
rect 258 249 317 265
rect 292 215 317 249
rect 351 249 464 255
rect 351 215 367 249
rect 401 215 464 249
rect 510 249 710 255
rect 510 215 535 249
rect 569 215 710 249
rect 258 199 317 215
rect 283 181 317 199
rect 17 117 70 147
rect 187 136 249 158
rect 283 147 611 181
rect 187 135 250 136
rect 17 83 35 117
rect 69 83 70 117
rect 194 120 250 135
rect 17 65 70 83
rect 126 97 160 113
rect 126 17 160 63
rect 194 86 216 120
rect 397 111 431 147
rect 194 52 250 86
rect 287 63 303 97
rect 337 63 363 97
rect 287 17 363 63
rect 577 111 611 147
rect 397 61 431 77
rect 477 63 493 97
rect 527 63 543 97
rect 477 17 543 63
rect 577 61 611 77
rect 645 83 661 117
rect 695 83 711 117
rect 645 17 711 83
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
flabel locali s 673 221 707 255 0 FreeSans 400 180 0 0 C
port 3 nsew signal input
flabel locali s 397 221 431 255 0 FreeSans 400 180 0 0 A
port 1 nsew signal input
flabel locali s 214 85 248 119 0 FreeSans 200 180 0 0 X
port 9 nsew signal output
flabel locali s 581 221 615 255 0 FreeSans 400 180 0 0 C
port 3 nsew signal input
flabel locali s 489 425 523 459 0 FreeSans 400 180 0 0 B
port 2 nsew signal input
flabel locali s 30 221 64 255 0 FreeSans 400 0 0 0 D_N
port 4 nsew signal input
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional abutment
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional abutment
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
rlabel comment s 0 0 0 0 4 or4b_2
rlabel metal1 s 0 -48 736 48 1 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 496 736 592 1 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 736 544
string GDS_END 1082032
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1075538
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 3.680 0.000 
<< end >>
