magic
tech sky130A
magscale 1 2
timestamp 1676037725
<< metal1 >>
tri 287 9440 321 9474 se
tri 317 9390 321 9394 ne
tri 2390 2540 2396 2546 ne
tri 2524 2540 2530 2546 nw
tri 9569 2540 9575 2546 ne
tri 9703 2540 9709 2546 nw
tri 1845 2490 1851 2496 se
tri 1979 2490 1985 2496 sw
tri 3519 2490 3525 2496 se
tri 3653 2490 3659 2496 sw
tri 8092 2490 8098 2496 se
tri 8228 2490 8234 2496 sw
tri 9764 2490 9770 2496 se
tri 9900 2490 9906 2496 sw
tri 245 1812 291 1858 sw
tri 2043 1812 2077 1846 se
tri 2129 1812 2163 1846 sw
rect 225 1760 3647 1812
rect 320 1680 9770 1732
tri 320 1646 354 1680 nw
tri 352 1383 386 1417 sw
rect 317 1331 14937 1383
<< metal2 >>
rect 12150 28507 12206 31368
tri 12206 28507 12226 28527 sw
rect 12150 28505 12226 28507
tri 12150 28429 12226 28505 ne
tri 12226 28429 12304 28507 sw
tri 12226 28351 12304 28429 ne
tri 12304 28351 12382 28429 sw
tri 12304 28273 12382 28351 ne
tri 12382 28273 12460 28351 sw
tri 12382 28217 12438 28273 ne
rect 12438 28239 12998 28273
tri 12998 28239 13032 28273 sw
rect 12438 28217 13032 28239
tri 12976 28161 13032 28217 ne
tri 13032 28161 13110 28239 sw
tri 13032 28083 13110 28161 ne
tri 13110 28083 13188 28161 sw
tri 13110 28061 13132 28083 ne
rect 13132 27538 13188 28083
tri 13132 27482 13188 27538 ne
tri 13188 27490 13258 27560 sw
rect 13188 27482 13258 27490
tri 13188 27412 13258 27482 ne
tri 13258 27412 13336 27490 sw
tri 14252 27477 14330 27555 se
rect 14330 27499 14393 27555
tri 14330 27477 14352 27499 nw
tri 13258 27334 13336 27412 ne
tri 13336 27334 13414 27412 sw
tri 14174 27399 14252 27477 se
tri 14252 27399 14330 27477 nw
tri 14109 27334 14174 27399 se
rect 14174 27334 14187 27399
tri 14187 27334 14252 27399 nw
tri 13336 27278 13392 27334 ne
rect 13392 27278 14131 27334
tri 14131 27278 14187 27334 nw
rect 321 9375 373 9390
rect 321 1986 352 9375
tri 352 9354 373 9375 nw
tri 715 3387 785 3457 se
rect 785 3387 915 3898
tri 1618 3844 1802 4028 se
rect 1802 3898 2265 4028
rect 5647 3904 6364 4028
tri 1802 3844 1856 3898 nw
rect 584 3257 915 3387
tri 1497 3723 1618 3844 se
rect 1618 3723 1627 3844
tri 524 2106 584 2166 se
rect 584 2106 714 3257
tri 714 3187 784 3257 nw
tri 714 2106 768 2160 sw
tri 1410 2106 1497 2193 se
rect 1497 2106 1627 3723
tri 1627 3669 1802 3844 nw
rect 2697 3319 2827 3898
tri 2827 3319 2852 3344 sw
rect 2697 3290 2852 3319
tri 2697 3135 2852 3290 ne
tri 2852 3135 3036 3319 sw
tri 2852 2951 3036 3135 ne
tri 3036 2951 3220 3135 sw
tri 3036 2897 3090 2951 ne
rect 1851 2401 1979 2496
tri 2396 2489 2447 2540 ne
tri 1851 2273 1979 2401 ne
tri 1979 2345 1981 2347 sw
rect 1979 2273 1981 2345
tri 1979 2271 1981 2273 ne
tri 1981 2271 2055 2345 sw
tri 1981 2197 2055 2271 ne
tri 2055 2197 2129 2271 sw
tri 1627 2106 1714 2193 sw
tri 2055 2175 2077 2197 ne
tri 321 1955 352 1986 ne
tri 352 1965 384 1997 sw
rect 352 1955 384 1965
tri 543 1958 577 1992 nw
tri 621 1958 655 1992 ne
tri 785 1958 819 1992 nw
tri 862 1958 896 1992 ne
tri 1390 1956 1426 1992 nw
tri 1528 1956 1564 1992 ne
tri 1694 1956 1730 1992 nw
tri 1811 1956 1847 1992 ne
tri 352 1953 354 1955 ne
tri 321 1551 354 1584 se
rect 354 1572 384 1955
rect 2077 1888 2129 2197
rect 2447 1652 2499 2540
tri 2499 2515 2524 2540 nw
tri 3003 2106 3090 2193 se
rect 3090 2106 3220 2951
rect 2790 1992 3220 2106
tri 2499 1652 2575 1728 sw
rect 354 1551 363 1572
tri 363 1551 384 1572 nw
rect 321 1372 352 1551
tri 352 1540 363 1551 nw
rect 2790 1478 2920 1992
tri 2920 1956 2956 1992 nw
rect 5647 1491 5978 3904
tri 5978 3769 6113 3904 nw
tri 7345 2106 7657 2418 se
rect 7657 2218 7787 3899
tri 7787 2218 7793 2224 sw
rect 7657 2106 7793 2218
tri 8505 2066 8589 2150 se
rect 8589 1992 8846 3903
tri 9575 2493 9622 2540 ne
tri 8846 2066 8936 2156 sw
tri 6933 1956 6969 1992 nw
tri 7197 1956 7233 1992 ne
tri 7363 1956 7399 1992 nw
tri 7627 1956 7663 1992 ne
tri 8635 1956 8671 1992 nw
tri 8899 1956 8935 1992 ne
tri 9065 1956 9101 1992 nw
tri 9329 1956 9365 1992 ne
tri 2790 1348 2920 1478 ne
rect 9622 1453 9674 2540
tri 9674 2511 9703 2540 nw
tri 10082 2106 10214 2238 se
rect 10214 2106 10736 3903
tri 10736 2106 10868 2238 sw
tri 11425 2106 11625 2306 se
rect 11625 2106 12079 3905
tri 12079 2106 12211 2238 sw
tri 12885 2106 13047 2268 se
rect 13047 2106 13513 3905
tri 13513 2106 13619 2212 sw
tri 10115 1956 10151 1992 nw
tri 10379 1956 10415 1992 ne
tri 10545 1956 10581 1992 nw
tri 10809 1956 10845 1992 ne
tri 11458 1956 11494 1992 nw
tri 11722 1956 11758 1992 ne
tri 11888 1956 11924 1992 nw
tri 12152 1956 12188 1992 ne
tri 12892 1956 12928 1992 nw
tri 13156 1956 13192 1992 ne
tri 13322 1956 13358 1992 nw
tri 13586 1956 13622 1992 ne
tri 14589 1732 14623 1766 se
tri 10180 1646 10214 1680 ne
tri 2920 1354 2988 1422 sw
tri 9622 1401 9674 1453 ne
tri 9674 1411 9738 1475 sw
rect 9674 1401 9738 1411
tri 9674 1354 9721 1401 ne
rect 9721 1367 9738 1401
tri 9738 1367 9782 1411 sw
tri 10155 1367 10214 1426 se
rect 10214 1404 10266 1680
tri 10266 1651 10295 1680 nw
tri 14675 1652 14703 1680 se
tri 14755 1543 14783 1571 se
tri 14835 1463 14863 1491 se
rect 10214 1367 10229 1404
tri 10229 1367 10266 1404 nw
tri 14915 1383 14943 1411 se
rect 9721 1354 10177 1367
rect 2920 1348 2988 1354
tri 2920 1280 2988 1348 ne
tri 2988 1280 3062 1354 sw
tri 9721 1315 9760 1354 ne
rect 9760 1315 10177 1354
tri 10177 1315 10229 1367 nw
tri 2988 1206 3062 1280 ne
tri 3062 1206 3136 1280 sw
tri 14470 1206 14506 1242 se
tri 3062 1154 3114 1206 ne
rect 3114 1154 14506 1206
tri 14488 1136 14506 1154 ne
<< metal3 >>
rect 14395 27494 14567 27560
tri 14395 27388 14501 27494 ne
rect 14501 1286 14567 27494
use sky130_fd_io__nfet_con_diff_wo_abt_270v2  sky130_fd_io__nfet_con_diff_wo_abt_270v2_0
timestamp 1676037725
transform -1 0 15088 0 -1 8404
box 0 423 15173 5493
use sky130_fd_io__tk_em2o_cdns_55959141808653  sky130_fd_io__tk_em2o_cdns_55959141808653_0
timestamp 1676037725
transform 0 -1 12892 1 0 1584
box 0 0 1 1
use sky130_fd_io__tk_em2o_cdns_55959141808653  sky130_fd_io__tk_em2o_cdns_55959141808653_1
timestamp 1676037725
transform 0 -1 11458 1 0 1584
box 0 0 1 1
use sky130_fd_io__tk_em2o_cdns_55959141808653  sky130_fd_io__tk_em2o_cdns_55959141808653_2
timestamp 1676037725
transform 0 -1 10115 1 0 1584
box 0 0 1 1
use sky130_fd_io__tk_em2o_cdns_55959141808653  sky130_fd_io__tk_em2o_cdns_55959141808653_3
timestamp 1676037725
transform 0 -1 8635 1 0 1584
box 0 0 1 1
use sky130_fd_io__tk_em2o_cdns_55959141808653  sky130_fd_io__tk_em2o_cdns_55959141808653_4
timestamp 1676037725
transform 0 -1 6933 1 0 1584
box 0 0 1 1
use sky130_fd_io__tk_em2o_cdns_55959141808653  sky130_fd_io__tk_em2o_cdns_55959141808653_5
timestamp 1676037725
transform 0 -1 13322 1 0 1584
box 0 0 1 1
use sky130_fd_io__tk_em2o_cdns_55959141808653  sky130_fd_io__tk_em2o_cdns_55959141808653_6
timestamp 1676037725
transform 0 -1 10975 1 0 1584
box 0 0 1 1
use sky130_fd_io__tk_em2o_cdns_55959141808653  sky130_fd_io__tk_em2o_cdns_55959141808653_7
timestamp 1676037725
transform 0 -1 9495 1 0 1584
box 0 0 1 1
use sky130_fd_io__tk_em2o_cdns_55959141808653  sky130_fd_io__tk_em2o_cdns_55959141808653_8
timestamp 1676037725
transform 0 -1 12318 1 0 1584
box 0 0 1 1
use sky130_fd_io__tk_em2o_cdns_55959141808653  sky130_fd_io__tk_em2o_cdns_55959141808653_9
timestamp 1676037725
transform 0 -1 7793 1 0 1584
box 0 0 1 1
use sky130_fd_io__tk_em2o_cdns_55959141808653  sky130_fd_io__tk_em2o_cdns_55959141808653_10
timestamp 1676037725
transform 0 -1 1977 1 0 1584
box 0 0 1 1
use sky130_fd_io__tk_em2o_cdns_55959141808653  sky130_fd_io__tk_em2o_cdns_55959141808653_11
timestamp 1676037725
transform 0 -1 1694 1 0 1584
box 0 0 1 1
use sky130_fd_io__tk_em2o_cdns_55959141808653  sky130_fd_io__tk_em2o_cdns_55959141808653_12
timestamp 1676037725
transform 0 1 413 1 0 1584
box 0 0 1 1
use sky130_fd_io__tk_em2o_cdns_55959141808653  sky130_fd_io__tk_em2o_cdns_55959141808653_13
timestamp 1676037725
transform 0 1 896 1 0 1584
box 0 0 1 1
use sky130_fd_io__tk_em2s_cdns_55959141808652  sky130_fd_io__tk_em2s_cdns_55959141808652_0
timestamp 1676037725
transform 0 -1 11888 1 0 1584
box 0 0 1 1
use sky130_fd_io__tk_em2s_cdns_55959141808652  sky130_fd_io__tk_em2s_cdns_55959141808652_1
timestamp 1676037725
transform 0 -1 7363 1 0 1584
box 0 0 1 1
use sky130_fd_io__tk_em2s_cdns_55959141808652  sky130_fd_io__tk_em2s_cdns_55959141808652_2
timestamp 1676037725
transform 0 -1 10545 1 0 1584
box 0 0 1 1
use sky130_fd_io__tk_em2s_cdns_55959141808652  sky130_fd_io__tk_em2s_cdns_55959141808652_3
timestamp 1676037725
transform 0 -1 9065 1 0 1584
box 0 0 1 1
use sky130_fd_io__tk_em2s_cdns_55959141808652  sky130_fd_io__tk_em2s_cdns_55959141808652_4
timestamp 1676037725
transform 0 -1 13752 1 0 1584
box 0 0 1 1
use sky130_fd_io__tk_em2s_cdns_55959141808652  sky130_fd_io__tk_em2s_cdns_55959141808652_5
timestamp 1676037725
transform 0 -1 1390 1 0 1584
box 0 0 1 1
use sky130_fd_io__tk_em2s_cdns_55959141808652  sky130_fd_io__tk_em2s_cdns_55959141808652_6
timestamp 1676037725
transform 0 1 655 1 0 1584
box 0 0 1 1
use sky130_fd_pr__res_generic_po__example_5595914180838  sky130_fd_pr__res_generic_po__example_5595914180838_0
timestamp 1676037725
transform 1 0 336 0 1 9367
box 15 17 2025 18
use sky130_fd_pr__via_pol1_centered__example_559591418081  sky130_fd_pr__via_pol1_centered__example_559591418081_0
timestamp 1676037725
transform -1 0 2461 0 -1 9417
box 0 0 1 1
use sky130_fd_pr__via_pol1_centered__example_559591418081  sky130_fd_pr__via_pol1_centered__example_559591418081_1
timestamp 1676037725
transform 1 0 251 0 -1 9417
box 0 0 1 1
<< properties >>
string GDS_END 46281392
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 46246244
<< end >>
