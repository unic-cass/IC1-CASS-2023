magic
tech sky130B
magscale 1 2
timestamp 1676037725
<< poly >>
rect 4432 33100 4566 33116
rect 4432 33066 4448 33100
rect 4482 33066 4516 33100
rect 4550 33066 4566 33100
rect 4432 33050 4566 33066
rect 5724 33100 5858 33116
rect 5724 33066 5740 33100
rect 5774 33066 5808 33100
rect 5842 33066 5858 33100
rect 5724 33050 5858 33066
rect 7720 33100 7854 33116
rect 7720 33066 7736 33100
rect 7770 33066 7804 33100
rect 7838 33066 7854 33100
rect 7720 33050 7854 33066
rect 9014 33100 9148 33116
rect 9014 33066 9030 33100
rect 9064 33066 9098 33100
rect 9132 33066 9148 33100
rect 9014 33050 9148 33066
rect 9526 33100 9660 33116
rect 9526 33066 9542 33100
rect 9576 33066 9610 33100
rect 9644 33066 9660 33100
rect 9526 33050 9660 33066
rect 10816 33100 10950 33116
rect 10816 33066 10832 33100
rect 10866 33066 10900 33100
rect 10934 33066 10950 33100
rect 10816 33050 10950 33066
rect 11331 33100 11465 33116
rect 11331 33066 11347 33100
rect 11381 33066 11415 33100
rect 11449 33066 11465 33100
rect 11331 33050 11465 33066
rect 12625 33100 12759 33116
rect 12625 33066 12641 33100
rect 12675 33066 12709 33100
rect 12743 33066 12759 33100
rect 12625 33050 12759 33066
rect 13132 33100 13266 33116
rect 13132 33066 13148 33100
rect 13182 33066 13216 33100
rect 13250 33066 13266 33100
rect 13132 33050 13266 33066
rect 14426 33100 14560 33116
rect 14426 33066 14442 33100
rect 14476 33066 14510 33100
rect 14544 33066 14560 33100
rect 14426 33050 14560 33066
rect 14940 33100 15074 33116
rect 14940 33066 14956 33100
rect 14990 33066 15024 33100
rect 15058 33066 15074 33100
rect 14940 33050 15074 33066
rect 16230 33100 16364 33116
rect 16230 33066 16246 33100
rect 16280 33066 16314 33100
rect 16348 33066 16364 33100
rect 16230 33050 16364 33066
<< polycont >>
rect 4448 33066 4482 33100
rect 4516 33066 4550 33100
rect 5740 33066 5774 33100
rect 5808 33066 5842 33100
rect 7736 33066 7770 33100
rect 7804 33066 7838 33100
rect 9030 33066 9064 33100
rect 9098 33066 9132 33100
rect 9542 33066 9576 33100
rect 9610 33066 9644 33100
rect 10832 33066 10866 33100
rect 10900 33066 10934 33100
rect 11347 33066 11381 33100
rect 11415 33066 11449 33100
rect 12641 33066 12675 33100
rect 12709 33066 12743 33100
rect 13148 33066 13182 33100
rect 13216 33066 13250 33100
rect 14442 33066 14476 33100
rect 14510 33066 14544 33100
rect 14956 33066 14990 33100
rect 15024 33066 15058 33100
rect 16246 33066 16280 33100
rect 16314 33066 16348 33100
<< locali >>
rect 4432 33404 4566 33418
rect 4432 33370 4444 33404
rect 4478 33370 4520 33404
rect 4554 33370 4566 33404
rect 4432 33100 4566 33370
rect 4432 33066 4448 33100
rect 4482 33066 4516 33100
rect 4550 33066 4566 33100
rect 4432 33050 4566 33066
rect 5724 33404 5858 33418
rect 5724 33370 5736 33404
rect 5770 33370 5812 33404
rect 5846 33370 5858 33404
rect 5724 33100 5858 33370
rect 5724 33066 5740 33100
rect 5774 33066 5808 33100
rect 5842 33066 5858 33100
rect 5724 33050 5858 33066
rect 7720 33404 7854 33418
rect 7720 33370 7732 33404
rect 7766 33370 7808 33404
rect 7842 33370 7854 33404
rect 7720 33100 7854 33370
rect 7720 33066 7736 33100
rect 7770 33066 7804 33100
rect 7838 33066 7854 33100
rect 7720 33050 7854 33066
rect 9014 33404 9148 33418
rect 9014 33370 9026 33404
rect 9060 33370 9102 33404
rect 9136 33370 9148 33404
rect 9014 33100 9148 33370
rect 9014 33066 9030 33100
rect 9064 33066 9098 33100
rect 9132 33066 9148 33100
rect 9014 33050 9148 33066
rect 9526 33404 9660 33418
rect 9526 33370 9538 33404
rect 9572 33370 9614 33404
rect 9648 33370 9660 33404
rect 9526 33100 9660 33370
rect 9526 33066 9542 33100
rect 9576 33066 9610 33100
rect 9644 33066 9660 33100
rect 9526 33050 9660 33066
rect 10816 33404 10950 33418
rect 10816 33370 10828 33404
rect 10862 33370 10904 33404
rect 10938 33370 10950 33404
rect 10816 33100 10950 33370
rect 10816 33066 10832 33100
rect 10866 33066 10900 33100
rect 10934 33066 10950 33100
rect 10816 33050 10950 33066
rect 11331 33404 11465 33418
rect 11331 33370 11343 33404
rect 11377 33370 11419 33404
rect 11453 33370 11465 33404
rect 11331 33100 11465 33370
rect 11331 33066 11347 33100
rect 11381 33066 11415 33100
rect 11449 33066 11465 33100
rect 11331 33050 11465 33066
rect 12625 33404 12759 33418
rect 12625 33370 12637 33404
rect 12671 33370 12713 33404
rect 12747 33370 12759 33404
rect 12625 33100 12759 33370
rect 12625 33066 12641 33100
rect 12675 33066 12709 33100
rect 12743 33066 12759 33100
rect 12625 33050 12759 33066
rect 13132 33404 13266 33418
rect 13132 33370 13144 33404
rect 13178 33370 13220 33404
rect 13254 33370 13266 33404
rect 13132 33100 13266 33370
rect 13132 33066 13148 33100
rect 13182 33066 13216 33100
rect 13250 33066 13266 33100
rect 13132 33050 13266 33066
rect 14426 33404 14560 33418
rect 14426 33370 14438 33404
rect 14472 33370 14514 33404
rect 14548 33370 14560 33404
rect 14426 33100 14560 33370
rect 14426 33066 14442 33100
rect 14476 33066 14510 33100
rect 14544 33066 14560 33100
rect 14426 33050 14560 33066
rect 14940 33404 15074 33418
rect 14940 33370 14952 33404
rect 14986 33370 15028 33404
rect 15062 33370 15074 33404
rect 14940 33100 15074 33370
rect 14940 33066 14956 33100
rect 14990 33066 15024 33100
rect 15058 33066 15074 33100
rect 14940 33050 15074 33066
rect 16230 33404 16364 33418
rect 16230 33370 16242 33404
rect 16276 33370 16318 33404
rect 16352 33370 16364 33404
rect 16230 33100 16364 33370
rect 16230 33066 16246 33100
rect 16280 33066 16314 33100
rect 16348 33066 16364 33100
rect 16230 33050 16364 33066
<< viali >>
rect 4444 33370 4478 33404
rect 4520 33370 4554 33404
rect 5736 33370 5770 33404
rect 5812 33370 5846 33404
rect 7732 33370 7766 33404
rect 7808 33370 7842 33404
rect 9026 33370 9060 33404
rect 9102 33370 9136 33404
rect 9538 33370 9572 33404
rect 9614 33370 9648 33404
rect 10828 33370 10862 33404
rect 10904 33370 10938 33404
rect 11343 33370 11377 33404
rect 11419 33370 11453 33404
rect 12637 33370 12671 33404
rect 12713 33370 12747 33404
rect 13144 33370 13178 33404
rect 13220 33370 13254 33404
rect 14438 33370 14472 33404
rect 14514 33370 14548 33404
rect 14952 33370 14986 33404
rect 15028 33370 15062 33404
rect 16242 33370 16276 33404
rect 16318 33370 16352 33404
<< metal1 >>
rect 12043 35241 12466 35287
rect 10299 35210 10429 35214
rect 10299 35158 10305 35210
rect 10357 35158 10371 35210
rect 10423 35158 10429 35210
rect 10299 35154 10429 35158
rect 12043 35130 12125 35241
rect 12193 35207 12323 35211
rect 12193 35155 12199 35207
rect 12251 35155 12265 35207
rect 12317 35155 12323 35207
rect 12193 35151 12323 35155
rect 12384 35130 12466 35241
rect 4848 35071 4978 35100
rect 4848 35019 4854 35071
rect 4906 35019 4920 35071
rect 4972 35019 4978 35071
rect 4848 34990 4978 35019
rect 2910 34926 3054 34932
rect 2962 34874 3002 34926
rect 2910 34826 3054 34874
rect 1930 34667 1936 34783
rect 2052 34667 2058 34783
rect 2099 34727 2105 34783
rect 1930 33356 2058 34667
rect 1930 33240 1936 33356
rect 2052 33240 2058 33356
rect 2098 34667 2105 34727
rect 2221 34667 2227 34783
rect 2962 34774 3002 34826
rect 2910 34726 3054 34774
rect 2962 34674 3002 34726
rect 2910 34668 3054 34674
rect 2098 33356 2227 34667
rect 5278 34465 5408 34592
rect 10729 34545 10859 34592
rect 10729 34493 10736 34545
rect 10788 34493 10800 34545
rect 10852 34493 10859 34545
rect 11763 34545 11893 34592
rect 11763 34493 11770 34545
rect 11822 34493 11834 34545
rect 11886 34493 11893 34545
rect 5278 34413 5285 34465
rect 5337 34413 5349 34465
rect 5401 34413 5408 34465
rect 2098 33325 2105 33356
rect 2099 33240 2105 33325
rect 2221 33240 2227 33356
rect 3857 33404 5858 33433
rect 3857 33370 4444 33404
rect 4478 33370 4520 33404
rect 4554 33370 5736 33404
rect 5770 33370 5812 33404
rect 5846 33370 5858 33404
rect 3857 33355 5858 33370
rect 7719 33420 7902 33433
rect 7719 33368 7725 33420
rect 7777 33368 7789 33420
rect 7841 33404 7902 33420
rect 7842 33370 7902 33404
rect 7841 33368 7902 33370
rect 7719 33355 7902 33368
rect 8930 33421 9148 33433
rect 8930 33369 8936 33421
rect 8988 33369 9000 33421
rect 9052 33404 9148 33421
rect 9060 33370 9102 33404
rect 9136 33370 9148 33404
rect 9052 33369 9148 33370
rect 8930 33355 9148 33369
rect 9500 33421 9656 33433
rect 9500 33369 9532 33421
rect 9584 33369 9596 33421
rect 9648 33418 9656 33421
rect 11091 33420 16551 33433
rect 9648 33369 9660 33418
rect 9500 33356 9660 33369
rect 10816 33404 10950 33418
rect 10816 33370 10828 33404
rect 10862 33370 10904 33404
rect 10938 33370 10950 33404
rect 10816 33356 10950 33370
rect 11091 33404 16300 33420
rect 11091 33370 11343 33404
rect 11377 33370 11419 33404
rect 11453 33370 12637 33404
rect 12671 33370 12713 33404
rect 12747 33370 13144 33404
rect 13178 33370 13220 33404
rect 13254 33370 14438 33404
rect 14472 33370 14514 33404
rect 14548 33370 14952 33404
rect 14986 33370 15028 33404
rect 15062 33370 16242 33404
rect 16276 33370 16300 33404
rect 11091 33368 16300 33370
rect 16352 33368 16365 33420
rect 16417 33368 16429 33420
rect 16481 33368 16493 33420
rect 16545 33368 16551 33420
rect 9500 33355 9656 33356
rect 11091 33355 16551 33368
rect 23032 32105 23084 32111
rect 23032 32041 23084 32053
rect 23032 31142 23084 31989
rect 23032 31078 23084 31090
rect 23032 31020 23084 31026
tri 3235 30281 3307 30353 sw
rect 3235 30275 3347 30281
rect 3235 30223 3268 30275
rect 3320 30223 3347 30275
rect 3235 30147 3347 30223
rect 3235 30095 3268 30147
rect 3320 30095 3347 30147
rect 3235 30019 3347 30095
rect 3235 29967 3268 30019
rect 3320 29967 3347 30019
rect 3235 29891 3347 29967
rect 3235 29839 3268 29891
rect 3320 29839 3347 29891
rect 3235 29763 3347 29839
rect 3235 29711 3268 29763
rect 3320 29711 3347 29763
rect 3235 29635 3347 29711
rect 3235 29583 3268 29635
rect 3320 29583 3347 29635
rect 3235 29506 3347 29583
rect 3235 29454 3268 29506
rect 3320 29454 3347 29506
rect 3235 29377 3347 29454
rect 3235 29325 3268 29377
rect 3320 29325 3347 29377
rect 3235 29248 3347 29325
rect 3235 29196 3268 29248
rect 3320 29196 3347 29248
rect 3235 29119 3347 29196
rect 3235 29067 3268 29119
rect 3320 29067 3347 29119
rect 3235 28990 3347 29067
rect 3235 28938 3268 28990
rect 3320 28938 3347 28990
rect 3235 28861 3347 28938
rect 3235 28809 3268 28861
rect 3320 28809 3347 28861
rect 3235 28732 3347 28809
rect 3235 28680 3268 28732
rect 3320 28680 3347 28732
rect 3235 28603 3347 28680
rect 3235 28551 3268 28603
rect 3320 28551 3347 28603
rect 3235 28474 3347 28551
rect 3235 28422 3268 28474
rect 3320 28422 3347 28474
rect 3235 28345 3347 28422
rect 3235 28293 3268 28345
rect 3320 28293 3347 28345
rect 3235 28216 3347 28293
rect 3235 28164 3268 28216
rect 3320 28164 3347 28216
rect 3235 28087 3347 28164
rect 3235 28035 3268 28087
rect 3320 28035 3347 28087
rect 3235 27958 3347 28035
rect 3235 27906 3268 27958
rect 3320 27906 3347 27958
rect 3235 27829 3347 27906
rect 3235 27777 3268 27829
rect 3320 27777 3347 27829
rect 3235 27700 3347 27777
rect 3235 27648 3268 27700
rect 3320 27648 3347 27700
rect 3235 27571 3347 27648
rect 3235 27519 3268 27571
rect 3320 27519 3347 27571
rect 3235 27442 3347 27519
rect 3235 27390 3268 27442
rect 3320 27390 3347 27442
rect 3235 27313 3347 27390
rect 3235 27261 3268 27313
rect 3320 27261 3347 27313
rect 3235 27184 3347 27261
rect 3235 27132 3268 27184
rect 3320 27132 3347 27184
rect 3235 27055 3347 27132
rect 3235 27003 3268 27055
rect 3320 27003 3347 27055
rect 3235 26926 3347 27003
rect 3235 26874 3268 26926
rect 3320 26874 3347 26926
rect 3235 26797 3347 26874
rect 3235 26745 3268 26797
rect 3320 26745 3347 26797
rect 3235 26668 3347 26745
rect 3235 26616 3268 26668
rect 3320 26616 3347 26668
rect 3235 26539 3347 26616
rect 3235 26487 3268 26539
rect 3320 26487 3347 26539
rect 3235 26410 3347 26487
rect 3235 26358 3268 26410
rect 3320 26358 3347 26410
rect 3235 26281 3347 26358
rect 3235 26229 3268 26281
rect 3320 26229 3347 26281
rect 3235 26152 3347 26229
rect 3235 26100 3268 26152
rect 3320 26100 3347 26152
rect 3235 26023 3347 26100
rect 3235 25971 3268 26023
rect 3320 25971 3347 26023
rect 3235 25894 3347 25971
rect 3235 25842 3268 25894
rect 3320 25842 3347 25894
rect 3235 25765 3347 25842
rect 3235 25713 3268 25765
rect 3320 25713 3347 25765
rect 3235 25636 3347 25713
rect 3235 25584 3268 25636
rect 3320 25584 3347 25636
rect 3235 25507 3347 25584
rect 3235 25455 3268 25507
rect 3320 25455 3347 25507
rect 3235 25378 3347 25455
rect 3235 25326 3268 25378
rect 3320 25326 3347 25378
rect 3235 25249 3347 25326
rect 3235 25197 3268 25249
rect 3320 25197 3347 25249
rect 3235 25120 3347 25197
rect 3235 25068 3268 25120
rect 3320 25068 3347 25120
rect 3235 24991 3347 25068
rect 3235 24939 3268 24991
rect 3320 24939 3347 24991
rect 3235 24862 3347 24939
rect 3235 24810 3268 24862
rect 3320 24810 3347 24862
rect 3235 24733 3347 24810
rect 3235 24681 3268 24733
rect 3320 24681 3347 24733
rect 3235 24604 3347 24681
rect 3235 24552 3268 24604
rect 3320 24552 3347 24604
rect 3235 24475 3347 24552
rect 3235 24423 3268 24475
rect 3320 24423 3347 24475
rect 3235 24346 3347 24423
rect 3954 24513 3960 24565
rect 4012 24513 4026 24565
rect 4078 24513 4092 24565
rect 4144 24513 4158 24565
rect 4210 24513 4224 24565
rect 4276 24513 4289 24565
rect 4341 24513 4354 24565
rect 4406 24513 4419 24565
rect 4471 24513 4484 24565
rect 4536 24513 4542 24565
rect 3954 24449 4542 24513
rect 3954 24397 3960 24449
rect 4012 24397 4026 24449
rect 4078 24397 4092 24449
rect 4144 24397 4158 24449
rect 4210 24397 4224 24449
rect 4276 24397 4289 24449
rect 4341 24397 4354 24449
rect 4406 24397 4419 24449
rect 4471 24397 4484 24449
rect 4536 24397 4542 24449
rect 5762 24513 5768 24565
rect 5820 24513 5833 24565
rect 5885 24513 5898 24565
rect 5950 24513 5963 24565
rect 6015 24513 6028 24565
rect 6080 24513 6093 24565
rect 6145 24513 6158 24565
rect 6210 24513 6223 24565
rect 6275 24513 6287 24565
rect 6339 24513 6345 24565
rect 5762 24449 6345 24513
rect 5762 24397 5768 24449
rect 5820 24397 5833 24449
rect 5885 24397 5898 24449
rect 5950 24397 5963 24449
rect 6015 24397 6028 24449
rect 6080 24397 6093 24449
rect 6145 24397 6158 24449
rect 6210 24397 6223 24449
rect 6275 24397 6287 24449
rect 6339 24397 6345 24449
rect 7241 24513 7247 24565
rect 7299 24513 7312 24565
rect 7364 24513 7377 24565
rect 7429 24513 7442 24565
rect 7494 24513 7507 24565
rect 7559 24513 7572 24565
rect 7624 24513 7637 24565
rect 7689 24513 7701 24565
rect 7753 24513 7765 24565
rect 7817 24513 7823 24565
rect 7241 24449 7823 24513
rect 7241 24397 7247 24449
rect 7299 24397 7312 24449
rect 7364 24397 7377 24449
rect 7429 24397 7442 24449
rect 7494 24397 7507 24449
rect 7559 24397 7572 24449
rect 7624 24397 7637 24449
rect 7689 24397 7701 24449
rect 7753 24397 7765 24449
rect 7817 24397 7823 24449
rect 9045 24513 9051 24565
rect 9103 24513 9116 24565
rect 9168 24513 9181 24565
rect 9233 24513 9246 24565
rect 9298 24513 9311 24565
rect 9363 24513 9376 24565
rect 9428 24513 9441 24565
rect 9493 24513 9506 24565
rect 9558 24513 9570 24565
rect 9622 24513 9628 24565
rect 9045 24449 9628 24513
rect 9045 24397 9051 24449
rect 9103 24397 9116 24449
rect 9168 24397 9181 24449
rect 9233 24397 9246 24449
rect 9298 24397 9311 24449
rect 9363 24397 9376 24449
rect 9428 24397 9441 24449
rect 9493 24397 9506 24449
rect 9558 24397 9570 24449
rect 9622 24397 9628 24449
rect 10849 24513 10855 24565
rect 10907 24513 10920 24565
rect 10972 24513 10985 24565
rect 11037 24513 11050 24565
rect 11102 24513 11115 24565
rect 11167 24513 11180 24565
rect 11232 24513 11245 24565
rect 11297 24513 11309 24565
rect 11361 24513 11373 24565
rect 11425 24513 11431 24565
rect 10849 24449 11431 24513
rect 10849 24397 10855 24449
rect 10907 24397 10920 24449
rect 10972 24397 10985 24449
rect 11037 24397 11050 24449
rect 11102 24397 11115 24449
rect 11167 24397 11180 24449
rect 11232 24397 11245 24449
rect 11297 24397 11309 24449
rect 11361 24397 11373 24449
rect 11425 24397 11431 24449
rect 12648 24513 12654 24565
rect 12706 24513 12720 24565
rect 12772 24513 12786 24565
rect 12838 24513 12852 24565
rect 12904 24513 12917 24565
rect 12969 24513 12982 24565
rect 13034 24513 13047 24565
rect 13099 24513 13112 24565
rect 13164 24513 13177 24565
rect 13229 24513 13235 24565
rect 12648 24449 13235 24513
rect 12648 24397 12654 24449
rect 12706 24397 12720 24449
rect 12772 24397 12786 24449
rect 12838 24397 12852 24449
rect 12904 24397 12917 24449
rect 12969 24397 12982 24449
rect 13034 24397 13047 24449
rect 13099 24397 13112 24449
rect 13164 24397 13177 24449
rect 13229 24397 13235 24449
rect 14457 24511 14463 24563
rect 14515 24511 14528 24563
rect 14580 24511 14593 24563
rect 14645 24511 14658 24563
rect 14710 24511 14723 24563
rect 14775 24511 14788 24563
rect 14840 24511 14853 24563
rect 14905 24511 14917 24563
rect 14969 24511 14981 24563
rect 15033 24511 15039 24563
rect 14457 24447 15039 24511
rect 14457 24395 14463 24447
rect 14515 24395 14528 24447
rect 14580 24395 14593 24447
rect 14645 24395 14658 24447
rect 14710 24395 14723 24447
rect 14775 24395 14788 24447
rect 14840 24395 14853 24447
rect 14905 24395 14917 24447
rect 14969 24395 14981 24447
rect 15033 24395 15039 24447
rect 16261 24513 16267 24565
rect 16319 24513 16334 24565
rect 16386 24513 16401 24565
rect 16453 24513 16467 24565
rect 16519 24513 16533 24565
rect 16585 24513 16599 24565
rect 16651 24513 16665 24565
rect 16717 24513 16731 24565
rect 16783 24513 16797 24565
rect 16849 24513 16855 24565
rect 16261 24449 16855 24513
rect 16261 24397 16267 24449
rect 16319 24397 16334 24449
rect 16386 24397 16401 24449
rect 16453 24397 16467 24449
rect 16519 24397 16533 24449
rect 16585 24397 16599 24449
rect 16651 24397 16665 24449
rect 16717 24397 16731 24449
rect 16783 24397 16797 24449
rect 16849 24397 16855 24449
rect 3235 24294 3268 24346
rect 3320 24294 3347 24346
rect 3235 24217 3347 24294
rect 3235 24165 3268 24217
rect 3320 24165 3347 24217
rect 3235 24088 3347 24165
rect 3235 24036 3268 24088
rect 3320 24036 3347 24088
tri 3347 24084 3449 24186 sw
rect 3235 23966 3347 24036
<< via1 >>
rect 10305 35158 10357 35210
rect 10371 35158 10423 35210
rect 12199 35155 12251 35207
rect 12265 35155 12317 35207
rect 4854 35019 4906 35071
rect 4920 35019 4972 35071
rect 2910 34874 2962 34926
rect 3002 34874 3054 34926
rect 1936 34667 2052 34783
rect 1936 33240 2052 33356
rect 2105 34667 2221 34783
rect 2910 34774 2962 34826
rect 3002 34774 3054 34826
rect 2910 34674 2962 34726
rect 3002 34674 3054 34726
rect 10736 34493 10788 34545
rect 10800 34493 10852 34545
rect 11770 34493 11822 34545
rect 11834 34493 11886 34545
rect 5285 34413 5337 34465
rect 5349 34413 5401 34465
rect 2105 33240 2221 33356
rect 7725 33404 7777 33420
rect 7725 33370 7732 33404
rect 7732 33370 7766 33404
rect 7766 33370 7777 33404
rect 7725 33368 7777 33370
rect 7789 33404 7841 33420
rect 7789 33370 7808 33404
rect 7808 33370 7841 33404
rect 7789 33368 7841 33370
rect 8936 33369 8988 33421
rect 9000 33404 9052 33421
rect 9000 33370 9026 33404
rect 9026 33370 9052 33404
rect 9000 33369 9052 33370
rect 9532 33404 9584 33421
rect 9532 33370 9538 33404
rect 9538 33370 9572 33404
rect 9572 33370 9584 33404
rect 9532 33369 9584 33370
rect 9596 33404 9648 33421
rect 9596 33370 9614 33404
rect 9614 33370 9648 33404
rect 9596 33369 9648 33370
rect 16300 33404 16352 33420
rect 16300 33370 16318 33404
rect 16318 33370 16352 33404
rect 16300 33368 16352 33370
rect 16365 33368 16417 33420
rect 16429 33368 16481 33420
rect 16493 33368 16545 33420
rect 23032 32053 23084 32105
rect 23032 31989 23084 32041
rect 23032 31090 23084 31142
rect 23032 31026 23084 31078
rect 3268 30223 3320 30275
rect 3268 30095 3320 30147
rect 3268 29967 3320 30019
rect 3268 29839 3320 29891
rect 3268 29711 3320 29763
rect 3268 29583 3320 29635
rect 3268 29454 3320 29506
rect 3268 29325 3320 29377
rect 3268 29196 3320 29248
rect 3268 29067 3320 29119
rect 3268 28938 3320 28990
rect 3268 28809 3320 28861
rect 3268 28680 3320 28732
rect 3268 28551 3320 28603
rect 3268 28422 3320 28474
rect 3268 28293 3320 28345
rect 3268 28164 3320 28216
rect 3268 28035 3320 28087
rect 3268 27906 3320 27958
rect 3268 27777 3320 27829
rect 3268 27648 3320 27700
rect 3268 27519 3320 27571
rect 3268 27390 3320 27442
rect 3268 27261 3320 27313
rect 3268 27132 3320 27184
rect 3268 27003 3320 27055
rect 3268 26874 3320 26926
rect 3268 26745 3320 26797
rect 3268 26616 3320 26668
rect 3268 26487 3320 26539
rect 3268 26358 3320 26410
rect 3268 26229 3320 26281
rect 3268 26100 3320 26152
rect 3268 25971 3320 26023
rect 3268 25842 3320 25894
rect 3268 25713 3320 25765
rect 3268 25584 3320 25636
rect 3268 25455 3320 25507
rect 3268 25326 3320 25378
rect 3268 25197 3320 25249
rect 3268 25068 3320 25120
rect 3268 24939 3320 24991
rect 3268 24810 3320 24862
rect 3268 24681 3320 24733
rect 3268 24552 3320 24604
rect 3268 24423 3320 24475
rect 3960 24513 4012 24565
rect 4026 24513 4078 24565
rect 4092 24513 4144 24565
rect 4158 24513 4210 24565
rect 4224 24513 4276 24565
rect 4289 24513 4341 24565
rect 4354 24513 4406 24565
rect 4419 24513 4471 24565
rect 4484 24513 4536 24565
rect 3960 24397 4012 24449
rect 4026 24397 4078 24449
rect 4092 24397 4144 24449
rect 4158 24397 4210 24449
rect 4224 24397 4276 24449
rect 4289 24397 4341 24449
rect 4354 24397 4406 24449
rect 4419 24397 4471 24449
rect 4484 24397 4536 24449
rect 5768 24513 5820 24565
rect 5833 24513 5885 24565
rect 5898 24513 5950 24565
rect 5963 24513 6015 24565
rect 6028 24513 6080 24565
rect 6093 24513 6145 24565
rect 6158 24513 6210 24565
rect 6223 24513 6275 24565
rect 6287 24513 6339 24565
rect 5768 24397 5820 24449
rect 5833 24397 5885 24449
rect 5898 24397 5950 24449
rect 5963 24397 6015 24449
rect 6028 24397 6080 24449
rect 6093 24397 6145 24449
rect 6158 24397 6210 24449
rect 6223 24397 6275 24449
rect 6287 24397 6339 24449
rect 7247 24513 7299 24565
rect 7312 24513 7364 24565
rect 7377 24513 7429 24565
rect 7442 24513 7494 24565
rect 7507 24513 7559 24565
rect 7572 24513 7624 24565
rect 7637 24513 7689 24565
rect 7701 24513 7753 24565
rect 7765 24513 7817 24565
rect 7247 24397 7299 24449
rect 7312 24397 7364 24449
rect 7377 24397 7429 24449
rect 7442 24397 7494 24449
rect 7507 24397 7559 24449
rect 7572 24397 7624 24449
rect 7637 24397 7689 24449
rect 7701 24397 7753 24449
rect 7765 24397 7817 24449
rect 9051 24513 9103 24565
rect 9116 24513 9168 24565
rect 9181 24513 9233 24565
rect 9246 24513 9298 24565
rect 9311 24513 9363 24565
rect 9376 24513 9428 24565
rect 9441 24513 9493 24565
rect 9506 24513 9558 24565
rect 9570 24513 9622 24565
rect 9051 24397 9103 24449
rect 9116 24397 9168 24449
rect 9181 24397 9233 24449
rect 9246 24397 9298 24449
rect 9311 24397 9363 24449
rect 9376 24397 9428 24449
rect 9441 24397 9493 24449
rect 9506 24397 9558 24449
rect 9570 24397 9622 24449
rect 10855 24513 10907 24565
rect 10920 24513 10972 24565
rect 10985 24513 11037 24565
rect 11050 24513 11102 24565
rect 11115 24513 11167 24565
rect 11180 24513 11232 24565
rect 11245 24513 11297 24565
rect 11309 24513 11361 24565
rect 11373 24513 11425 24565
rect 10855 24397 10907 24449
rect 10920 24397 10972 24449
rect 10985 24397 11037 24449
rect 11050 24397 11102 24449
rect 11115 24397 11167 24449
rect 11180 24397 11232 24449
rect 11245 24397 11297 24449
rect 11309 24397 11361 24449
rect 11373 24397 11425 24449
rect 12654 24513 12706 24565
rect 12720 24513 12772 24565
rect 12786 24513 12838 24565
rect 12852 24513 12904 24565
rect 12917 24513 12969 24565
rect 12982 24513 13034 24565
rect 13047 24513 13099 24565
rect 13112 24513 13164 24565
rect 13177 24513 13229 24565
rect 12654 24397 12706 24449
rect 12720 24397 12772 24449
rect 12786 24397 12838 24449
rect 12852 24397 12904 24449
rect 12917 24397 12969 24449
rect 12982 24397 13034 24449
rect 13047 24397 13099 24449
rect 13112 24397 13164 24449
rect 13177 24397 13229 24449
rect 14463 24511 14515 24563
rect 14528 24511 14580 24563
rect 14593 24511 14645 24563
rect 14658 24511 14710 24563
rect 14723 24511 14775 24563
rect 14788 24511 14840 24563
rect 14853 24511 14905 24563
rect 14917 24511 14969 24563
rect 14981 24511 15033 24563
rect 14463 24395 14515 24447
rect 14528 24395 14580 24447
rect 14593 24395 14645 24447
rect 14658 24395 14710 24447
rect 14723 24395 14775 24447
rect 14788 24395 14840 24447
rect 14853 24395 14905 24447
rect 14917 24395 14969 24447
rect 14981 24395 15033 24447
rect 16267 24513 16319 24565
rect 16334 24513 16386 24565
rect 16401 24513 16453 24565
rect 16467 24513 16519 24565
rect 16533 24513 16585 24565
rect 16599 24513 16651 24565
rect 16665 24513 16717 24565
rect 16731 24513 16783 24565
rect 16797 24513 16849 24565
rect 16267 24397 16319 24449
rect 16334 24397 16386 24449
rect 16401 24397 16453 24449
rect 16467 24397 16519 24449
rect 16533 24397 16585 24449
rect 16599 24397 16651 24449
rect 16665 24397 16717 24449
rect 16731 24397 16783 24449
rect 16797 24397 16849 24449
rect 3268 24294 3320 24346
rect 3268 24165 3320 24217
rect 3268 24036 3320 24088
<< metal2 >>
rect 22471 36563 22527 36572
rect 22471 36483 22527 36507
tri 1930 35194 1990 35254 se
rect 1990 35210 12323 35254
rect 1990 35194 10305 35210
rect 1930 35158 10305 35194
rect 10357 35158 10371 35210
rect 10423 35207 12323 35210
rect 10423 35158 12199 35207
rect 1930 35155 12199 35158
rect 12251 35155 12265 35207
rect 12317 35155 12323 35207
rect 1930 35145 12323 35155
rect 1930 34783 2058 35145
tri 2058 35093 2110 35145 nw
tri 2149 35093 2161 35105 se
rect 2161 35093 4978 35105
rect 1930 34667 1936 34783
rect 2052 34667 2058 34783
tri 2098 35042 2149 35093 se
rect 2149 35071 4978 35093
rect 2149 35042 4854 35071
rect 2098 35019 4854 35042
rect 4906 35019 4920 35071
rect 4972 35019 4978 35071
rect 2098 34985 4978 35019
rect 2098 34783 2227 34985
tri 2227 34942 2270 34985 nw
rect 18252 34976 18308 34985
rect 2098 34667 2105 34783
rect 2221 34667 2227 34783
rect 2910 34926 3082 34932
rect 2962 34923 3002 34926
rect 3054 34923 3082 34926
rect 2968 34874 3002 34923
rect 2910 34867 2912 34874
rect 2968 34867 3026 34874
rect 2910 34828 3082 34867
rect 2910 34826 2912 34828
rect 2968 34826 3026 34828
rect 2968 34774 3002 34826
rect 10942 34794 11438 34950
tri 10942 34792 10944 34794 ne
rect 10944 34792 11438 34794
rect 12744 34794 13240 34950
rect 18252 34896 18308 34920
tri 12744 34792 12746 34794 ne
rect 12746 34792 13240 34794
rect 18126 34886 18182 34895
rect 18126 34806 18182 34830
rect 2910 34772 2912 34774
rect 2968 34772 3026 34774
rect 2910 34733 3082 34772
rect 2910 34726 2912 34733
rect 2968 34726 3026 34733
rect 2968 34677 3002 34726
rect 2962 34674 3002 34677
rect 3054 34674 3082 34677
rect 2910 34668 3082 34674
tri 18087 34545 18126 34584 se
rect 18126 34545 18182 34750
rect 10730 34493 10736 34545
rect 10788 34493 10800 34545
rect 10852 34493 11770 34545
rect 11822 34493 11834 34545
rect 11886 34524 18182 34545
rect 11886 34493 18151 34524
tri 18151 34493 18182 34524 nw
tri 18227 34703 18252 34728 se
rect 18252 34706 18308 34840
rect 18380 34976 18436 34985
rect 18380 34896 18436 34920
rect 18252 34703 18283 34706
rect 5279 34413 5285 34465
rect 5337 34413 5349 34465
rect 5401 34453 5407 34465
tri 5407 34453 5419 34465 sw
tri 18198 34453 18227 34482 se
rect 18227 34453 18283 34703
tri 18283 34681 18308 34706 nw
rect 5401 34442 18283 34453
rect 5401 34413 18254 34442
tri 18254 34413 18283 34442 nw
tri 18316 34658 18380 34722 se
rect 18380 34706 18436 34840
rect 18506 34976 18562 34985
rect 18506 34896 18562 34920
rect 18380 34658 18388 34706
tri 18388 34658 18436 34706 nw
tri 18445 34658 18506 34719 se
rect 18506 34703 18562 34840
tri 18285 34074 18316 34105 se
rect 18316 34074 18372 34658
tri 18372 34642 18388 34658 nw
rect 7719 34050 18372 34074
rect 7719 34022 18344 34050
tri 18344 34022 18372 34050 nw
tri 18405 34618 18445 34658 se
rect 18445 34647 18506 34658
tri 18506 34647 18562 34703 nw
rect 18445 34618 18461 34647
rect 1930 33240 1936 33356
rect 2052 33240 2058 33356
tri 1878 33178 1930 33230 se
rect 1930 33178 2058 33240
rect 380 33106 2058 33178
rect 380 33058 2010 33106
tri 2010 33058 2058 33106 nw
rect 2099 33240 2105 33356
rect 2221 33240 2227 33356
tri 2079 33058 2099 33078 se
rect 2099 33058 2227 33240
tri 2039 33018 2079 33058 se
rect 2079 33018 2227 33058
rect 380 32953 2227 33018
rect 380 32898 2172 32953
tri 2172 32898 2227 32953 nw
rect 3245 30275 3347 30281
rect 3245 30216 3268 30275
rect 3320 30272 3347 30275
rect 3324 30216 3347 30272
rect 3245 30171 3347 30216
rect 3245 30095 3268 30171
rect 3324 30115 3347 30171
rect 3320 30095 3347 30115
rect 3245 30070 3347 30095
rect 3245 29913 3268 30070
rect 3324 30014 3347 30070
rect 3320 29969 3347 30014
rect 3324 29913 3347 29969
rect 3245 29891 3347 29913
rect 3245 29812 3268 29891
rect 3320 29868 3347 29891
rect 3324 29812 3347 29868
rect 3245 29767 3347 29812
rect 3245 29711 3268 29767
rect 3324 29711 3347 29767
rect 3245 29666 3347 29711
rect 3245 29583 3268 29666
rect 3324 29610 3347 29666
rect 3320 29583 3347 29610
rect 3245 29565 3347 29583
rect 3245 29509 3268 29565
rect 3324 29509 3347 29565
rect 3245 29506 3347 29509
rect 3245 29408 3268 29506
rect 3320 29464 3347 29506
rect 3324 29408 3347 29464
rect 3245 29377 3347 29408
rect 3245 29307 3268 29377
rect 3320 29363 3347 29377
rect 3324 29307 3347 29363
rect 3245 29262 3347 29307
rect 3245 29196 3268 29262
rect 3324 29206 3347 29262
rect 3320 29196 3347 29206
rect 3245 29161 3347 29196
rect 3245 29067 3268 29161
rect 3324 29105 3347 29161
rect 3320 29067 3347 29105
rect 3245 29060 3347 29067
rect 3245 29004 3268 29060
rect 3324 29004 3347 29060
rect 3245 28990 3347 29004
rect 3245 28903 3268 28990
rect 3320 28959 3347 28990
rect 3324 28903 3347 28959
rect 3245 28861 3347 28903
rect 3245 28802 3268 28861
rect 3320 28858 3347 28861
rect 3324 28802 3347 28858
rect 3245 28757 3347 28802
rect 3245 28680 3268 28757
rect 3324 28701 3347 28757
rect 3320 28680 3347 28701
rect 3245 28656 3347 28680
rect 3245 28499 3268 28656
rect 3324 28600 3347 28656
rect 3320 28555 3347 28600
rect 3324 28499 3347 28555
rect 3245 28474 3347 28499
rect 3245 28398 3268 28474
rect 3320 28454 3347 28474
rect 3324 28398 3347 28454
rect 3245 28353 3347 28398
rect 3245 28293 3268 28353
rect 3324 28297 3347 28353
rect 3320 28293 3347 28297
rect 3245 28252 3347 28293
rect 3245 28164 3268 28252
rect 3324 28196 3347 28252
rect 3320 28164 3347 28196
rect 3245 28151 3347 28164
rect 3245 28095 3268 28151
rect 3324 28095 3347 28151
rect 3245 28087 3347 28095
rect 3245 27994 3268 28087
rect 3320 28050 3347 28087
rect 3324 27994 3347 28050
rect 3245 27958 3347 27994
rect 3245 27893 3268 27958
rect 3320 27949 3347 27958
rect 3324 27893 3347 27949
rect 3245 27848 3347 27893
rect 3245 27777 3268 27848
rect 3324 27792 3347 27848
rect 3320 27777 3347 27792
rect 3245 27747 3347 27777
rect 3245 27648 3268 27747
rect 3324 27691 3347 27747
rect 3320 27648 3347 27691
rect 3245 27646 3347 27648
rect 3245 27590 3268 27646
rect 3324 27590 3347 27646
rect 3245 27571 3347 27590
rect 3245 27489 3268 27571
rect 3320 27545 3347 27571
rect 3324 27489 3347 27545
rect 3245 27444 3347 27489
rect 3245 27388 3268 27444
rect 3324 27388 3347 27444
rect 3245 27343 3347 27388
rect 3245 27261 3268 27343
rect 3324 27287 3347 27343
rect 3320 27261 3347 27287
rect 3245 27242 3347 27261
rect 3245 27186 3268 27242
rect 3324 27186 3347 27242
rect 3245 27184 3347 27186
rect 3245 27085 3268 27184
rect 3320 27141 3347 27184
rect 3324 27085 3347 27141
rect 3245 27055 3347 27085
rect 3245 26984 3268 27055
rect 3320 27040 3347 27055
rect 3324 26984 3347 27040
rect 3245 26939 3347 26984
rect 3245 26874 3268 26939
rect 3324 26883 3347 26939
rect 3320 26874 3347 26883
rect 3245 26838 3347 26874
rect 3245 26745 3268 26838
rect 3324 26782 3347 26838
rect 3320 26745 3347 26782
rect 3245 26737 3347 26745
rect 3245 26681 3268 26737
rect 3324 26681 3347 26737
rect 3245 26668 3347 26681
rect 3245 26580 3268 26668
rect 3320 26636 3347 26668
rect 3324 26580 3347 26636
rect 3245 26539 3347 26580
rect 3245 26479 3268 26539
rect 3320 26535 3347 26539
rect 3324 26479 3347 26535
rect 3245 26434 3347 26479
rect 3245 26358 3268 26434
rect 3324 26378 3347 26434
rect 3320 26358 3347 26378
rect 3245 26333 3347 26358
rect 3245 26176 3268 26333
rect 3324 26277 3347 26333
rect 3320 26232 3347 26277
rect 3324 26176 3347 26232
rect 3245 26152 3347 26176
rect 3245 26075 3268 26152
rect 3320 26131 3347 26152
rect 3324 26075 3347 26131
rect 3245 26030 3347 26075
rect 3245 25971 3268 26030
rect 3324 25974 3347 26030
rect 3320 25971 3347 25974
rect 3245 25929 3347 25971
rect 3245 25842 3268 25929
rect 3324 25873 3347 25929
rect 3320 25842 3347 25873
rect 3245 25827 3347 25842
rect 3245 25771 3268 25827
rect 3324 25771 3347 25827
rect 3245 25765 3347 25771
rect 3245 25669 3268 25765
rect 3320 25725 3347 25765
rect 3324 25669 3347 25725
rect 3245 25636 3347 25669
rect 3245 25567 3268 25636
rect 3320 25623 3347 25636
rect 3324 25567 3347 25623
rect 3245 25521 3347 25567
rect 3245 25455 3268 25521
rect 3324 25465 3347 25521
rect 3320 25455 3347 25465
rect 3245 25419 3347 25455
rect 3245 25326 3268 25419
rect 3324 25363 3347 25419
rect 3320 25326 3347 25363
rect 3245 25317 3347 25326
rect 3245 25261 3268 25317
rect 3324 25261 3347 25317
rect 3245 25249 3347 25261
rect 3245 25159 3268 25249
rect 3320 25215 3347 25249
rect 3324 25159 3347 25215
rect 3245 25120 3347 25159
rect 3245 25057 3268 25120
rect 3320 25113 3347 25120
rect 3324 25057 3347 25113
rect 3245 25011 3347 25057
rect 3245 24939 3268 25011
rect 3324 24955 3347 25011
rect 3320 24939 3347 24955
rect 3245 24909 3347 24939
rect 3245 24810 3268 24909
rect 3324 24853 3347 24909
rect 3320 24810 3347 24853
rect 3245 24807 3347 24810
rect 3245 24751 3268 24807
rect 3324 24751 3347 24807
rect 3245 24733 3347 24751
rect 3245 24649 3268 24733
rect 3320 24705 3347 24733
rect 3324 24649 3347 24705
rect 3245 24604 3347 24649
rect 3245 24547 3268 24604
rect 3320 24603 3347 24604
rect 3324 24547 3347 24603
rect 3245 24501 3347 24547
rect 3245 24423 3268 24501
rect 3324 24445 3347 24501
rect 3320 24423 3347 24445
rect 3245 24399 3347 24423
rect 3245 24241 3268 24399
rect 3324 24343 3347 24399
rect 3954 24565 4542 33921
rect 3954 24513 3960 24565
rect 4019 24513 4026 24565
rect 4210 24513 4221 24565
rect 4277 24513 4289 24565
rect 4471 24513 4477 24565
rect 4536 24513 4542 24565
rect 3954 24509 3963 24513
rect 4019 24509 4049 24513
rect 4105 24509 4135 24513
rect 4191 24509 4221 24513
rect 4277 24509 4307 24513
rect 4363 24509 4392 24513
rect 4448 24509 4477 24513
rect 4533 24509 4542 24513
rect 3954 24453 4542 24509
rect 3954 24449 3963 24453
rect 4019 24449 4049 24453
rect 4105 24449 4135 24453
rect 4191 24449 4221 24453
rect 4277 24449 4307 24453
rect 4363 24449 4392 24453
rect 4448 24449 4477 24453
rect 4533 24449 4542 24453
rect 3954 24397 3960 24449
rect 4019 24397 4026 24449
rect 4210 24397 4221 24449
rect 4277 24397 4289 24449
rect 4471 24397 4477 24449
rect 4536 24397 4542 24449
rect 5762 24565 6345 33739
rect 7719 33420 7847 34022
tri 7847 33997 7872 34022 nw
tri 8930 33998 8954 34022 ne
rect 7719 33368 7725 33420
rect 7777 33368 7789 33420
rect 7841 33368 7847 33420
tri 8930 33421 8954 33445 se
rect 8954 33421 9032 34022
tri 9032 33997 9057 34022 nw
tri 9506 33978 9550 34022 ne
tri 9032 33421 9058 33447 sw
rect 8930 33369 8936 33421
rect 8988 33369 9000 33421
rect 9052 33369 9058 33421
tri 9526 33421 9550 33445 se
rect 9550 33421 9628 34022
tri 9628 33997 9653 34022 nw
rect 10806 33980 18370 33989
rect 10806 33957 18314 33980
tri 18136 33931 18162 33957 ne
rect 18162 33931 18314 33957
rect 18216 33924 18314 33931
rect 18216 33900 18370 33924
rect 18216 33844 18314 33900
rect 18216 33835 18370 33844
tri 18216 33737 18314 33835 nw
tri 9628 33421 9654 33447 sw
tri 18342 33433 18405 33496 se
rect 18405 33433 18461 34618
tri 18461 34602 18506 34647 nw
rect 9526 33369 9532 33421
rect 9584 33369 9596 33421
rect 9648 33369 9654 33421
rect 16294 33420 18461 33433
rect 7719 33355 7847 33368
rect 16294 33368 16300 33420
rect 16352 33368 16365 33420
rect 16417 33368 16429 33420
rect 16481 33368 16493 33420
rect 16545 33404 18461 33420
rect 16545 33368 18412 33404
rect 16294 33355 18412 33368
tri 18412 33355 18461 33404 nw
rect 5762 24513 5768 24565
rect 5827 24513 5833 24565
rect 6015 24513 6026 24565
rect 6082 24513 6093 24565
rect 6275 24513 6280 24565
rect 6339 24513 6345 24565
rect 5762 24509 5771 24513
rect 5827 24509 5856 24513
rect 5912 24509 5941 24513
rect 5997 24509 6026 24513
rect 6082 24509 6111 24513
rect 6167 24509 6196 24513
rect 6252 24509 6280 24513
rect 6336 24509 6345 24513
rect 5762 24453 6345 24509
rect 5762 24449 5771 24453
rect 5827 24449 5856 24453
rect 5912 24449 5941 24453
rect 5997 24449 6026 24453
rect 6082 24449 6111 24453
rect 6167 24449 6196 24453
rect 6252 24449 6280 24453
rect 6336 24449 6345 24453
rect 5762 24397 5768 24449
rect 5827 24397 5833 24449
rect 6015 24397 6026 24449
rect 6082 24397 6093 24449
rect 6275 24397 6280 24449
rect 6339 24397 6345 24449
rect 7241 24565 7823 32943
rect 7241 24513 7247 24565
rect 7306 24513 7312 24565
rect 7494 24513 7505 24565
rect 7561 24513 7572 24565
rect 7753 24513 7757 24565
rect 7817 24513 7823 24565
rect 7241 24509 7250 24513
rect 7306 24509 7335 24513
rect 7391 24509 7420 24513
rect 7476 24509 7505 24513
rect 7561 24509 7589 24513
rect 7645 24509 7673 24513
rect 7729 24509 7757 24513
rect 7813 24509 7823 24513
rect 7241 24453 7823 24509
rect 7241 24449 7250 24453
rect 7306 24449 7335 24453
rect 7391 24449 7420 24453
rect 7476 24449 7505 24453
rect 7561 24449 7589 24453
rect 7645 24449 7673 24453
rect 7729 24449 7757 24453
rect 7813 24449 7823 24453
rect 7241 24397 7247 24449
rect 7306 24397 7312 24449
rect 7494 24397 7505 24449
rect 7561 24397 7572 24449
rect 7753 24397 7757 24449
rect 7817 24397 7823 24449
rect 9045 24565 9628 32943
rect 9045 24513 9051 24565
rect 9110 24513 9116 24565
rect 9298 24513 9309 24565
rect 9365 24513 9376 24565
rect 9558 24513 9562 24565
rect 9622 24513 9628 24565
rect 9045 24509 9054 24513
rect 9110 24509 9139 24513
rect 9195 24509 9224 24513
rect 9280 24509 9309 24513
rect 9365 24509 9394 24513
rect 9450 24509 9478 24513
rect 9534 24509 9562 24513
rect 9618 24509 9628 24513
rect 9045 24453 9628 24509
rect 9045 24449 9054 24453
rect 9110 24449 9139 24453
rect 9195 24449 9224 24453
rect 9280 24449 9309 24453
rect 9365 24449 9394 24453
rect 9450 24449 9478 24453
rect 9534 24449 9562 24453
rect 9618 24449 9628 24453
rect 9045 24397 9051 24449
rect 9110 24397 9116 24449
rect 9298 24397 9309 24449
rect 9365 24397 9376 24449
rect 9558 24397 9562 24449
rect 9622 24397 9628 24449
rect 10849 24565 11431 32943
rect 10849 24513 10855 24565
rect 10914 24513 10920 24565
rect 11102 24513 11113 24565
rect 11169 24513 11180 24565
rect 11361 24513 11365 24565
rect 11425 24513 11431 24565
rect 10849 24509 10858 24513
rect 10914 24509 10943 24513
rect 10999 24509 11028 24513
rect 11084 24509 11113 24513
rect 11169 24509 11197 24513
rect 11253 24509 11281 24513
rect 11337 24509 11365 24513
rect 11421 24509 11431 24513
rect 10849 24453 11431 24509
rect 10849 24449 10858 24453
rect 10914 24449 10943 24453
rect 10999 24449 11028 24453
rect 11084 24449 11113 24453
rect 11169 24449 11197 24453
rect 11253 24449 11281 24453
rect 11337 24449 11365 24453
rect 11421 24449 11431 24453
rect 10849 24397 10855 24449
rect 10914 24397 10920 24449
rect 11102 24397 11113 24449
rect 11169 24397 11180 24449
rect 11361 24397 11365 24449
rect 11425 24397 11431 24449
rect 12648 24565 13235 32943
rect 12648 24513 12654 24565
rect 12713 24513 12720 24565
rect 12904 24513 12915 24565
rect 12971 24513 12982 24565
rect 13164 24513 13170 24565
rect 13229 24513 13235 24565
rect 12648 24509 12657 24513
rect 12713 24509 12743 24513
rect 12799 24509 12829 24513
rect 12885 24509 12915 24513
rect 12971 24509 13000 24513
rect 13056 24509 13085 24513
rect 13141 24509 13170 24513
rect 13226 24509 13235 24513
rect 12648 24453 13235 24509
rect 12648 24449 12657 24453
rect 12713 24449 12743 24453
rect 12799 24449 12829 24453
rect 12885 24449 12915 24453
rect 12971 24449 13000 24453
rect 13056 24449 13085 24453
rect 13141 24449 13170 24453
rect 13226 24449 13235 24453
rect 12648 24397 12654 24449
rect 12713 24397 12720 24449
rect 12904 24397 12915 24449
rect 12971 24397 12982 24449
rect 13164 24397 13170 24449
rect 13229 24397 13235 24449
rect 14457 24563 15039 32943
rect 14457 24511 14463 24563
rect 14522 24511 14528 24563
rect 14710 24511 14721 24563
rect 14777 24511 14788 24563
rect 14969 24511 14973 24563
rect 15033 24511 15039 24563
rect 14457 24507 14466 24511
rect 14522 24507 14551 24511
rect 14607 24507 14636 24511
rect 14692 24507 14721 24511
rect 14777 24507 14805 24511
rect 14861 24507 14889 24511
rect 14945 24507 14973 24511
rect 15029 24507 15039 24511
rect 14457 24451 15039 24507
rect 14457 24447 14466 24451
rect 14522 24447 14551 24451
rect 14607 24447 14636 24451
rect 14692 24447 14721 24451
rect 14777 24447 14805 24451
rect 14861 24447 14889 24451
rect 14945 24447 14973 24451
rect 15029 24447 15039 24451
rect 14457 24395 14463 24447
rect 14522 24395 14528 24447
rect 14710 24395 14721 24447
rect 14777 24395 14788 24447
rect 14969 24395 14973 24447
rect 15033 24395 15039 24447
rect 16261 24565 16856 32943
rect 22471 26809 22527 36427
rect 22603 36563 22659 36572
rect 22603 36483 22659 36507
tri 22571 35395 22603 35427 se
rect 22603 35395 22659 36427
rect 22571 35389 22659 35395
rect 22571 27523 22627 35389
tri 22627 35357 22659 35389 nw
rect 22731 36563 22787 36572
rect 22731 36483 22787 36507
tri 22671 35309 22731 35369 se
rect 22731 35343 22787 36427
rect 22731 35309 22745 35343
rect 22671 35301 22745 35309
tri 22745 35301 22787 35343 nw
rect 22857 36563 22913 36572
rect 22857 36483 22913 36507
tri 22831 35301 22857 35327 se
rect 22857 35301 22913 36427
rect 22671 28696 22727 35301
tri 22727 35283 22745 35301 nw
tri 22797 35267 22831 35301 se
rect 22831 35267 22853 35301
rect 22797 32111 22853 35267
tri 22853 35241 22913 35301 nw
tri 22853 32111 22893 32151 sw
rect 22797 32105 23084 32111
rect 22797 32053 23032 32105
rect 22797 32041 23084 32053
rect 22797 31989 23032 32041
rect 22797 31983 23084 31989
rect 23032 31142 23084 31148
rect 23032 31078 23084 31090
tri 22994 31011 23032 31049 se
rect 23032 31011 23084 31026
tri 22937 30954 22994 31011 se
rect 22994 30954 23027 31011
tri 23027 30954 23084 31011 nw
tri 22847 30864 22937 30954 se
tri 22937 30864 23027 30954 nw
tri 22774 30791 22847 30864 se
rect 22774 29574 22847 30791
tri 22847 30774 22937 30864 nw
tri 22774 29501 22847 29574 ne
tri 22847 29525 22931 29609 sw
rect 22847 29501 23112 29525
tri 22847 29453 22895 29501 ne
rect 22895 29453 23112 29501
tri 22727 28696 22819 28788 sw
rect 22671 28568 23032 28696
tri 22627 27523 22719 27615 sw
rect 22571 27395 22950 27523
tri 22527 26809 22619 26901 sw
rect 22471 26655 22869 26809
rect 16261 24513 16267 24565
rect 16326 24513 16334 24565
rect 16519 24513 16531 24565
rect 16587 24513 16599 24565
rect 16783 24513 16791 24565
rect 16849 24513 16856 24565
rect 16261 24509 16270 24513
rect 16326 24509 16357 24513
rect 16413 24509 16444 24513
rect 16500 24509 16531 24513
rect 16587 24509 16618 24513
rect 16674 24509 16705 24513
rect 16761 24509 16791 24513
rect 16847 24509 16856 24513
rect 16261 24453 16856 24509
rect 16261 24449 16270 24453
rect 16326 24449 16357 24453
rect 16413 24449 16444 24453
rect 16500 24449 16531 24453
rect 16587 24449 16618 24453
rect 16674 24449 16705 24453
rect 16761 24449 16791 24453
rect 16847 24449 16856 24453
rect 16261 24397 16267 24449
rect 16326 24397 16334 24449
rect 16519 24397 16531 24449
rect 16587 24397 16599 24449
rect 16783 24397 16791 24449
rect 16849 24397 16856 24449
rect 3320 24297 3347 24343
rect 3324 24241 3347 24297
rect 3245 24217 3347 24241
rect 3245 24139 3268 24217
rect 3320 24195 3347 24217
rect 3324 24139 3347 24195
rect 3245 24093 3347 24139
rect 3245 24036 3268 24093
rect 3324 24037 3347 24093
rect 3320 24036 3347 24037
rect 3245 24028 3347 24036
<< via2 >>
rect 22471 36507 22527 36563
rect 22471 36427 22527 36483
rect 2912 34874 2962 34923
rect 2962 34874 2968 34923
rect 3026 34874 3054 34923
rect 3054 34874 3082 34923
rect 2912 34867 2968 34874
rect 3026 34867 3082 34874
rect 2912 34826 2968 34828
rect 3026 34826 3082 34828
rect 2912 34774 2962 34826
rect 2962 34774 2968 34826
rect 3026 34774 3054 34826
rect 3054 34774 3082 34826
rect 18252 34920 18308 34976
rect 18126 34830 18182 34886
rect 2912 34772 2968 34774
rect 3026 34772 3082 34774
rect 2912 34726 2968 34733
rect 3026 34726 3082 34733
rect 2912 34677 2962 34726
rect 2962 34677 2968 34726
rect 3026 34677 3054 34726
rect 3054 34677 3082 34726
rect 18126 34750 18182 34806
rect 18252 34840 18308 34896
rect 18380 34920 18436 34976
rect 18380 34840 18436 34896
rect 18506 34920 18562 34976
rect 18506 34840 18562 34896
rect 3268 30223 3320 30272
rect 3320 30223 3324 30272
rect 3268 30216 3324 30223
rect 3268 30147 3324 30171
rect 3268 30115 3320 30147
rect 3320 30115 3324 30147
rect 3268 30019 3324 30070
rect 3268 30014 3320 30019
rect 3320 30014 3324 30019
rect 3268 29967 3320 29969
rect 3320 29967 3324 29969
rect 3268 29913 3324 29967
rect 3268 29839 3320 29868
rect 3320 29839 3324 29868
rect 3268 29812 3324 29839
rect 3268 29763 3324 29767
rect 3268 29711 3320 29763
rect 3320 29711 3324 29763
rect 3268 29635 3324 29666
rect 3268 29610 3320 29635
rect 3320 29610 3324 29635
rect 3268 29509 3324 29565
rect 3268 29454 3320 29464
rect 3320 29454 3324 29464
rect 3268 29408 3324 29454
rect 3268 29325 3320 29363
rect 3320 29325 3324 29363
rect 3268 29307 3324 29325
rect 3268 29248 3324 29262
rect 3268 29206 3320 29248
rect 3320 29206 3324 29248
rect 3268 29119 3324 29161
rect 3268 29105 3320 29119
rect 3320 29105 3324 29119
rect 3268 29004 3324 29060
rect 3268 28938 3320 28959
rect 3320 28938 3324 28959
rect 3268 28903 3324 28938
rect 3268 28809 3320 28858
rect 3320 28809 3324 28858
rect 3268 28802 3324 28809
rect 3268 28732 3324 28757
rect 3268 28701 3320 28732
rect 3320 28701 3324 28732
rect 3268 28603 3324 28656
rect 3268 28600 3320 28603
rect 3320 28600 3324 28603
rect 3268 28551 3320 28555
rect 3320 28551 3324 28555
rect 3268 28499 3324 28551
rect 3268 28422 3320 28454
rect 3320 28422 3324 28454
rect 3268 28398 3324 28422
rect 3268 28345 3324 28353
rect 3268 28297 3320 28345
rect 3320 28297 3324 28345
rect 3268 28216 3324 28252
rect 3268 28196 3320 28216
rect 3320 28196 3324 28216
rect 3268 28095 3324 28151
rect 3268 28035 3320 28050
rect 3320 28035 3324 28050
rect 3268 27994 3324 28035
rect 3268 27906 3320 27949
rect 3320 27906 3324 27949
rect 3268 27893 3324 27906
rect 3268 27829 3324 27848
rect 3268 27792 3320 27829
rect 3320 27792 3324 27829
rect 3268 27700 3324 27747
rect 3268 27691 3320 27700
rect 3320 27691 3324 27700
rect 3268 27590 3324 27646
rect 3268 27519 3320 27545
rect 3320 27519 3324 27545
rect 3268 27489 3324 27519
rect 3268 27442 3324 27444
rect 3268 27390 3320 27442
rect 3320 27390 3324 27442
rect 3268 27388 3324 27390
rect 3268 27313 3324 27343
rect 3268 27287 3320 27313
rect 3320 27287 3324 27313
rect 3268 27186 3324 27242
rect 3268 27132 3320 27141
rect 3320 27132 3324 27141
rect 3268 27085 3324 27132
rect 3268 27003 3320 27040
rect 3320 27003 3324 27040
rect 3268 26984 3324 27003
rect 3268 26926 3324 26939
rect 3268 26883 3320 26926
rect 3320 26883 3324 26926
rect 3268 26797 3324 26838
rect 3268 26782 3320 26797
rect 3320 26782 3324 26797
rect 3268 26681 3324 26737
rect 3268 26616 3320 26636
rect 3320 26616 3324 26636
rect 3268 26580 3324 26616
rect 3268 26487 3320 26535
rect 3320 26487 3324 26535
rect 3268 26479 3324 26487
rect 3268 26410 3324 26434
rect 3268 26378 3320 26410
rect 3320 26378 3324 26410
rect 3268 26281 3324 26333
rect 3268 26277 3320 26281
rect 3320 26277 3324 26281
rect 3268 26229 3320 26232
rect 3320 26229 3324 26232
rect 3268 26176 3324 26229
rect 3268 26100 3320 26131
rect 3320 26100 3324 26131
rect 3268 26075 3324 26100
rect 3268 26023 3324 26030
rect 3268 25974 3320 26023
rect 3320 25974 3324 26023
rect 3268 25894 3324 25929
rect 3268 25873 3320 25894
rect 3320 25873 3324 25894
rect 3268 25771 3324 25827
rect 3268 25713 3320 25725
rect 3320 25713 3324 25725
rect 3268 25669 3324 25713
rect 3268 25584 3320 25623
rect 3320 25584 3324 25623
rect 3268 25567 3324 25584
rect 3268 25507 3324 25521
rect 3268 25465 3320 25507
rect 3320 25465 3324 25507
rect 3268 25378 3324 25419
rect 3268 25363 3320 25378
rect 3320 25363 3324 25378
rect 3268 25261 3324 25317
rect 3268 25197 3320 25215
rect 3320 25197 3324 25215
rect 3268 25159 3324 25197
rect 3268 25068 3320 25113
rect 3320 25068 3324 25113
rect 3268 25057 3324 25068
rect 3268 24991 3324 25011
rect 3268 24955 3320 24991
rect 3320 24955 3324 24991
rect 3268 24862 3324 24909
rect 3268 24853 3320 24862
rect 3320 24853 3324 24862
rect 3268 24751 3324 24807
rect 3268 24681 3320 24705
rect 3320 24681 3324 24705
rect 3268 24649 3324 24681
rect 3268 24552 3320 24603
rect 3320 24552 3324 24603
rect 3268 24547 3324 24552
rect 3268 24475 3324 24501
rect 3268 24445 3320 24475
rect 3320 24445 3324 24475
rect 3268 24346 3324 24399
rect 3268 24343 3320 24346
rect 3320 24343 3324 24346
rect 3963 24513 4012 24565
rect 4012 24513 4019 24565
rect 4049 24513 4078 24565
rect 4078 24513 4092 24565
rect 4092 24513 4105 24565
rect 4135 24513 4144 24565
rect 4144 24513 4158 24565
rect 4158 24513 4191 24565
rect 4221 24513 4224 24565
rect 4224 24513 4276 24565
rect 4276 24513 4277 24565
rect 4307 24513 4341 24565
rect 4341 24513 4354 24565
rect 4354 24513 4363 24565
rect 4392 24513 4406 24565
rect 4406 24513 4419 24565
rect 4419 24513 4448 24565
rect 4477 24513 4484 24565
rect 4484 24513 4533 24565
rect 3963 24509 4019 24513
rect 4049 24509 4105 24513
rect 4135 24509 4191 24513
rect 4221 24509 4277 24513
rect 4307 24509 4363 24513
rect 4392 24509 4448 24513
rect 4477 24509 4533 24513
rect 3963 24449 4019 24453
rect 4049 24449 4105 24453
rect 4135 24449 4191 24453
rect 4221 24449 4277 24453
rect 4307 24449 4363 24453
rect 4392 24449 4448 24453
rect 4477 24449 4533 24453
rect 3963 24397 4012 24449
rect 4012 24397 4019 24449
rect 4049 24397 4078 24449
rect 4078 24397 4092 24449
rect 4092 24397 4105 24449
rect 4135 24397 4144 24449
rect 4144 24397 4158 24449
rect 4158 24397 4191 24449
rect 4221 24397 4224 24449
rect 4224 24397 4276 24449
rect 4276 24397 4277 24449
rect 4307 24397 4341 24449
rect 4341 24397 4354 24449
rect 4354 24397 4363 24449
rect 4392 24397 4406 24449
rect 4406 24397 4419 24449
rect 4419 24397 4448 24449
rect 4477 24397 4484 24449
rect 4484 24397 4533 24449
rect 18314 33924 18370 33980
rect 18314 33844 18370 33900
rect 5771 24513 5820 24565
rect 5820 24513 5827 24565
rect 5856 24513 5885 24565
rect 5885 24513 5898 24565
rect 5898 24513 5912 24565
rect 5941 24513 5950 24565
rect 5950 24513 5963 24565
rect 5963 24513 5997 24565
rect 6026 24513 6028 24565
rect 6028 24513 6080 24565
rect 6080 24513 6082 24565
rect 6111 24513 6145 24565
rect 6145 24513 6158 24565
rect 6158 24513 6167 24565
rect 6196 24513 6210 24565
rect 6210 24513 6223 24565
rect 6223 24513 6252 24565
rect 6280 24513 6287 24565
rect 6287 24513 6336 24565
rect 5771 24509 5827 24513
rect 5856 24509 5912 24513
rect 5941 24509 5997 24513
rect 6026 24509 6082 24513
rect 6111 24509 6167 24513
rect 6196 24509 6252 24513
rect 6280 24509 6336 24513
rect 5771 24449 5827 24453
rect 5856 24449 5912 24453
rect 5941 24449 5997 24453
rect 6026 24449 6082 24453
rect 6111 24449 6167 24453
rect 6196 24449 6252 24453
rect 6280 24449 6336 24453
rect 5771 24397 5820 24449
rect 5820 24397 5827 24449
rect 5856 24397 5885 24449
rect 5885 24397 5898 24449
rect 5898 24397 5912 24449
rect 5941 24397 5950 24449
rect 5950 24397 5963 24449
rect 5963 24397 5997 24449
rect 6026 24397 6028 24449
rect 6028 24397 6080 24449
rect 6080 24397 6082 24449
rect 6111 24397 6145 24449
rect 6145 24397 6158 24449
rect 6158 24397 6167 24449
rect 6196 24397 6210 24449
rect 6210 24397 6223 24449
rect 6223 24397 6252 24449
rect 6280 24397 6287 24449
rect 6287 24397 6336 24449
rect 7250 24513 7299 24565
rect 7299 24513 7306 24565
rect 7335 24513 7364 24565
rect 7364 24513 7377 24565
rect 7377 24513 7391 24565
rect 7420 24513 7429 24565
rect 7429 24513 7442 24565
rect 7442 24513 7476 24565
rect 7505 24513 7507 24565
rect 7507 24513 7559 24565
rect 7559 24513 7561 24565
rect 7589 24513 7624 24565
rect 7624 24513 7637 24565
rect 7637 24513 7645 24565
rect 7673 24513 7689 24565
rect 7689 24513 7701 24565
rect 7701 24513 7729 24565
rect 7757 24513 7765 24565
rect 7765 24513 7813 24565
rect 7250 24509 7306 24513
rect 7335 24509 7391 24513
rect 7420 24509 7476 24513
rect 7505 24509 7561 24513
rect 7589 24509 7645 24513
rect 7673 24509 7729 24513
rect 7757 24509 7813 24513
rect 7250 24449 7306 24453
rect 7335 24449 7391 24453
rect 7420 24449 7476 24453
rect 7505 24449 7561 24453
rect 7589 24449 7645 24453
rect 7673 24449 7729 24453
rect 7757 24449 7813 24453
rect 7250 24397 7299 24449
rect 7299 24397 7306 24449
rect 7335 24397 7364 24449
rect 7364 24397 7377 24449
rect 7377 24397 7391 24449
rect 7420 24397 7429 24449
rect 7429 24397 7442 24449
rect 7442 24397 7476 24449
rect 7505 24397 7507 24449
rect 7507 24397 7559 24449
rect 7559 24397 7561 24449
rect 7589 24397 7624 24449
rect 7624 24397 7637 24449
rect 7637 24397 7645 24449
rect 7673 24397 7689 24449
rect 7689 24397 7701 24449
rect 7701 24397 7729 24449
rect 7757 24397 7765 24449
rect 7765 24397 7813 24449
rect 9054 24513 9103 24565
rect 9103 24513 9110 24565
rect 9139 24513 9168 24565
rect 9168 24513 9181 24565
rect 9181 24513 9195 24565
rect 9224 24513 9233 24565
rect 9233 24513 9246 24565
rect 9246 24513 9280 24565
rect 9309 24513 9311 24565
rect 9311 24513 9363 24565
rect 9363 24513 9365 24565
rect 9394 24513 9428 24565
rect 9428 24513 9441 24565
rect 9441 24513 9450 24565
rect 9478 24513 9493 24565
rect 9493 24513 9506 24565
rect 9506 24513 9534 24565
rect 9562 24513 9570 24565
rect 9570 24513 9618 24565
rect 9054 24509 9110 24513
rect 9139 24509 9195 24513
rect 9224 24509 9280 24513
rect 9309 24509 9365 24513
rect 9394 24509 9450 24513
rect 9478 24509 9534 24513
rect 9562 24509 9618 24513
rect 9054 24449 9110 24453
rect 9139 24449 9195 24453
rect 9224 24449 9280 24453
rect 9309 24449 9365 24453
rect 9394 24449 9450 24453
rect 9478 24449 9534 24453
rect 9562 24449 9618 24453
rect 9054 24397 9103 24449
rect 9103 24397 9110 24449
rect 9139 24397 9168 24449
rect 9168 24397 9181 24449
rect 9181 24397 9195 24449
rect 9224 24397 9233 24449
rect 9233 24397 9246 24449
rect 9246 24397 9280 24449
rect 9309 24397 9311 24449
rect 9311 24397 9363 24449
rect 9363 24397 9365 24449
rect 9394 24397 9428 24449
rect 9428 24397 9441 24449
rect 9441 24397 9450 24449
rect 9478 24397 9493 24449
rect 9493 24397 9506 24449
rect 9506 24397 9534 24449
rect 9562 24397 9570 24449
rect 9570 24397 9618 24449
rect 10858 24513 10907 24565
rect 10907 24513 10914 24565
rect 10943 24513 10972 24565
rect 10972 24513 10985 24565
rect 10985 24513 10999 24565
rect 11028 24513 11037 24565
rect 11037 24513 11050 24565
rect 11050 24513 11084 24565
rect 11113 24513 11115 24565
rect 11115 24513 11167 24565
rect 11167 24513 11169 24565
rect 11197 24513 11232 24565
rect 11232 24513 11245 24565
rect 11245 24513 11253 24565
rect 11281 24513 11297 24565
rect 11297 24513 11309 24565
rect 11309 24513 11337 24565
rect 11365 24513 11373 24565
rect 11373 24513 11421 24565
rect 10858 24509 10914 24513
rect 10943 24509 10999 24513
rect 11028 24509 11084 24513
rect 11113 24509 11169 24513
rect 11197 24509 11253 24513
rect 11281 24509 11337 24513
rect 11365 24509 11421 24513
rect 10858 24449 10914 24453
rect 10943 24449 10999 24453
rect 11028 24449 11084 24453
rect 11113 24449 11169 24453
rect 11197 24449 11253 24453
rect 11281 24449 11337 24453
rect 11365 24449 11421 24453
rect 10858 24397 10907 24449
rect 10907 24397 10914 24449
rect 10943 24397 10972 24449
rect 10972 24397 10985 24449
rect 10985 24397 10999 24449
rect 11028 24397 11037 24449
rect 11037 24397 11050 24449
rect 11050 24397 11084 24449
rect 11113 24397 11115 24449
rect 11115 24397 11167 24449
rect 11167 24397 11169 24449
rect 11197 24397 11232 24449
rect 11232 24397 11245 24449
rect 11245 24397 11253 24449
rect 11281 24397 11297 24449
rect 11297 24397 11309 24449
rect 11309 24397 11337 24449
rect 11365 24397 11373 24449
rect 11373 24397 11421 24449
rect 12657 24513 12706 24565
rect 12706 24513 12713 24565
rect 12743 24513 12772 24565
rect 12772 24513 12786 24565
rect 12786 24513 12799 24565
rect 12829 24513 12838 24565
rect 12838 24513 12852 24565
rect 12852 24513 12885 24565
rect 12915 24513 12917 24565
rect 12917 24513 12969 24565
rect 12969 24513 12971 24565
rect 13000 24513 13034 24565
rect 13034 24513 13047 24565
rect 13047 24513 13056 24565
rect 13085 24513 13099 24565
rect 13099 24513 13112 24565
rect 13112 24513 13141 24565
rect 13170 24513 13177 24565
rect 13177 24513 13226 24565
rect 12657 24509 12713 24513
rect 12743 24509 12799 24513
rect 12829 24509 12885 24513
rect 12915 24509 12971 24513
rect 13000 24509 13056 24513
rect 13085 24509 13141 24513
rect 13170 24509 13226 24513
rect 12657 24449 12713 24453
rect 12743 24449 12799 24453
rect 12829 24449 12885 24453
rect 12915 24449 12971 24453
rect 13000 24449 13056 24453
rect 13085 24449 13141 24453
rect 13170 24449 13226 24453
rect 12657 24397 12706 24449
rect 12706 24397 12713 24449
rect 12743 24397 12772 24449
rect 12772 24397 12786 24449
rect 12786 24397 12799 24449
rect 12829 24397 12838 24449
rect 12838 24397 12852 24449
rect 12852 24397 12885 24449
rect 12915 24397 12917 24449
rect 12917 24397 12969 24449
rect 12969 24397 12971 24449
rect 13000 24397 13034 24449
rect 13034 24397 13047 24449
rect 13047 24397 13056 24449
rect 13085 24397 13099 24449
rect 13099 24397 13112 24449
rect 13112 24397 13141 24449
rect 13170 24397 13177 24449
rect 13177 24397 13226 24449
rect 14466 24511 14515 24563
rect 14515 24511 14522 24563
rect 14551 24511 14580 24563
rect 14580 24511 14593 24563
rect 14593 24511 14607 24563
rect 14636 24511 14645 24563
rect 14645 24511 14658 24563
rect 14658 24511 14692 24563
rect 14721 24511 14723 24563
rect 14723 24511 14775 24563
rect 14775 24511 14777 24563
rect 14805 24511 14840 24563
rect 14840 24511 14853 24563
rect 14853 24511 14861 24563
rect 14889 24511 14905 24563
rect 14905 24511 14917 24563
rect 14917 24511 14945 24563
rect 14973 24511 14981 24563
rect 14981 24511 15029 24563
rect 14466 24507 14522 24511
rect 14551 24507 14607 24511
rect 14636 24507 14692 24511
rect 14721 24507 14777 24511
rect 14805 24507 14861 24511
rect 14889 24507 14945 24511
rect 14973 24507 15029 24511
rect 14466 24447 14522 24451
rect 14551 24447 14607 24451
rect 14636 24447 14692 24451
rect 14721 24447 14777 24451
rect 14805 24447 14861 24451
rect 14889 24447 14945 24451
rect 14973 24447 15029 24451
rect 14466 24395 14515 24447
rect 14515 24395 14522 24447
rect 14551 24395 14580 24447
rect 14580 24395 14593 24447
rect 14593 24395 14607 24447
rect 14636 24395 14645 24447
rect 14645 24395 14658 24447
rect 14658 24395 14692 24447
rect 14721 24395 14723 24447
rect 14723 24395 14775 24447
rect 14775 24395 14777 24447
rect 14805 24395 14840 24447
rect 14840 24395 14853 24447
rect 14853 24395 14861 24447
rect 14889 24395 14905 24447
rect 14905 24395 14917 24447
rect 14917 24395 14945 24447
rect 14973 24395 14981 24447
rect 14981 24395 15029 24447
rect 22603 36507 22659 36563
rect 22603 36427 22659 36483
rect 22731 36507 22787 36563
rect 22731 36427 22787 36483
rect 22857 36507 22913 36563
rect 22857 36427 22913 36483
rect 16270 24513 16319 24565
rect 16319 24513 16326 24565
rect 16357 24513 16386 24565
rect 16386 24513 16401 24565
rect 16401 24513 16413 24565
rect 16444 24513 16453 24565
rect 16453 24513 16467 24565
rect 16467 24513 16500 24565
rect 16531 24513 16533 24565
rect 16533 24513 16585 24565
rect 16585 24513 16587 24565
rect 16618 24513 16651 24565
rect 16651 24513 16665 24565
rect 16665 24513 16674 24565
rect 16705 24513 16717 24565
rect 16717 24513 16731 24565
rect 16731 24513 16761 24565
rect 16791 24513 16797 24565
rect 16797 24513 16847 24565
rect 16270 24509 16326 24513
rect 16357 24509 16413 24513
rect 16444 24509 16500 24513
rect 16531 24509 16587 24513
rect 16618 24509 16674 24513
rect 16705 24509 16761 24513
rect 16791 24509 16847 24513
rect 16270 24449 16326 24453
rect 16357 24449 16413 24453
rect 16444 24449 16500 24453
rect 16531 24449 16587 24453
rect 16618 24449 16674 24453
rect 16705 24449 16761 24453
rect 16791 24449 16847 24453
rect 16270 24397 16319 24449
rect 16319 24397 16326 24449
rect 16357 24397 16386 24449
rect 16386 24397 16401 24449
rect 16401 24397 16413 24449
rect 16444 24397 16453 24449
rect 16453 24397 16467 24449
rect 16467 24397 16500 24449
rect 16531 24397 16533 24449
rect 16533 24397 16585 24449
rect 16585 24397 16587 24449
rect 16618 24397 16651 24449
rect 16651 24397 16665 24449
rect 16665 24397 16674 24449
rect 16705 24397 16717 24449
rect 16717 24397 16731 24449
rect 16731 24397 16761 24449
rect 16791 24397 16797 24449
rect 16797 24397 16847 24449
rect 3268 24294 3320 24297
rect 3320 24294 3324 24297
rect 3268 24241 3324 24294
rect 3268 24165 3320 24195
rect 3320 24165 3324 24195
rect 3268 24139 3324 24165
rect 3268 24088 3324 24093
rect 3268 24037 3320 24088
rect 3320 24037 3324 24088
<< metal3 >>
tri 18121 36947 18222 37048 se
rect 18222 36978 22817 37048
rect 18222 36947 18248 36978
tri 18248 36947 18279 36978 nw
tri 14612 36745 14769 36902 ne
rect 2907 34923 3087 34928
rect 2907 34867 2912 34923
rect 2968 34867 3026 34923
rect 3082 34867 3087 34923
rect 2907 34828 3087 34867
rect 2907 34772 2912 34828
rect 2968 34772 3026 34828
rect 3082 34772 3087 34828
rect 2907 34733 3087 34772
rect 18121 34886 18187 36947
tri 18187 36886 18248 36947 nw
tri 22760 36921 22817 36978 ne
tri 22817 36947 22918 37048 sw
rect 22817 36921 22918 36947
tri 18317 36886 18348 36917 se
rect 18348 36886 22691 36917
rect 18121 34830 18126 34886
rect 18182 34830 18187 34886
tri 18247 36816 18317 36886 se
rect 18317 36847 22691 36886
rect 18317 36816 18344 36847
rect 18247 36786 18344 36816
tri 18344 36786 18405 36847 nw
tri 22634 36790 22691 36847 ne
tri 22691 36816 22792 36917 sw
tri 22817 36886 22852 36921 ne
rect 22691 36790 22792 36816
rect 18247 34976 18313 36786
tri 18313 36755 18344 36786 nw
rect 18247 34920 18252 34976
rect 18308 34920 18313 34976
rect 18247 34896 18313 34920
rect 18247 34840 18252 34896
rect 18308 34840 18313 34896
rect 18247 34835 18313 34840
tri 18375 36685 18476 36786 se
rect 18476 36716 22563 36786
rect 18476 36685 18502 36716
tri 18502 36685 18533 36716 nw
rect 18375 34976 18441 36685
tri 18441 36624 18502 36685 nw
tri 22506 36659 22563 36716 ne
tri 22563 36685 22664 36786 sw
tri 22691 36755 22726 36790 ne
rect 22563 36659 22664 36685
tri 18514 36554 18615 36655 se
rect 18615 36585 22431 36655
rect 18615 36554 18628 36585
rect 18375 34920 18380 34976
rect 18436 34920 18441 34976
rect 18375 34896 18441 34920
rect 18375 34840 18380 34896
rect 18436 34840 18441 34896
rect 18375 34835 18441 34840
tri 18501 36541 18514 36554 se
rect 18514 36541 18628 36554
tri 18628 36541 18672 36585 nw
rect 18501 34976 18567 36541
tri 18567 36480 18628 36541 nw
tri 22374 36528 22431 36585 ne
tri 22431 36568 22518 36655 sw
tri 22563 36624 22598 36659 ne
rect 22431 36563 22532 36568
rect 22431 36528 22471 36563
rect 18501 34920 18506 34976
rect 18562 34920 18567 34976
rect 18501 34896 18567 34920
rect 18501 34840 18506 34896
rect 18562 34840 18567 34896
rect 18501 34835 18567 34840
tri 18629 36416 18733 36520 se
rect 18733 36493 22263 36520
tri 22263 36493 22290 36520 sw
tri 22431 36493 22466 36528 ne
rect 22466 36507 22471 36528
rect 22527 36507 22532 36563
rect 18733 36416 22290 36493
rect 18629 36400 22290 36416
rect 18121 34806 18187 34830
rect 18121 34750 18126 34806
rect 18182 34750 18187 34806
rect 18121 34745 18187 34750
rect 2907 34677 2912 34733
rect 2968 34677 3026 34733
rect 3082 34677 3087 34733
rect 2907 34672 3087 34677
rect 3240 30272 3352 30277
rect 3240 30216 3268 30272
rect 3324 30216 3352 30272
rect 3240 30171 3352 30216
rect 3240 30115 3268 30171
rect 3324 30115 3352 30171
rect 3240 30070 3352 30115
rect 3240 30014 3268 30070
rect 3324 30014 3352 30070
rect 3240 29969 3352 30014
rect 3240 29913 3268 29969
rect 3324 29913 3352 29969
rect 3240 29868 3352 29913
rect 3240 29812 3268 29868
rect 3324 29812 3352 29868
rect 3240 29767 3352 29812
rect 3240 29711 3268 29767
rect 3324 29711 3352 29767
rect 3240 29666 3352 29711
rect 3240 29610 3268 29666
rect 3324 29610 3352 29666
rect 3240 29565 3352 29610
rect 3240 29509 3268 29565
rect 3324 29509 3352 29565
rect 3240 29464 3352 29509
rect 3240 29408 3268 29464
rect 3324 29408 3352 29464
rect 3240 29363 3352 29408
rect 3240 29307 3268 29363
rect 3324 29307 3352 29363
rect 3240 29262 3352 29307
rect 3240 29206 3268 29262
rect 3324 29206 3352 29262
rect 3240 29161 3352 29206
rect 3240 29105 3268 29161
rect 3324 29105 3352 29161
rect 3240 29060 3352 29105
rect 3240 29004 3268 29060
rect 3324 29004 3352 29060
rect 3240 28959 3352 29004
rect 3240 28903 3268 28959
rect 3324 28903 3352 28959
rect 3240 28858 3352 28903
rect 3240 28802 3268 28858
rect 3324 28802 3352 28858
rect 3240 28757 3352 28802
rect 3240 28701 3268 28757
rect 3324 28701 3352 28757
rect 3240 28656 3352 28701
rect 3240 28600 3268 28656
rect 3324 28600 3352 28656
rect 3240 28555 3352 28600
rect 3240 28499 3268 28555
rect 3324 28499 3352 28555
rect 3240 28454 3352 28499
rect 3240 28398 3268 28454
rect 3324 28398 3352 28454
rect 3240 28353 3352 28398
rect 3240 28297 3268 28353
rect 3324 28297 3352 28353
rect 3240 28252 3352 28297
rect 3240 28196 3268 28252
rect 3324 28196 3352 28252
rect 3240 28151 3352 28196
rect 3240 28095 3268 28151
rect 3324 28095 3352 28151
rect 3240 28050 3352 28095
rect 3240 27994 3268 28050
rect 3324 27994 3352 28050
rect 3240 27949 3352 27994
rect 3240 27893 3268 27949
rect 3324 27893 3352 27949
rect 3240 27848 3352 27893
rect 3240 27792 3268 27848
rect 3324 27792 3352 27848
rect 3240 27747 3352 27792
rect 3240 27691 3268 27747
rect 3324 27691 3352 27747
rect 3240 27646 3352 27691
rect 3240 27590 3268 27646
rect 3324 27590 3352 27646
rect 3240 27545 3352 27590
rect 3240 27489 3268 27545
rect 3324 27489 3352 27545
rect 3240 27444 3352 27489
rect 3240 27388 3268 27444
rect 3324 27388 3352 27444
rect 3240 27343 3352 27388
rect 3240 27287 3268 27343
rect 3324 27287 3352 27343
rect 3240 27242 3352 27287
rect 3240 27186 3268 27242
rect 3324 27186 3352 27242
rect 3240 27141 3352 27186
rect 3240 27085 3268 27141
rect 3324 27085 3352 27141
rect 3240 27040 3352 27085
rect 3240 26984 3268 27040
rect 3324 26984 3352 27040
rect 3240 26939 3352 26984
rect 3240 26883 3268 26939
rect 3324 26883 3352 26939
rect 3240 26838 3352 26883
rect 3240 26782 3268 26838
rect 3324 26782 3352 26838
rect 3240 26737 3352 26782
rect 3240 26681 3268 26737
rect 3324 26681 3352 26737
rect 3240 26636 3352 26681
rect 3240 26580 3268 26636
rect 3324 26580 3352 26636
rect 3240 26535 3352 26580
rect 3240 26479 3268 26535
rect 3324 26479 3352 26535
rect 3240 26434 3352 26479
rect 3240 26378 3268 26434
rect 3324 26378 3352 26434
rect 3240 26333 3352 26378
rect 3240 26277 3268 26333
rect 3324 26277 3352 26333
rect 3240 26232 3352 26277
rect 3240 26176 3268 26232
rect 3324 26176 3352 26232
rect 3240 26131 3352 26176
rect 3240 26075 3268 26131
rect 3324 26075 3352 26131
rect 3240 26030 3352 26075
rect 3240 25974 3268 26030
rect 3324 25974 3352 26030
rect 3240 25929 3352 25974
rect 3240 25873 3268 25929
rect 3324 25873 3352 25929
rect 3240 25827 3352 25873
rect 3240 25771 3268 25827
rect 3324 25771 3352 25827
rect 3240 25725 3352 25771
rect 3240 25669 3268 25725
rect 3324 25669 3352 25725
rect 3240 25623 3352 25669
rect 3240 25567 3268 25623
rect 3324 25567 3352 25623
rect 3240 25521 3352 25567
rect 3240 25465 3268 25521
rect 3324 25465 3352 25521
rect 3240 25419 3352 25465
rect 3240 25363 3268 25419
rect 3324 25363 3352 25419
rect 3240 25317 3352 25363
rect 3240 25261 3268 25317
rect 3324 25261 3352 25317
rect 3240 25215 3352 25261
rect 3240 25159 3268 25215
rect 3324 25159 3352 25215
rect 3240 25113 3352 25159
rect 3240 25057 3268 25113
rect 3324 25057 3352 25113
rect 3240 25011 3352 25057
rect 3240 24955 3268 25011
rect 3324 24955 3352 25011
rect 3240 24909 3352 24955
rect 3240 24853 3268 24909
rect 3324 24853 3352 24909
rect 3240 24807 3352 24853
rect 3240 24751 3268 24807
rect 3324 24751 3352 24807
rect 3240 24705 3352 24751
rect 3240 24649 3268 24705
rect 3324 24649 3352 24705
rect 3240 24603 3352 24649
rect 3240 24547 3268 24603
rect 3324 24547 3352 24603
rect 3240 24501 3352 24547
rect 3240 24445 3268 24501
rect 3324 24445 3352 24501
rect 3240 24399 3352 24445
rect 3240 24343 3268 24399
rect 3324 24343 3352 24399
rect 3949 24565 4541 33890
rect 3949 24509 3963 24565
rect 4019 24509 4049 24565
rect 4105 24509 4135 24565
rect 4191 24509 4221 24565
rect 4277 24509 4307 24565
rect 4363 24509 4392 24565
rect 4448 24509 4477 24565
rect 4533 24509 4541 24565
rect 3949 24453 4541 24509
rect 3949 24397 3963 24453
rect 4019 24397 4049 24453
rect 4105 24397 4135 24453
rect 4191 24397 4221 24453
rect 4277 24397 4307 24453
rect 4363 24397 4392 24453
rect 4448 24397 4477 24453
rect 4533 24397 4541 24453
rect 3949 24367 4541 24397
rect 3240 24297 3352 24343
rect 3240 24241 3268 24297
rect 3324 24241 3352 24297
rect 3240 24195 3352 24241
rect 3240 24139 3268 24195
rect 3324 24139 3352 24195
rect 3240 24093 3352 24139
rect 3240 24037 3268 24093
rect 3324 24037 3352 24093
rect 3240 24032 3352 24037
rect 4853 21949 5445 33634
rect 5758 24946 6352 33921
rect 5758 24565 6347 24946
tri 6347 24941 6352 24946 nw
rect 5758 24509 5771 24565
rect 5827 24509 5856 24565
rect 5912 24509 5941 24565
rect 5997 24509 6026 24565
rect 6082 24509 6111 24565
rect 6167 24509 6196 24565
rect 6252 24509 6280 24565
rect 6336 24509 6347 24565
rect 5758 24453 6347 24509
rect 5758 24397 5771 24453
rect 5827 24397 5856 24453
rect 5912 24397 5941 24453
rect 5997 24397 6026 24453
rect 6082 24397 6111 24453
rect 6167 24397 6196 24453
rect 6252 24397 6280 24453
rect 6336 24397 6347 24453
rect 5758 24392 6347 24397
rect 7236 24565 7828 33634
rect 8138 24620 8730 34496
tri 18471 34303 18629 34461 se
rect 18629 34392 18718 36400
tri 18718 36336 18782 36400 nw
tri 22182 36319 22263 36400 ne
rect 22263 36345 22290 36400
tri 22290 36345 22438 36493 sw
rect 22466 36483 22532 36507
rect 22466 36427 22471 36483
rect 22527 36427 22532 36483
rect 22466 36422 22532 36427
rect 22598 36563 22664 36659
rect 22598 36507 22603 36563
rect 22659 36507 22664 36563
rect 22598 36483 22664 36507
rect 22598 36427 22603 36483
rect 22659 36427 22664 36483
rect 22598 36422 22664 36427
rect 22726 36563 22792 36790
rect 22726 36507 22731 36563
rect 22787 36507 22792 36563
rect 22726 36483 22792 36507
rect 22726 36427 22731 36483
rect 22787 36427 22792 36483
rect 22726 36422 22792 36427
rect 22852 36563 22918 36921
rect 22852 36507 22857 36563
rect 22913 36507 22918 36563
rect 22852 36483 22918 36507
rect 22852 36427 22857 36483
rect 22913 36427 22918 36483
rect 22852 36422 22918 36427
rect 22263 36319 22438 36345
tri 22263 36144 22438 36319 ne
tri 22438 36144 22639 36345 sw
tri 22438 36066 22516 36144 ne
tri 18629 34303 18718 34392 nw
tri 18313 34145 18471 34303 se
tri 18471 34145 18629 34303 nw
tri 18309 34141 18313 34145 se
rect 18313 34141 18419 34145
rect 18309 33980 18419 34141
tri 18419 34093 18471 34145 nw
rect 18309 33924 18314 33980
rect 18370 33924 18419 33980
rect 18309 33900 18419 33924
rect 18309 33844 18314 33900
rect 18370 33844 18419 33900
rect 18309 33839 18419 33844
tri 9942 33634 9947 33639 se
tri 11746 33634 11751 33639 se
tri 13550 33634 13555 33639 se
tri 15354 33634 15359 33639 se
tri 8138 24614 8144 24620 ne
rect 7236 24509 7250 24565
rect 7306 24509 7335 24565
rect 7391 24509 7420 24565
rect 7476 24509 7505 24565
rect 7561 24509 7589 24565
rect 7645 24509 7673 24565
rect 7729 24509 7757 24565
rect 7813 24509 7828 24565
rect 7236 24453 7828 24509
rect 7236 24397 7250 24453
rect 7306 24397 7335 24453
rect 7391 24397 7420 24453
rect 7476 24397 7505 24453
rect 7561 24397 7589 24453
rect 7645 24397 7673 24453
rect 7729 24397 7757 24453
rect 7813 24397 7828 24453
rect 7236 24385 7828 24397
rect 9040 24565 9632 33634
rect 9942 24620 10534 33634
tri 9942 24614 9948 24620 ne
rect 9040 24509 9054 24565
rect 9110 24509 9139 24565
rect 9195 24509 9224 24565
rect 9280 24509 9309 24565
rect 9365 24509 9394 24565
rect 9450 24509 9478 24565
rect 9534 24509 9562 24565
rect 9618 24509 9632 24565
rect 9040 24453 9632 24509
rect 9040 24397 9054 24453
rect 9110 24397 9139 24453
rect 9195 24397 9224 24453
rect 9280 24397 9309 24453
rect 9365 24397 9394 24453
rect 9450 24397 9478 24453
rect 9534 24397 9562 24453
rect 9618 24397 9632 24453
rect 9040 24392 9632 24397
rect 10844 24565 11436 33634
rect 11746 24620 12338 33634
tri 11746 24614 11752 24620 ne
rect 10844 24509 10858 24565
rect 10914 24509 10943 24565
rect 10999 24509 11028 24565
rect 11084 24509 11113 24565
rect 11169 24509 11197 24565
rect 11253 24509 11281 24565
rect 11337 24509 11365 24565
rect 11421 24509 11436 24565
rect 10844 24453 11436 24509
rect 10844 24397 10858 24453
rect 10914 24397 10943 24453
rect 10999 24397 11028 24453
rect 11084 24397 11113 24453
rect 11169 24397 11197 24453
rect 11253 24397 11281 24453
rect 11337 24397 11365 24453
rect 11421 24397 11436 24453
rect 10844 24392 11436 24397
rect 12648 24565 13240 33634
rect 13550 24620 14142 33634
tri 13870 24614 13876 24620 ne
rect 12648 24509 12657 24565
rect 12713 24509 12743 24565
rect 12799 24509 12829 24565
rect 12885 24509 12915 24565
rect 12971 24509 13000 24565
rect 13056 24509 13085 24565
rect 13141 24509 13170 24565
rect 13226 24509 13240 24565
rect 12648 24453 13240 24509
rect 12648 24397 12657 24453
rect 12713 24397 12743 24453
rect 12799 24397 12829 24453
rect 12885 24397 12915 24453
rect 12971 24397 13000 24453
rect 13056 24397 13085 24453
rect 13141 24397 13170 24453
rect 13226 24397 13240 24453
rect 12648 24392 13240 24397
rect 14452 24563 15044 33634
rect 15354 24620 15946 33634
tri 15354 24614 15360 24620 ne
rect 14452 24507 14466 24563
rect 14522 24507 14551 24563
rect 14607 24507 14636 24563
rect 14692 24507 14721 24563
rect 14777 24507 14805 24563
rect 14861 24507 14889 24563
rect 14945 24507 14973 24563
rect 15029 24507 15044 24563
rect 14452 24451 15044 24507
rect 14452 24395 14466 24451
rect 14522 24395 14551 24451
rect 14607 24395 14636 24451
rect 14692 24395 14721 24451
rect 14777 24395 14805 24451
rect 14861 24395 14889 24451
rect 14945 24395 14973 24451
rect 15029 24395 15044 24451
rect 14452 24389 15044 24395
rect 16265 24565 16852 24570
rect 16265 24509 16270 24565
rect 16326 24509 16357 24565
rect 16413 24509 16444 24565
rect 16500 24509 16531 24565
rect 16587 24509 16618 24565
rect 16674 24509 16705 24565
rect 16761 24509 16791 24565
rect 16847 24509 16852 24565
rect 16265 24453 16852 24509
rect 16265 24397 16270 24453
rect 16326 24397 16357 24453
rect 16413 24397 16444 24453
rect 16500 24397 16531 24453
rect 16587 24397 16618 24453
rect 16674 24397 16705 24453
rect 16761 24397 16791 24453
rect 16847 24397 16852 24453
rect 16265 24392 16852 24397
rect 22516 22730 22639 36144
tri 4792 21844 4853 21905 sw
rect 4853 21844 5674 21949
rect 4792 21638 5674 21844
use sky130_fd_io__gpio_ovtv2_pddrvr  sky130_fd_io__gpio_ovtv2_pddrvr_0
timestamp 1676037725
transform 1 0 170 0 1 0
box 658 12107 23573 39298
use sky130_fd_io__gpio_ovtv2_pddrvr_strong_slow  sky130_fd_io__gpio_ovtv2_pddrvr_strong_slow_0
timestamp 1676037725
transform 0 1 2950 -1 0 35104
box -191 -134 1152 12303
use sky130_fd_io__gpio_ovtv2_pddrvr_weak  sky130_fd_io__gpio_ovtv2_pddrvr_weak_0
timestamp 1676037725
transform 0 -1 15177 -1 0 35104
box -118 -108 1119 7520
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_0
timestamp 1676037725
transform 1 0 16230 0 1 33050
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_1
timestamp 1676037725
transform 1 0 9526 0 1 33050
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_2
timestamp 1676037725
transform 1 0 9014 0 1 33050
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_3
timestamp 1676037725
transform 1 0 10816 0 1 33050
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_4
timestamp 1676037725
transform 1 0 11331 0 1 33050
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_5
timestamp 1676037725
transform 1 0 12625 0 1 33050
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_6
timestamp 1676037725
transform 1 0 13132 0 1 33050
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_7
timestamp 1676037725
transform 1 0 14426 0 1 33050
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_8
timestamp 1676037725
transform 1 0 14940 0 1 33050
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_9
timestamp 1676037725
transform 1 0 7720 0 1 33050
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_10
timestamp 1676037725
transform -1 0 4566 0 1 33050
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_11
timestamp 1676037725
transform -1 0 5858 0 1 33050
box 0 0 1 1
<< labels >>
flabel comment s 658 31742 658 31742 0 FreeSans 400 180 0 0 P1G
flabel comment s 618 33116 618 33116 0 FreeSans 600 0 0 0 WEAK_PAD
flabel comment s 787 32965 787 32965 0 FreeSans 600 0 0 0 STRONG_SLOW_PAD
flabel metal2 s 17422 34493 17614 34533 3 FreeSans 520 0 0 0 PD_H[0]
port 1 nsew
flabel metal2 s 17501 34428 17501 34428 3 FreeSans 520 0 0 0 PD_H[1]
flabel metal2 s 17422 34022 17614 34074 3 FreeSans 520 0 0 0 PD_H[2]
port 2 nsew
flabel metal2 s 17422 33355 17614 33433 3 FreeSans 520 0 0 0 PD_H[3]
port 3 nsew
<< properties >>
string GDS_END 42014948
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 41969956
<< end >>
