magic
tech sky130A
magscale 1 2
timestamp 1676037725
<< nwell >>
rect 2470 420 2634 752
<< poly >>
rect 4396 970 4462 986
rect 2730 933 2796 949
rect 2730 899 2746 933
rect 2780 899 2796 933
rect 2730 865 2796 899
rect 2730 831 2746 865
rect 2780 831 2796 865
rect 2730 796 2796 831
rect 2730 762 2746 796
rect 2780 762 2796 796
rect 2730 746 2796 762
rect 2946 933 3012 949
rect 2946 899 2962 933
rect 2996 899 3012 933
rect 2946 865 3012 899
rect 2946 831 2962 865
rect 2996 831 3012 865
rect 2946 796 3012 831
rect 2946 762 2962 796
rect 2996 762 3012 796
rect 2946 746 3012 762
rect 3101 933 3167 949
rect 3101 899 3117 933
rect 3151 899 3167 933
rect 3101 865 3167 899
rect 3101 831 3117 865
rect 3151 831 3167 865
rect 3101 796 3167 831
rect 3101 762 3117 796
rect 3151 762 3167 796
rect 3101 746 3167 762
rect 3368 933 3434 949
rect 3368 899 3384 933
rect 3418 899 3434 933
rect 3368 865 3434 899
rect 3368 831 3384 865
rect 3418 831 3434 865
rect 3368 796 3434 831
rect 3368 762 3384 796
rect 3418 762 3434 796
rect 3368 746 3434 762
rect 3584 933 3650 949
rect 3584 899 3600 933
rect 3634 899 3650 933
rect 3584 865 3650 899
rect 3584 831 3600 865
rect 3634 831 3650 865
rect 3584 796 3650 831
rect 3584 762 3600 796
rect 3634 762 3650 796
rect 3584 746 3650 762
rect 3739 933 3805 949
rect 3739 899 3755 933
rect 3789 899 3805 933
rect 3739 865 3805 899
rect 3739 831 3755 865
rect 3789 831 3805 865
rect 3739 796 3805 831
rect 3739 762 3755 796
rect 3789 762 3805 796
rect 3739 746 3805 762
rect 4027 933 4093 949
rect 4027 899 4043 933
rect 4077 899 4093 933
rect 4027 865 4093 899
rect 4027 831 4043 865
rect 4077 831 4093 865
rect 4027 796 4093 831
rect 4027 762 4043 796
rect 4077 762 4093 796
rect 4027 746 4093 762
rect 4182 933 4248 949
rect 4182 899 4198 933
rect 4232 899 4248 933
rect 4182 865 4248 899
rect 4182 831 4198 865
rect 4232 831 4248 865
rect 4182 796 4248 831
rect 4182 762 4198 796
rect 4232 762 4248 796
rect 4396 936 4412 970
rect 4446 936 4462 970
rect 4396 902 4462 936
rect 4396 868 4412 902
rect 4446 868 4462 902
rect 4396 834 4462 868
rect 4396 800 4412 834
rect 4446 800 4462 834
rect 4396 784 4462 800
rect 4564 970 4630 986
rect 4564 936 4580 970
rect 4614 936 4630 970
rect 4564 902 4630 936
rect 4564 868 4580 902
rect 4614 868 4630 902
rect 4564 834 4630 868
rect 4564 800 4580 834
rect 4614 800 4630 834
rect 4564 784 4630 800
rect 4848 933 4914 949
rect 4848 899 4864 933
rect 4898 899 4914 933
rect 4848 865 4914 899
rect 4848 831 4864 865
rect 4898 831 4914 865
rect 4848 796 4914 831
rect 4182 746 4248 762
rect 4848 762 4864 796
rect 4898 762 4914 796
rect 4848 746 4914 762
rect 5064 933 5130 949
rect 5064 899 5080 933
rect 5114 899 5130 933
rect 5064 865 5130 899
rect 5064 831 5080 865
rect 5114 831 5130 865
rect 5064 796 5130 831
rect 5064 762 5080 796
rect 5114 762 5130 796
rect 5064 746 5130 762
rect 5310 933 5376 949
rect 5310 899 5326 933
rect 5360 899 5376 933
rect 5310 865 5376 899
rect 5310 831 5326 865
rect 5360 831 5376 865
rect 5310 796 5376 831
rect 5310 762 5326 796
rect 5360 762 5376 796
rect 5310 746 5376 762
rect 5526 933 5592 949
rect 5526 899 5542 933
rect 5576 899 5592 933
rect 5526 865 5592 899
rect 5526 831 5542 865
rect 5576 831 5592 865
rect 5526 796 5592 831
rect 5526 762 5542 796
rect 5576 762 5592 796
rect 5526 746 5592 762
rect 5820 933 5886 949
rect 5820 899 5836 933
rect 5870 899 5886 933
rect 5820 865 5886 899
rect 5820 831 5836 865
rect 5870 831 5886 865
rect 5820 796 5886 831
rect 5820 762 5836 796
rect 5870 762 5886 796
rect 5820 746 5886 762
rect 5956 933 6022 949
rect 5956 899 5972 933
rect 6006 899 6022 933
rect 5956 865 6022 899
rect 5956 831 5972 865
rect 6006 831 6022 865
rect 5956 796 6022 831
rect 5956 762 5972 796
rect 6006 762 6022 796
rect 5956 746 6022 762
rect 6172 933 6238 949
rect 6172 899 6188 933
rect 6222 899 6238 933
rect 6172 865 6238 899
rect 6172 831 6188 865
rect 6222 831 6238 865
rect 6172 796 6238 831
rect 6172 762 6188 796
rect 6222 762 6238 796
rect 6172 746 6238 762
rect 6308 933 6374 949
rect 6308 899 6324 933
rect 6358 899 6374 933
rect 6308 865 6374 899
rect 6308 831 6324 865
rect 6358 831 6374 865
rect 6308 796 6374 831
rect 6308 762 6324 796
rect 6358 762 6374 796
rect 6308 746 6374 762
<< polycont >>
rect 2746 899 2780 933
rect 2746 831 2780 865
rect 2746 762 2780 796
rect 2962 899 2996 933
rect 2962 831 2996 865
rect 2962 762 2996 796
rect 3117 899 3151 933
rect 3117 831 3151 865
rect 3117 762 3151 796
rect 3384 899 3418 933
rect 3384 831 3418 865
rect 3384 762 3418 796
rect 3600 899 3634 933
rect 3600 831 3634 865
rect 3600 762 3634 796
rect 3755 899 3789 933
rect 3755 831 3789 865
rect 3755 762 3789 796
rect 4043 899 4077 933
rect 4043 831 4077 865
rect 4043 762 4077 796
rect 4198 899 4232 933
rect 4198 831 4232 865
rect 4198 762 4232 796
rect 4412 936 4446 970
rect 4412 868 4446 902
rect 4412 800 4446 834
rect 4580 936 4614 970
rect 4580 868 4614 902
rect 4580 800 4614 834
rect 4864 899 4898 933
rect 4864 831 4898 865
rect 4864 762 4898 796
rect 5080 899 5114 933
rect 5080 831 5114 865
rect 5080 762 5114 796
rect 5326 899 5360 933
rect 5326 831 5360 865
rect 5326 762 5360 796
rect 5542 899 5576 933
rect 5542 831 5576 865
rect 5542 762 5576 796
rect 5836 899 5870 933
rect 5836 831 5870 865
rect 5836 762 5870 796
rect 5972 899 6006 933
rect 5972 831 6006 865
rect 5972 762 6006 796
rect 6188 899 6222 933
rect 6188 831 6222 865
rect 6188 762 6222 796
rect 6324 899 6358 933
rect 6324 831 6358 865
rect 6324 762 6358 796
<< locali >>
rect 5128 1270 5278 1336
rect 2254 850 2328 1090
rect 2746 933 2780 949
rect 2746 865 2780 899
rect 2854 908 2888 946
rect 2962 933 2996 949
rect 3117 933 3151 949
rect 2746 796 2780 831
rect 2746 746 2780 762
rect 2962 865 2996 899
rect 2962 796 2996 831
rect 3030 834 3064 872
rect 3117 865 3151 899
rect 2962 746 2996 762
rect 3117 798 3122 831
rect 3156 798 3194 832
rect 3117 796 3151 798
rect 3117 746 3151 762
rect 2943 308 2977 346
rect 3030 376 3064 414
rect 2678 234 2712 272
rect 3274 114 3316 1236
rect 3384 933 3418 949
rect 3384 865 3418 899
rect 3492 908 3526 946
rect 3600 933 3634 949
rect 3755 933 3789 949
rect 3384 796 3418 831
rect 3384 746 3418 762
rect 3600 865 3634 899
rect 3600 796 3634 831
rect 3668 834 3702 872
rect 3940 906 3974 1236
rect 4412 970 4446 986
rect 4043 933 4077 949
rect 3755 865 3789 899
rect 3600 746 3634 762
rect 3755 796 3789 831
rect 3844 834 3878 872
rect 3940 872 3954 906
rect 3940 834 3988 872
rect 3940 800 3954 834
rect 4198 933 4232 949
rect 4043 865 4077 899
rect 3755 746 3789 762
rect 4043 796 4077 831
rect 4130 834 4164 872
rect 4198 865 4232 899
rect 4043 746 4077 762
rect 4198 796 4232 831
rect 4412 905 4446 936
rect 4412 834 4446 868
rect 4198 746 4232 762
rect 4306 758 4340 796
rect 4412 784 4446 799
rect 4580 970 4614 986
rect 4580 902 4614 936
rect 4580 834 4614 868
rect 4864 933 4898 949
rect 4864 865 4898 899
rect 4580 784 4614 800
rect 4686 758 4720 796
rect 4864 796 4898 831
rect 5080 933 5114 949
rect 5080 865 5114 899
rect 4864 746 4898 762
rect 4972 758 5006 796
rect 5080 796 5114 831
rect 5080 746 5114 762
rect 5244 905 5278 1270
rect 5326 933 5360 949
rect 5244 871 5249 905
rect 5244 833 5283 871
rect 5244 799 5249 833
rect 5326 865 5360 899
rect 3405 376 3439 414
rect 4130 308 4164 346
rect 4883 296 4917 334
rect 3578 234 3612 272
rect 5148 296 5182 334
rect 3245 87 3316 114
rect 4796 138 4830 176
rect 3245 -11 3311 87
rect 3370 -12 3472 54
rect 3718 -12 3722 54
rect 3758 -3 3796 31
rect 4038 20 4076 54
rect 4584 21 4622 55
rect 5244 53 5278 799
rect 5326 796 5360 831
rect 5326 746 5360 762
rect 5542 933 5576 949
rect 5542 865 5576 899
rect 5542 796 5576 831
rect 5542 746 5576 762
rect 5836 933 5870 949
rect 5836 865 5870 899
rect 5836 796 5870 831
rect 5836 746 5870 762
rect 5972 933 6006 949
rect 5972 865 6006 899
rect 5972 796 6006 831
rect 5972 746 6006 762
rect 6188 933 6222 949
rect 6188 865 6222 899
rect 6188 796 6222 831
rect 6188 746 6222 762
rect 6324 933 6358 949
rect 6324 865 6358 899
rect 6324 796 6358 831
rect 6324 746 6358 762
rect 5343 58 5377 96
rect 4004 -12 4008 20
rect 5128 -12 5278 53
rect 5312 24 5343 54
rect 5377 24 5414 54
rect 5312 -12 5414 24
rect 2732 -29 2834 -12
rect 2762 -63 2800 -29
rect 2732 -77 2834 -63
rect 4184 -49 4286 -12
rect 4218 -83 4256 -49
<< viali >>
rect 2854 946 2888 980
rect 2854 874 2888 908
rect 3030 872 3064 906
rect 3030 800 3064 834
rect 3122 831 3151 832
rect 3151 831 3156 832
rect 3122 798 3156 831
rect 3194 798 3228 832
rect 3030 414 3064 448
rect 2943 346 2977 380
rect 3030 342 3064 376
rect 2678 272 2712 306
rect 2943 274 2977 308
rect 2678 200 2712 234
rect 3492 946 3526 980
rect 3492 874 3526 908
rect 3668 872 3702 906
rect 3668 800 3702 834
rect 3844 872 3878 906
rect 3844 800 3878 834
rect 3954 872 3988 906
rect 3954 800 3988 834
rect 4130 872 4164 906
rect 4130 800 4164 834
rect 4412 902 4446 905
rect 4412 871 4446 902
rect 4306 796 4340 830
rect 4412 800 4446 833
rect 4412 799 4446 800
rect 4686 796 4720 830
rect 4306 724 4340 758
rect 4686 724 4720 758
rect 4972 796 5006 830
rect 4972 724 5006 758
rect 5249 871 5283 905
rect 5249 799 5283 833
rect 3405 414 3439 448
rect 3405 342 3439 376
rect 4130 346 4164 380
rect 3578 272 3612 306
rect 4130 274 4164 308
rect 4883 334 4917 368
rect 4883 262 4917 296
rect 5148 334 5182 368
rect 5148 262 5182 296
rect 3578 200 3612 234
rect 4796 176 4830 210
rect 4796 104 4830 138
rect 3724 -3 3758 31
rect 3796 -3 3830 31
rect 4004 20 4038 54
rect 4076 20 4110 54
rect 4550 21 4584 55
rect 4622 21 4656 55
rect 5343 96 5377 130
rect 5343 24 5377 58
rect 2728 -63 2762 -29
rect 2800 -63 2834 -29
rect 4184 -83 4218 -49
rect 4256 -83 4290 -49
<< metal1 >>
rect 1183 1014 1210 1216
rect 2408 1014 2695 1216
rect 3252 1014 3333 1216
rect 3480 1014 3538 1216
rect 3890 1014 3942 1216
rect 4732 1014 4813 1216
rect 5165 1014 5275 1216
rect 5451 1014 5480 1216
rect 3480 986 5480 1014
rect 1051 940 2761 986
rect 2842 980 2900 986
rect 2842 946 2854 980
rect 2888 946 2900 980
tri 2817 915 2842 940 ne
rect 2190 884 2447 912
rect 2441 860 2447 884
rect 2499 860 2511 912
rect 2563 860 2569 912
rect 2842 908 2900 946
rect 3252 940 3333 986
rect 3480 980 3538 986
rect 3480 946 3492 980
rect 3526 946 3538 980
tri 2900 915 2925 940 nw
rect 2356 810 2403 856
tri 2403 810 2449 856 sw
tri 2603 852 2642 891 se
rect 2642 852 2648 904
rect 2700 852 2712 904
rect 2764 852 2770 904
rect 2842 874 2854 908
rect 2888 874 2900 908
rect 2842 868 2900 874
rect 3018 906 3076 912
rect 3018 872 3030 906
rect 3064 872 3076 906
tri 3432 892 3480 940 ne
rect 3480 908 3538 946
rect 3890 940 3942 986
rect 4732 940 4813 986
rect 5165 940 5275 986
rect 5451 940 5480 986
tri 2390 756 2444 810 ne
rect 2444 802 2449 810
tri 2449 802 2457 810 sw
tri 2553 802 2603 852 se
rect 2603 802 2606 852
rect 2444 789 2606 802
tri 2606 789 2669 852 nw
rect 3018 834 3076 872
rect 3480 874 3492 908
rect 3526 874 3538 908
rect 3480 868 3538 874
rect 3656 906 3714 912
rect 3656 872 3668 906
rect 3702 872 3714 906
rect 3018 800 3030 834
rect 3064 800 3076 834
rect 3018 794 3076 800
rect 3110 832 3240 838
rect 3110 798 3122 832
rect 3156 798 3194 832
rect 3228 829 3240 832
rect 3656 834 3714 872
rect 3832 906 3890 912
rect 3832 872 3844 906
rect 3878 872 3890 906
tri 3714 841 3739 866 nw
tri 3807 841 3832 866 ne
rect 3656 829 3668 834
rect 3228 800 3668 829
rect 3702 800 3714 834
rect 3228 798 3714 800
rect 3110 792 3240 798
rect 3656 794 3714 798
rect 3832 834 3890 872
rect 3832 800 3844 834
rect 3878 800 3890 834
rect 3832 794 3890 800
rect 3942 906 4000 912
rect 3942 872 3954 906
rect 3988 872 4000 906
rect 3942 834 4000 872
rect 4118 906 4176 912
rect 4118 872 4130 906
rect 4164 872 4176 906
tri 4000 841 4025 866 nw
tri 4093 841 4118 866 ne
rect 3942 800 3954 834
rect 3988 800 4000 834
rect 3942 794 4000 800
rect 4118 834 4176 872
rect 4400 905 5295 911
rect 4400 904 4412 905
rect 4446 904 5249 905
rect 4400 852 4406 904
rect 4458 852 4470 904
rect 4522 883 5249 904
rect 4522 852 4528 883
tri 4528 852 4559 883 nw
tri 5212 858 5237 883 ne
rect 5237 871 5249 883
rect 5283 871 5295 905
rect 4118 800 4130 834
rect 4164 800 4176 834
rect 4118 794 4176 800
rect 4294 830 4352 836
rect 4294 796 4306 830
rect 4340 796 4352 830
rect 2444 756 2573 789
tri 2573 756 2606 789 nw
tri 4269 764 4294 789 se
rect 2622 718 3538 764
rect 3890 718 3942 764
rect 4294 758 4352 796
rect 4400 833 4458 852
rect 4400 799 4412 833
rect 4446 799 4458 833
rect 4400 793 4458 799
rect 4674 830 4732 836
rect 4674 796 4686 830
rect 4720 796 4732 830
tri 4352 764 4377 789 sw
tri 4649 764 4674 789 se
rect 4674 764 4732 796
rect 4960 830 5018 836
rect 4960 796 4972 830
rect 5006 796 5018 830
tri 4732 764 4757 789 sw
tri 4935 764 4960 789 se
rect 4294 724 4306 758
rect 4340 724 4352 758
rect 4294 718 4352 724
rect 4674 758 4813 764
rect 4674 724 4686 758
rect 4720 724 4813 758
rect 4674 718 4813 724
rect 4960 758 5018 796
rect 5237 833 5295 871
rect 5237 799 5249 833
rect 5283 799 5295 833
rect 5237 793 5295 799
tri 5018 764 5043 789 sw
rect 4960 724 4972 758
rect 5006 724 5018 758
rect 4960 718 5018 724
rect 5165 718 5275 764
rect 5451 718 5480 764
rect 2622 690 5480 718
rect 2622 676 2695 690
rect 2341 488 2695 676
rect 3252 488 3333 690
rect 3480 488 3538 690
rect 3890 488 3942 690
rect 4732 488 4813 690
rect 5165 488 5275 690
rect 5451 488 5480 690
rect 3024 448 3445 460
rect 3024 414 3030 448
rect 3064 414 3405 448
rect 3439 414 3445 448
rect 3024 408 3445 414
rect 4516 408 5480 460
rect 2937 380 2983 392
rect 2937 346 2943 380
rect 2977 346 2983 380
rect 2672 306 2718 318
rect 2672 272 2678 306
rect 2712 272 2718 306
rect 2672 234 2718 272
rect 2937 308 2983 346
rect 3024 376 3070 408
tri 3070 383 3095 408 nw
tri 3374 383 3399 408 ne
rect 3024 342 3030 376
rect 3064 342 3070 376
rect 3024 330 3070 342
rect 3399 376 3445 408
rect 3399 342 3405 376
rect 3439 342 3445 376
tri 3516 360 3544 388 se
rect 3544 360 3710 388
tri 3710 360 3738 388 sw
rect 4124 380 4170 392
tri 4726 383 4751 408 nw
rect 3399 330 3445 342
tri 3490 334 3516 360 se
rect 3516 348 3738 360
rect 3516 334 3528 348
rect 2937 274 2943 308
rect 2977 302 2983 308
tri 3458 302 3490 334 se
rect 3490 318 3528 334
tri 3528 318 3558 348 nw
rect 3490 302 3512 318
tri 3512 302 3528 318 nw
rect 3572 306 3618 318
rect 2977 274 3472 302
rect 2937 262 3472 274
tri 3472 262 3512 302 nw
rect 3572 272 3578 306
rect 3612 272 3618 306
tri 3692 302 3738 348 ne
tri 3738 302 3796 360 sw
rect 4124 346 4130 380
rect 4164 346 4170 380
rect 4124 308 4170 346
rect 4877 368 4923 380
rect 4877 334 4883 368
rect 4917 334 4923 368
rect 4124 302 4130 308
rect 3572 234 3618 272
tri 3738 262 3778 302 ne
rect 3778 274 4130 302
rect 4164 274 4170 308
tri 4852 302 4877 327 se
rect 4877 302 4923 334
rect 5142 368 5188 380
rect 5142 334 5148 368
rect 5182 334 5188 368
tri 4923 302 4948 327 sw
tri 5117 302 5142 327 se
rect 5142 302 5188 334
tri 5188 302 5213 327 sw
rect 3778 262 4170 274
rect 4548 296 5480 302
rect 4548 262 4883 296
rect 4917 262 5148 296
rect 5182 262 5480 296
rect 4548 250 5480 262
rect 2672 200 2678 234
rect 2712 200 3578 234
rect 3612 200 3618 234
rect 2672 188 3618 200
rect 4548 210 5480 222
rect 2441 127 2447 179
rect 2499 127 2511 179
rect 2563 160 2569 179
rect 4548 176 4796 210
rect 4830 176 5480 210
rect 4548 170 5480 176
rect 2563 127 4359 160
tri 4330 98 4359 127 ne
tri 4359 123 4396 160 sw
tri 4765 145 4790 170 ne
rect 4790 138 4836 170
tri 4836 145 4861 170 nw
rect 4359 98 4396 123
rect 3991 54 4126 68
tri 4359 61 4396 98 ne
tri 4396 61 4458 123 sw
rect 4790 104 4796 138
rect 4830 104 4836 138
rect 4790 92 4836 104
rect 5337 130 5383 142
rect 5337 96 5343 130
rect 5377 96 5383 130
rect 3712 31 3842 43
rect 3712 -3 3724 31
rect 3758 -3 3796 31
rect 3830 -3 3842 31
rect 3991 20 4004 54
rect 4038 20 4076 54
rect 4110 20 4126 54
rect 3991 8 4126 20
tri 4396 15 4442 61 ne
rect 4442 55 4668 61
rect 4442 21 4550 55
rect 4584 21 4622 55
rect 4656 21 4668 55
rect 4442 15 4668 21
rect 5337 58 5383 96
rect 5337 24 5343 58
rect 5377 24 5383 58
rect 5337 12 5383 24
rect 3712 -9 3842 -3
rect 2716 -29 2846 -23
rect 2716 -63 2728 -29
rect 2762 -63 2800 -29
rect 2834 -37 2846 -29
rect 2834 -49 5418 -37
rect 2834 -63 4184 -49
rect 2716 -69 4184 -63
rect 4178 -83 4184 -69
rect 4218 -83 4256 -49
rect 4290 -69 5418 -49
rect 4290 -83 4296 -69
rect 4178 -95 4296 -83
<< via1 >>
rect 2447 860 2499 912
rect 2511 860 2563 912
rect 2648 852 2700 904
rect 2712 852 2764 904
rect 4406 871 4412 904
rect 4412 871 4446 904
rect 4446 871 4458 904
rect 4406 852 4458 871
rect 4470 852 4522 904
rect 2447 127 2499 179
rect 2511 127 2563 179
<< metal2 >>
rect 2441 860 2447 912
rect 2499 860 2511 912
rect 2563 860 2569 912
rect 2441 179 2569 860
rect 2642 852 2648 904
rect 2700 852 2712 904
rect 2764 852 4406 904
rect 4458 852 4470 904
rect 4522 852 4528 904
rect 2441 127 2447 179
rect 2499 127 2511 179
rect 2563 127 2569 179
use sky130_fd_io__sio_hotswap_dly_ovtv2  sky130_fd_io__sio_hotswap_dly_ovtv2_0
timestamp 1676037725
transform -1 0 2576 0 -1 1264
box 88 0 2560 844
use sky130_fd_io__sio_hvsbt_inv_x1  sky130_fd_io__sio_hvsbt_inv_x1_0
timestamp 1676037725
transform -1 0 2871 0 -1 1357
box -107 21 267 1369
use sky130_fd_io__sio_hvsbt_inv_x1  sky130_fd_io__sio_hvsbt_inv_x1_1
timestamp 1676037725
transform -1 0 3509 0 -1 1357
box -107 21 267 1369
use sky130_fd_io__sio_hvsbt_inv_x1  sky130_fd_io__sio_hvsbt_inv_x1_2
timestamp 1676037725
transform -1 0 4989 0 -1 1357
box -107 21 267 1369
use sky130_fd_io__sio_hvsbt_inv_x1  sky130_fd_io__sio_hvsbt_inv_x1_3
timestamp 1676037725
transform 1 0 4989 0 -1 1357
box -107 21 267 1369
use sky130_fd_io__sio_hvsbt_inv_x1  sky130_fd_io__sio_hvsbt_inv_x1_4
timestamp 1676037725
transform -1 0 5451 0 -1 1357
box -107 21 267 1369
use sky130_fd_io__sio_hvsbt_nand2  sky130_fd_io__sio_hvsbt_nand2_0
timestamp 1676037725
transform 1 0 2871 0 -1 1357
box -107 21 459 1369
use sky130_fd_io__sio_hvsbt_nand2  sky130_fd_io__sio_hvsbt_nand2_1
timestamp 1676037725
transform -1 0 4323 0 -1 1357
box -107 21 459 1369
use sky130_fd_io__sio_hvsbt_nand2  sky130_fd_io__sio_hvsbt_nand2_2
timestamp 1676037725
transform 1 0 3509 0 -1 1357
box -107 21 459 1369
use sky130_fd_io__sio_hvsbt_nor  sky130_fd_io__sio_hvsbt_nor_0
timestamp 1676037725
transform 1 0 4323 0 -1 1357
box -107 21 487 1369
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_0
timestamp 1676037725
transform 0 1 3030 -1 0 448
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_1
timestamp 1676037725
transform 0 1 3405 -1 0 448
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_2
timestamp 1676037725
transform 0 -1 4830 1 0 104
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_3
timestamp 1676037725
transform 0 -1 4917 1 0 262
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_4
timestamp 1676037725
transform 0 -1 5182 1 0 262
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180878  sky130_fd_pr__via_l1m1__example_5595914180878_0
timestamp 1676037725
transform -1 0 3526 0 1 874
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180878  sky130_fd_pr__via_l1m1__example_5595914180878_1
timestamp 1676037725
transform -1 0 2888 0 1 874
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180878  sky130_fd_pr__via_l1m1__example_5595914180878_2
timestamp 1676037725
transform 1 0 3030 0 1 800
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180878  sky130_fd_pr__via_l1m1__example_5595914180878_3
timestamp 1676037725
transform -1 0 5006 0 1 724
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180878  sky130_fd_pr__via_l1m1__example_5595914180878_4
timestamp 1676037725
transform -1 0 4720 0 1 724
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180878  sky130_fd_pr__via_l1m1__example_5595914180878_5
timestamp 1676037725
transform 0 1 4004 -1 0 54
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180878  sky130_fd_pr__via_l1m1__example_5595914180878_6
timestamp 1676037725
transform 0 1 4184 -1 0 -49
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180878  sky130_fd_pr__via_l1m1__example_5595914180878_7
timestamp 1676037725
transform -1 0 4340 0 1 724
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180878  sky130_fd_pr__via_l1m1__example_5595914180878_8
timestamp 1676037725
transform -1 0 4446 0 1 799
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180878  sky130_fd_pr__via_l1m1__example_5595914180878_9
timestamp 1676037725
transform -1 0 5283 0 1 799
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180878  sky130_fd_pr__via_l1m1__example_5595914180878_10
timestamp 1676037725
transform 1 0 4130 0 1 800
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180878  sky130_fd_pr__via_l1m1__example_5595914180878_11
timestamp 1676037725
transform -1 0 3702 0 1 800
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180878  sky130_fd_pr__via_l1m1__example_5595914180878_12
timestamp 1676037725
transform 1 0 3954 0 1 800
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180878  sky130_fd_pr__via_l1m1__example_5595914180878_13
timestamp 1676037725
transform 1 0 3844 0 1 800
box 0 0 1 1
<< labels >>
flabel metal1 s 5451 940 5480 986 0 FreeSans 200 0 0 0 VGND
port 2 nsew
flabel metal1 s 5434 408 5480 460 0 FreeSans 200 0 0 0 EXITHS_H
port 3 nsew
flabel metal1 s 4019 29 4058 57 0 FreeSans 200 0 0 0 EN_H
port 4 nsew
flabel metal1 s 3759 -9 3801 19 0 FreeSans 200 0 0 0 FORCEHI_H[1]
port 5 nsew
flabel metal1 s 5316 -69 5418 -37 0 FreeSans 200 0 0 0 OD_H
port 6 nsew
flabel metal1 s 3480 488 3509 764 0 FreeSans 200 0 0 0 VCC_IO
port 7 nsew
flabel metal1 s 5451 488 5480 764 0 FreeSans 200 0 0 0 VCC_IO
port 7 nsew
flabel metal1 s 5451 1014 5480 1216 0 FreeSans 200 0 0 0 VGND
port 2 nsew
flabel metal1 s 3480 1014 3509 1216 0 FreeSans 200 0 0 0 VGND
port 2 nsew
flabel metal1 s 3480 940 3509 986 0 FreeSans 200 0 0 0 VGND
port 2 nsew
flabel metal1 s 4548 170 4594 222 0 FreeSans 200 0 0 0 ENHS_H
port 8 nsew
flabel metal1 s 5434 170 5480 222 0 FreeSans 200 0 0 0 ENHS_H
port 8 nsew
flabel metal1 s 5434 250 5480 302 0 FreeSans 200 0 0 0 ENHS_H_N
port 9 nsew
flabel metal1 s 4548 250 4594 302 0 FreeSans 200 0 0 0 ENHS_H_N
port 9 nsew
flabel metal1 s 4548 408 4594 460 0 FreeSans 200 0 0 0 EXITHS_H
port 3 nsew
flabel metal1 s 3509 940 3538 986 0 FreeSans 200 0 0 0 VGND
port 2 nsew
flabel metal1 s 3509 1014 3538 1216 0 FreeSans 200 0 0 0 VGND
port 2 nsew
flabel metal1 s 2080 718 2080 718 0 FreeSans 440 0 0 0 ENHS_DLY_H
flabel metal1 s 2602 940 2622 986 0 FreeSans 200 0 0 0 VGND
port 2 nsew
flabel metal1 s 2602 1014 2622 1216 0 FreeSans 200 0 0 0 VGND
port 2 nsew
flabel metal1 s 2635 488 2661 764 0 FreeSans 200 0 0 0 VCC_IO
port 7 nsew
flabel locali s 3245 -11 3311 50 0 FreeSans 200 180 0 0 DISHS_H_N
port 10 nsew
flabel locali s 5312 -12 5414 54 0 FreeSans 200 0 0 0 ENHS_LAT_H_N
port 11 nsew
flabel locali s 3370 -12 3472 54 0 FreeSans 200 180 0 0 DISHS_H
port 12 nsew
flabel locali s 3421 21 3421 21 0 FreeSans 200 0 0 0 DISHS_H
<< properties >>
string GDS_END 34133412
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 34112488
<< end >>
