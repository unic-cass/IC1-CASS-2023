* NGSPICE file created from wb_buttons_leds.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_2 abstract view
.subckt sky130_fd_sc_hd__a311oi_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_4 abstract view
.subckt sky130_fd_sc_hd__o32ai_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_4 abstract view
.subckt sky130_fd_sc_hd__a21bo_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_2 abstract view
.subckt sky130_fd_sc_hd__a32oi_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_4 abstract view
.subckt sky130_fd_sc_hd__o32a_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_1 abstract view
.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_1 abstract view
.subckt sky130_fd_sc_hd__nor2b_1 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_2 abstract view
.subckt sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_1 abstract view
.subckt sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_2 abstract view
.subckt sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd1_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd1_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s4s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s4s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_4 abstract view
.subckt sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_4 abstract view
.subckt sky130_fd_sc_hd__or2b_4 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_4 abstract view
.subckt sky130_fd_sc_hd__o311a_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_4 abstract view
.subckt sky130_fd_sc_hd__o311ai_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

.subckt wb_buttons_leds VGND VPWR buttons clk i_wb_addr[0] i_wb_addr[10] i_wb_addr[11]
+ i_wb_addr[12] i_wb_addr[13] i_wb_addr[14] i_wb_addr[15] i_wb_addr[16] i_wb_addr[17]
+ i_wb_addr[18] i_wb_addr[19] i_wb_addr[1] i_wb_addr[20] i_wb_addr[21] i_wb_addr[22]
+ i_wb_addr[23] i_wb_addr[24] i_wb_addr[25] i_wb_addr[26] i_wb_addr[27] i_wb_addr[28]
+ i_wb_addr[29] i_wb_addr[2] i_wb_addr[30] i_wb_addr[31] i_wb_addr[3] i_wb_addr[4]
+ i_wb_addr[5] i_wb_addr[6] i_wb_addr[7] i_wb_addr[8] i_wb_addr[9] i_wb_cyc i_wb_data[0]
+ i_wb_data[10] i_wb_data[11] i_wb_data[12] i_wb_data[13] i_wb_data[14] i_wb_data[15]
+ i_wb_data[16] i_wb_data[17] i_wb_data[18] i_wb_data[19] i_wb_data[1] i_wb_data[20]
+ i_wb_data[21] i_wb_data[22] i_wb_data[23] i_wb_data[24] i_wb_data[25] i_wb_data[26]
+ i_wb_data[27] i_wb_data[28] i_wb_data[29] i_wb_data[2] i_wb_data[30] i_wb_data[31]
+ i_wb_data[3] i_wb_data[4] i_wb_data[5] i_wb_data[6] i_wb_data[7] i_wb_data[8] i_wb_data[9]
+ i_wb_stb i_wb_we led_enb[0] led_enb[1] led_enb[2] led_enb[3] led_enb[4] led_enb[5]
+ led_enb[6] led_enb[7] led_enb[8] led_enb[9] leds[0] leds[10] leds[11] leds[1] leds[2]
+ leds[3] leds[4] leds[5] leds[6] leds[7] leds[8] leds[9] o_wb_ack o_wb_data[0] o_wb_data[10]
+ o_wb_data[11] o_wb_data[12] o_wb_data[13] o_wb_data[14] o_wb_data[15] o_wb_data[16]
+ o_wb_data[17] o_wb_data[18] o_wb_data[19] o_wb_data[1] o_wb_data[20] o_wb_data[21]
+ o_wb_data[22] o_wb_data[23] o_wb_data[24] o_wb_data[25] o_wb_data[26] o_wb_data[27]
+ o_wb_data[28] o_wb_data[29] o_wb_data[2] o_wb_data[30] o_wb_data[31] o_wb_data[3]
+ o_wb_data[4] o_wb_data[5] o_wb_data[6] o_wb_data[7] o_wb_data[8] o_wb_data[9] o_wb_stall
+ reset led_enb[11] led_enb[10]
XFILLER_0_94_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09671_ _05834_ _05888_ _05899_ _05910_ _05921_ VGND VGND VPWR VPWR _05932_ sky130_fd_sc_hd__a32o_1
X_18869_ clknet_4_7_0_clk _00035_ VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_474 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_143_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09938_ _05573_ _05649_ _06722_ _05693_ VGND VGND VPWR VPWR _08832_ sky130_fd_sc_hd__and4_1
X_09869_ _08060_ _08071_ _05682_ _06062_ VGND VGND VPWR VPWR _08082_ sky130_fd_sc_hd__and4b_1
XFILLER_0_99_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11900_ _01902_ _01901_ VGND VGND VPWR VPWR _01993_ sky130_fd_sc_hd__nand2_1
X_12880_ _02972_ VGND VGND VPWR VPWR _02973_ sky130_fd_sc_hd__clkbuf_4
XTAP_2501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11831_ _05399_ _05355_ _00217_ _00909_ VGND VGND VPWR VPWR _01924_ sky130_fd_sc_hd__nand4_1
XTAP_2534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14550_ _04773_ _04774_ VGND VGND VPWR VPWR _04775_ sky130_fd_sc_hd__xor2_2
XFILLER_0_67_133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11762_ _01853_ _01854_ VGND VGND VPWR VPWR _01855_ sky130_fd_sc_hd__xnor2_2
XTAP_1844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13501_ _06711_ _00509_ VGND VGND VPWR VPWR _03628_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10713_ ApproximateM_inst.lob_16.lob2.genblk1\[10\].genblk1.mux.sel VGND VGND VPWR
+ VPWR _00806_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_95_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14481_ _04608_ _04609_ _04625_ VGND VGND VPWR VPWR _04699_ sky130_fd_sc_hd__nand3_1
XFILLER_0_82_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11693_ _01781_ _01782_ _01741_ _01756_ VGND VGND VPWR VPWR _01786_ sky130_fd_sc_hd__o211ai_2
XTAP_1899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16220_ _03239_ _06418_ VGND VGND VPWR VPWR _06589_ sky130_fd_sc_hd__or2_1
X_13432_ _03043_ _03113_ _01677_ VGND VGND VPWR VPWR _03554_ sky130_fd_sc_hd__mux2_1
X_10644_ _00719_ _00720_ _00735_ _00736_ VGND VGND VPWR VPWR _00737_ sky130_fd_sc_hd__o211a_1
XFILLER_0_36_564 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_125_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16151_ _03126_ _06512_ _06513_ VGND VGND VPWR VPWR _06514_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_141_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10575_ _07080_ cla_inst.in1\[30\] _07755_ _07047_ VGND VGND VPWR VPWR _00668_ sky130_fd_sc_hd__a22o_1
XFILLER_0_51_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13363_ _03475_ _03477_ VGND VGND VPWR VPWR _03478_ sky130_fd_sc_hd__xor2_1
XFILLER_0_24_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer7 net169 VGND VGND VPWR VPWR net170 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_106_452 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15102_ _05375_ _05376_ VGND VGND VPWR VPWR _05378_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_2_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12314_ _02357_ VGND VGND VPWR VPWR _02407_ sky130_fd_sc_hd__inv_2
X_16082_ _03311_ _06368_ _06438_ VGND VGND VPWR VPWR _06440_ sky130_fd_sc_hd__and3_1
X_13294_ _03396_ _03400_ _03401_ VGND VGND VPWR VPWR _03402_ sky130_fd_sc_hd__and3_1
XFILLER_0_106_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15033_ _05198_ _05202_ _05196_ VGND VGND VPWR VPWR _05303_ sky130_fd_sc_hd__o21a_1
X_12245_ _05747_ _00878_ _02337_ _02245_ VGND VGND VPWR VPWR _02338_ sky130_fd_sc_hd__a22oi_1
X_12176_ _02265_ _02267_ VGND VGND VPWR VPWR _02269_ sky130_fd_sc_hd__nand2_1
X_11127_ _00514_ _00813_ VGND VGND VPWR VPWR _01220_ sky130_fd_sc_hd__nor2_2
X_16984_ _06874_ _06957_ VGND VGND VPWR VPWR _07420_ sky130_fd_sc_hd__or2_1
X_11058_ ApproximateM_inst.lob_16.lob2.genblk2.mux_final.sel VGND VGND VPWR VPWR _01151_
+ sky130_fd_sc_hd__clkbuf_4
X_18723_ _00516_ _09183_ net69 VGND VGND VPWR VPWR _09249_ sky130_fd_sc_hd__a21oi_1
X_15935_ _06272_ _06280_ VGND VGND VPWR VPWR _06281_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_3_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10009_ cla_inst.in2\[25\] VGND VGND VPWR VPWR _09352_ sky130_fd_sc_hd__buf_2
X_18654_ net62 _03086_ _09193_ VGND VGND VPWR VPWR _09199_ sky130_fd_sc_hd__mux2_1
X_15866_ _06157_ _06205_ _06206_ VGND VGND VPWR VPWR _06207_ sky130_fd_sc_hd__or3_1
X_17605_ _08086_ _08096_ VGND VGND VPWR VPWR _08097_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_149_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14817_ _04965_ _04966_ _05065_ _05066_ VGND VGND VPWR VPWR _05067_ sky130_fd_sc_hd__o211ai_4
X_18585_ salida\[12\] _09141_ _09142_ salida\[44\] _09146_ VGND VGND VPWR VPWR _09148_
+ sky130_fd_sc_hd__a221o_1
X_15797_ _06131_ _06132_ VGND VGND VPWR VPWR _06133_ sky130_fd_sc_hd__and2_1
XFILLER_0_58_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17536_ _02846_ _02847_ _08021_ VGND VGND VPWR VPWR _08022_ sky130_fd_sc_hd__o21a_2
XFILLER_0_147_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14748_ _04854_ _04859_ _04852_ VGND VGND VPWR VPWR _04991_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_58_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_522 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17467_ _06969_ net145 VGND VGND VPWR VPWR _07946_ sky130_fd_sc_hd__nand2_1
X_14679_ _04750_ _04915_ VGND VGND VPWR VPWR _04916_ sky130_fd_sc_hd__xor2_1
XFILLER_0_7_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16418_ sel_op\[2\] sel_op\[3\] sel_op\[1\] VGND VGND VPWR VPWR _06804_ sky130_fd_sc_hd__nor3_1
X_17398_ _07869_ _07870_ VGND VGND VPWR VPWR _07871_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_54_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16349_ _03049_ _06612_ _06728_ _06626_ VGND VGND VPWR VPWR _06729_ sky130_fd_sc_hd__o211a_1
XFILLER_0_54_383 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_759 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_770 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_898 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18019_ _08464_ _08545_ _08532_ VGND VGND VPWR VPWR _08547_ sky130_fd_sc_hd__and3_1
XFILLER_0_2_675 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_112_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_83 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09723_ _06460_ _06482_ _05083_ _05072_ VGND VGND VPWR VPWR _06493_ sky130_fd_sc_hd__a31oi_4
X_09654_ _05736_ VGND VGND VPWR VPWR _05747_ sky130_fd_sc_hd__buf_4
X_09585_ _04984_ _03750_ VGND VGND VPWR VPWR _04995_ sky130_fd_sc_hd__and2_4
XTAP_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_135_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10360_ _05017_ _06062_ _00451_ _00452_ VGND VGND VPWR VPWR _00453_ sky130_fd_sc_hd__nand4_2
XFILLER_0_143_591 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10291_ _09240_ _09326_ _09287_ VGND VGND VPWR VPWR _00384_ sky130_fd_sc_hd__o21a_1
X_12030_ _02108_ _02121_ VGND VGND VPWR VPWR _02123_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_103_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13981_ _09172_ _04154_ _00563_ _00358_ VGND VGND VPWR VPWR _04153_ sky130_fd_sc_hd__a22o_1
X_15720_ _05890_ _05983_ VGND VGND VPWR VPWR _06049_ sky130_fd_sc_hd__and2b_1
X_12932_ _01113_ VGND VGND VPWR VPWR _03025_ sky130_fd_sc_hd__buf_2
X_15651_ _09351_ _09311_ _07744_ _02991_ VGND VGND VPWR VPWR _05974_ sky130_fd_sc_hd__a22o_1
XTAP_2320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12863_ _02954_ _02955_ VGND VGND VPWR VPWR _02956_ sky130_fd_sc_hd__and2_1
XTAP_2331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14602_ _00592_ _01112_ _04773_ _04771_ VGND VGND VPWR VPWR _04832_ sky130_fd_sc_hd__a31oi_1
XTAP_2353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18370_ _08835_ _08837_ _08833_ VGND VGND VPWR VPWR _08928_ sky130_fd_sc_hd__a21bo_1
X_11814_ _01906_ _01822_ VGND VGND VPWR VPWR _01907_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_96_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_818 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15582_ _05897_ _05898_ VGND VGND VPWR VPWR _05900_ sky130_fd_sc_hd__nor2_1
XTAP_1630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12794_ _02884_ _02886_ VGND VGND VPWR VPWR _02887_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_28_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17321_ _07654_ _07658_ _07785_ VGND VGND VPWR VPWR _07787_ sky130_fd_sc_hd__or3b_1
X_14533_ _04756_ VGND VGND VPWR VPWR _04757_ sky130_fd_sc_hd__inv_2
XTAP_1663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11745_ _01660_ _01662_ VGND VGND VPWR VPWR _01838_ sky130_fd_sc_hd__xor2_1
XTAP_1674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17252_ _07113_ _06655_ _07489_ _07595_ VGND VGND VPWR VPWR _07712_ sky130_fd_sc_hd__and4_1
XFILLER_0_153_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14464_ _04678_ _04680_ _04533_ _04535_ VGND VGND VPWR VPWR _04682_ sky130_fd_sc_hd__o211a_1
XFILLER_0_43_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11676_ _01760_ _01761_ _01768_ VGND VGND VPWR VPWR _01769_ sky130_fd_sc_hd__nor3b_2
XFILLER_0_71_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16203_ _06567_ _06570_ _00357_ VGND VGND VPWR VPWR _06571_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_37_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13415_ _07047_ VGND VGND VPWR VPWR _03535_ sky130_fd_sc_hd__inv_2
X_10627_ _00553_ _00542_ VGND VGND VPWR VPWR _00720_ sky130_fd_sc_hd__and2b_1
X_17183_ _07634_ _07636_ VGND VGND VPWR VPWR _07637_ sky130_fd_sc_hd__nand2_1
X_14395_ _04598_ _04599_ _04605_ VGND VGND VPWR VPWR _04606_ sky130_fd_sc_hd__and3_1
XFILLER_0_70_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_141_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16134_ _01672_ _03188_ VGND VGND VPWR VPWR _06496_ sky130_fd_sc_hd__or2_1
X_13346_ _03453_ _03458_ VGND VGND VPWR VPWR _03459_ sky130_fd_sc_hd__xnor2_1
X_10558_ _00646_ _00472_ _00649_ _00650_ VGND VGND VPWR VPWR _00651_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_59_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16065_ _06420_ VGND VGND VPWR VPWR _06421_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13277_ _03379_ _03380_ _03381_ VGND VGND VPWR VPWR _03383_ sky130_fd_sc_hd__a21o_1
XFILLER_0_121_252 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10489_ _00535_ _00536_ net186 _00375_ VGND VGND VPWR VPWR _00582_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_59_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15016_ _05262_ _05282_ VGND VGND VPWR VPWR _05284_ sky130_fd_sc_hd__or2_1
X_12228_ _02320_ _02312_ VGND VGND VPWR VPWR _02321_ sky130_fd_sc_hd__and2b_1
XFILLER_0_121_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12159_ _02247_ _02250_ VGND VGND VPWR VPWR _02252_ sky130_fd_sc_hd__and2_1
XFILLER_0_75_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16967_ _07399_ _07400_ VGND VGND VPWR VPWR _07401_ sky130_fd_sc_hd__and2_1
X_18706_ _09235_ VGND VGND VPWR VPWR _00061_ sky130_fd_sc_hd__buf_1
X_15918_ _06260_ _06262_ VGND VGND VPWR VPWR _06263_ sky130_fd_sc_hd__xor2_1
X_16898_ _07212_ _07214_ _07325_ VGND VGND VPWR VPWR _07326_ sky130_fd_sc_hd__o21a_1
XFILLER_0_79_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15849_ _06183_ _06187_ _06188_ VGND VGND VPWR VPWR _06189_ sky130_fd_sc_hd__a21oi_1
X_18637_ _09176_ _09184_ VGND VGND VPWR VPWR _09185_ sky130_fd_sc_hd__and2_1
XFILLER_0_149_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_148_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18568_ salida\[6\] _09114_ _09118_ salida\[38\] _09128_ VGND VGND VPWR VPWR _09135_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_86_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_475 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17519_ _08001_ _08002_ VGND VGND VPWR VPWR _08003_ sky130_fd_sc_hd__xor2_1
XFILLER_0_129_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18499_ _03197_ _06317_ VGND VGND VPWR VPWR _09067_ sky130_fd_sc_hd__nand2_1
XFILLER_0_129_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_712 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_144_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_12_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_12_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_145_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_125_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_578 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09706_ _06288_ _06298_ VGND VGND VPWR VPWR _06309_ sky130_fd_sc_hd__nor2_1
X_09637_ ApproximateM_inst.lob_16.lob2.genblk1\[7\].genblk1.mux.sel VGND VGND VPWR
+ VPWR _05562_ sky130_fd_sc_hd__buf_2
X_09568_ _04777_ _04788_ _04799_ VGND VGND VPWR VPWR _04810_ sky130_fd_sc_hd__nand3_1
XFILLER_0_84_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_423 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09499_ _03399_ VGND VGND VPWR VPWR _04056_ sky130_fd_sc_hd__buf_4
X_11530_ _01185_ _01184_ _01183_ VGND VGND VPWR VPWR _01623_ sky130_fd_sc_hd__a21o_1
XFILLER_0_93_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11461_ _03892_ _00180_ _00130_ _03881_ VGND VGND VPWR VPWR _01554_ sky130_fd_sc_hd__a22o_1
X_13200_ _01504_ _00557_ VGND VGND VPWR VPWR _03301_ sky130_fd_sc_hd__nand2_1
X_10412_ _00497_ _00504_ VGND VGND VPWR VPWR _00505_ sky130_fd_sc_hd__xor2_2
X_14180_ _04369_ _04370_ VGND VGND VPWR VPWR _04371_ sky130_fd_sc_hd__and2_1
X_11392_ _01483_ _01484_ VGND VGND VPWR VPWR _01485_ sky130_fd_sc_hd__nor2_1
XFILLER_0_61_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13131_ _04984_ _05845_ _00613_ _00612_ _00443_ VGND VGND VPWR VPWR _03227_ sky130_fd_sc_hd__a32o_1
X_10343_ _00432_ _00434_ _00433_ VGND VGND VPWR VPWR _00436_ sky130_fd_sc_hd__a21o_1
XFILLER_0_131_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10274_ _00365_ _00366_ VGND VGND VPWR VPWR _00367_ sky130_fd_sc_hd__nor2_2
X_13062_ _03153_ VGND VGND VPWR VPWR _03154_ sky130_fd_sc_hd__clkbuf_4
X_12013_ _02047_ _02048_ _02049_ net328 VGND VGND VPWR VPWR _02106_ sky130_fd_sc_hd__o31ai_2
X_17870_ _08383_ _08384_ VGND VGND VPWR VPWR _08385_ sky130_fd_sc_hd__xnor2_1
X_16821_ _07103_ _07138_ VGND VGND VPWR VPWR _07242_ sky130_fd_sc_hd__and2_1
X_16752_ _07165_ _07166_ VGND VGND VPWR VPWR _07168_ sky130_fd_sc_hd__and2_1
X_13964_ _05834_ _03455_ VGND VGND VPWR VPWR _04135_ sky130_fd_sc_hd__nand2_1
X_15703_ _06028_ _06030_ VGND VGND VPWR VPWR _06031_ sky130_fd_sc_hd__nor2_1
Xmax_cap5 _02383_ VGND VGND VPWR VPWR net323 sky130_fd_sc_hd__clkbuf_1
X_12915_ _09166_ VGND VGND VPWR VPWR _03008_ sky130_fd_sc_hd__buf_2
X_16683_ _02975_ _07089_ _07092_ _06645_ VGND VGND VPWR VPWR _07093_ sky130_fd_sc_hd__a211o_1
X_13895_ _04058_ _04059_ VGND VGND VPWR VPWR _04060_ sky130_fd_sc_hd__xor2_1
X_15634_ _05934_ _05936_ VGND VGND VPWR VPWR _05956_ sky130_fd_sc_hd__or2_1
X_18422_ _01502_ _02891_ _02894_ VGND VGND VPWR VPWR _08985_ sky130_fd_sc_hd__nor3_1
XFILLER_0_0_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12846_ _02920_ _02938_ VGND VGND VPWR VPWR _02939_ sky130_fd_sc_hd__or2_1
XTAP_2150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18353_ _03108_ _07390_ _08845_ _04668_ _07592_ VGND VGND VPWR VPWR _08910_ sky130_fd_sc_hd__a32o_1
XTAP_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15565_ _04076_ _04084_ _03536_ VGND VGND VPWR VPWR _05881_ sky130_fd_sc_hd__mux2_1
X_12777_ _02866_ _02868_ VGND VGND VPWR VPWR _02870_ sky130_fd_sc_hd__nand2_1
XTAP_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17304_ _07767_ _07768_ VGND VGND VPWR VPWR _07769_ sky130_fd_sc_hd__nor2_1
X_14516_ _04735_ _04736_ _04584_ _04704_ VGND VGND VPWR VPWR _04738_ sky130_fd_sc_hd__a211oi_2
XTAP_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18284_ _08833_ _08834_ VGND VGND VPWR VPWR _08835_ sky130_fd_sc_hd__and2_1
X_11728_ _04416_ _00179_ _00129_ _04340_ VGND VGND VPWR VPWR _01821_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_16_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15496_ _03537_ _03913_ _05082_ VGND VGND VPWR VPWR _05806_ sky130_fd_sc_hd__or3_1
XFILLER_0_126_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17235_ _06368_ _06438_ _06425_ VGND VGND VPWR VPWR _07694_ sky130_fd_sc_hd__a21oi_1
X_14447_ _04480_ _04662_ VGND VGND VPWR VPWR _04663_ sky130_fd_sc_hd__xor2_1
XFILLER_0_127_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11659_ _01702_ _01704_ _01750_ VGND VGND VPWR VPWR _01752_ sky130_fd_sc_hd__nor3_1
XFILLER_0_114_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17166_ _07494_ _07588_ _07616_ VGND VGND VPWR VPWR _07618_ sky130_fd_sc_hd__nor3_1
X_14378_ _02059_ _08224_ _04439_ _04437_ VGND VGND VPWR VPWR _04587_ sky130_fd_sc_hd__a31o_1
XFILLER_0_40_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_684 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16117_ _03028_ VGND VGND VPWR VPWR _06477_ sky130_fd_sc_hd__buf_4
X_13329_ _09166_ _09172_ _00218_ _00178_ VGND VGND VPWR VPWR _03440_ sky130_fd_sc_hd__and4_1
X_17097_ _07541_ _07542_ VGND VGND VPWR VPWR _07543_ sky130_fd_sc_hd__and2b_1
XFILLER_0_150_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16048_ _06400_ _06401_ _05557_ VGND VGND VPWR VPWR _06402_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_19_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17999_ _03198_ _05807_ VGND VGND VPWR VPWR _08526_ sky130_fd_sc_hd__nand2_1
XFILLER_0_126_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_414 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09422_ op_code\[1\] VGND VGND VPWR VPWR _03217_ sky130_fd_sc_hd__buf_2
XFILLER_0_19_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_724 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_118_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_94 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_144_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_712 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10961_ _05399_ _05355_ _03804_ _03914_ VGND VGND VPWR VPWR _01054_ sky130_fd_sc_hd__nand4_4
X_12700_ _02764_ _02765_ VGND VGND VPWR VPWR _02793_ sky130_fd_sc_hd__xnor2_1
X_13680_ _03820_ _03822_ _03817_ VGND VGND VPWR VPWR _03824_ sky130_fd_sc_hd__o21ai_1
X_10892_ _00981_ _00984_ VGND VGND VPWR VPWR _00985_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_97_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12631_ _02686_ _02721_ VGND VGND VPWR VPWR _02724_ sky130_fd_sc_hd__nor2_1
XFILLER_0_65_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_823 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15350_ _05452_ _05566_ VGND VGND VPWR VPWR _05647_ sky130_fd_sc_hd__and2b_1
XFILLER_0_31_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12562_ _02611_ _02654_ VGND VGND VPWR VPWR _02655_ sky130_fd_sc_hd__nor2_1
XFILLER_0_93_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14301_ _04501_ _04502_ VGND VGND VPWR VPWR _04503_ sky130_fd_sc_hd__nand2_2
XFILLER_0_81_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11513_ _01550_ _01561_ VGND VGND VPWR VPWR _01606_ sky130_fd_sc_hd__or2_1
X_15281_ _05554_ _05555_ _05570_ VGND VGND VPWR VPWR _05572_ sky130_fd_sc_hd__or3_1
XFILLER_0_25_139 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_109_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12493_ _02585_ _02527_ VGND VGND VPWR VPWR _02586_ sky130_fd_sc_hd__xnor2_1
Xwire133 _04284_ VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__buf_1
XFILLER_0_124_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17020_ _00593_ _07355_ VGND VGND VPWR VPWR _07459_ sky130_fd_sc_hd__nor2_1
X_14232_ _04299_ _04300_ _04312_ VGND VGND VPWR VPWR _04428_ sky130_fd_sc_hd__nor3_1
XFILLER_0_135_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11444_ _04635_ _04362_ _00176_ VGND VGND VPWR VPWR _01537_ sky130_fd_sc_hd__and3_1
XFILLER_0_22_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14163_ _04350_ _04352_ VGND VGND VPWR VPWR _04353_ sky130_fd_sc_hd__and2_2
XFILLER_0_1_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11375_ _01394_ _01413_ _01466_ _01467_ VGND VGND VPWR VPWR _01468_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_132_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13114_ _03465_ _00439_ VGND VGND VPWR VPWR _03209_ sky130_fd_sc_hd__and2_1
X_10326_ _00417_ _00416_ _09342_ _00379_ VGND VGND VPWR VPWR _00419_ sky130_fd_sc_hd__o211ai_2
X_14094_ _04099_ _04132_ _07962_ VGND VGND VPWR VPWR _04277_ sky130_fd_sc_hd__and3_1
X_18971_ clknet_4_5_0_clk _09402_ VGND VGND VPWR VPWR salida\[24\] sky130_fd_sc_hd__dfxtp_1
XTAP_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17922_ _06680_ _08441_ VGND VGND VPWR VPWR _08443_ sky130_fd_sc_hd__nor2_1
X_13045_ _01220_ _03136_ _03040_ VGND VGND VPWR VPWR _03137_ sky130_fd_sc_hd__o21a_1
X_10257_ _00348_ _00337_ _00338_ VGND VGND VPWR VPWR _00350_ sky130_fd_sc_hd__nand3_1
XFILLER_0_147_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10188_ _00278_ _00279_ _00280_ VGND VGND VPWR VPWR _00281_ sky130_fd_sc_hd__nand3_1
X_17853_ _08283_ _08284_ _08282_ VGND VGND VPWR VPWR _08367_ sky130_fd_sc_hd__o21ai_1
X_16804_ _07215_ _07223_ VGND VGND VPWR VPWR _07224_ sky130_fd_sc_hd__xor2_1
X_17784_ _08257_ _08258_ _08291_ VGND VGND VPWR VPWR _08292_ sky130_fd_sc_hd__a21oi_1
X_14996_ _05260_ _05261_ VGND VGND VPWR VPWR _05262_ sky130_fd_sc_hd__and2_1
X_13947_ _04109_ _04115_ VGND VGND VPWR VPWR _04116_ sky130_fd_sc_hd__xnor2_1
X_16735_ _07139_ _07148_ VGND VGND VPWR VPWR _07149_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_72_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_58 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16666_ _02800_ _07073_ _04238_ VGND VGND VPWR VPWR _07074_ sky130_fd_sc_hd__a21oi_1
X_13878_ _04025_ _04026_ _04040_ VGND VGND VPWR VPWR _04041_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_88_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15617_ _05861_ net118 _05937_ VGND VGND VPWR VPWR _05938_ sky130_fd_sc_hd__o21bai_1
X_18405_ _08912_ _08915_ VGND VGND VPWR VPWR _08966_ sky130_fd_sc_hd__nand2_1
X_12829_ _02903_ _02904_ VGND VGND VPWR VPWR _02922_ sky130_fd_sc_hd__and2_2
X_16597_ _00494_ _02983_ _06487_ _06485_ VGND VGND VPWR VPWR _06999_ sky130_fd_sc_hd__or4_2
XFILLER_0_146_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_754 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15548_ _05757_ _05861_ _05862_ VGND VGND VPWR VPWR _05863_ sky130_fd_sc_hd__nor3_1
XFILLER_0_56_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18336_ _03206_ _08873_ _08874_ _08891_ VGND VGND VPWR VPWR _08892_ sky130_fd_sc_hd__o31ai_1
XTAP_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_139_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18267_ _08815_ _08816_ _06508_ VGND VGND VPWR VPWR _08817_ sky130_fd_sc_hd__o21a_1
XFILLER_0_126_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15479_ _05700_ _05702_ _05787_ VGND VGND VPWR VPWR _05788_ sky130_fd_sc_hd__o21ba_2
XFILLER_0_72_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_826 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_612 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17218_ _07673_ _07674_ _06649_ VGND VGND VPWR VPWR _07675_ sky130_fd_sc_hd__and3b_2
XFILLER_0_71_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18198_ _08586_ _08668_ VGND VGND VPWR VPWR _08742_ sky130_fd_sc_hd__or2b_1
XFILLER_0_114_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17149_ _06657_ net145 VGND VGND VPWR VPWR _07599_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09971_ cla_inst.in2\[30\] VGND VGND VPWR VPWR _09166_ sky130_fd_sc_hd__buf_2
XFILLER_0_79_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_367 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_137_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_743 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_153_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_117_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_826 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_132_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_114_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11160_ _00203_ _00134_ VGND VGND VPWR VPWR _01253_ sky130_fd_sc_hd__nand2_1
XFILLER_0_101_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10111_ _00203_ VGND VGND VPWR VPWR _00204_ sky130_fd_sc_hd__clkbuf_4
X_11091_ _05464_ _03837_ _04056_ _05508_ VGND VGND VPWR VPWR _01184_ sky130_fd_sc_hd__a22o_1
XFILLER_0_101_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10042_ _00126_ VGND VGND VPWR VPWR _00135_ sky130_fd_sc_hd__inv_2
X_14850_ _03651_ _03662_ _07755_ _08169_ VGND VGND VPWR VPWR _05102_ sky130_fd_sc_hd__nand4_2
Xhold85 op_code\[0\] VGND VGND VPWR VPWR net248 sky130_fd_sc_hd__buf_1
X_13801_ _04548_ _08169_ _03953_ _03954_ VGND VGND VPWR VPWR _03956_ sky130_fd_sc_hd__o2bb2a_1
Xhold96 net108 VGND VGND VPWR VPWR net259 sky130_fd_sc_hd__dlygate4sd3_1
X_14781_ _05025_ _05026_ VGND VGND VPWR VPWR _05027_ sky130_fd_sc_hd__nor2_1
X_11993_ _04351_ _04373_ _07548_ _07581_ VGND VGND VPWR VPWR _02086_ sky130_fd_sc_hd__and4_1
XFILLER_0_97_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16520_ _06913_ _06914_ _04247_ VGND VGND VPWR VPWR _06915_ sky130_fd_sc_hd__mux2_2
X_13732_ _03836_ _03715_ _03879_ _03880_ VGND VGND VPWR VPWR _03882_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_97_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10944_ _01029_ _01030_ _01035_ VGND VGND VPWR VPWR _01037_ sky130_fd_sc_hd__nand3_1
XFILLER_0_98_687 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16451_ _06781_ _06782_ _06780_ VGND VGND VPWR VPWR _06840_ sky130_fd_sc_hd__a21bo_1
X_13663_ _03802_ _03803_ _03789_ VGND VGND VPWR VPWR _03806_ sky130_fd_sc_hd__a21o_1
X_10875_ _04001_ _00165_ _00921_ _00920_ VGND VGND VPWR VPWR _00968_ sky130_fd_sc_hd__a31o_1
XFILLER_0_128_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15402_ _05575_ _05576_ _05587_ VGND VGND VPWR VPWR _05705_ sky130_fd_sc_hd__and3_1
X_12614_ _02701_ _02704_ _02705_ _02706_ VGND VGND VPWR VPWR _02707_ sky130_fd_sc_hd__a211oi_1
X_16382_ _06764_ VGND VGND VPWR VPWR _06766_ sky130_fd_sc_hd__clkbuf_4
X_13594_ _03518_ _03521_ _03730_ VGND VGND VPWR VPWR _03731_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_54_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_109_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18121_ _08654_ _08657_ VGND VGND VPWR VPWR _08658_ sky130_fd_sc_hd__xnor2_1
X_15333_ _05574_ _05592_ VGND VGND VPWR VPWR _05629_ sky130_fd_sc_hd__or2_1
XFILLER_0_108_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12545_ _07036_ _07973_ _00871_ _09179_ VGND VGND VPWR VPWR _02638_ sky130_fd_sc_hd__nand4_2
XFILLER_0_108_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18052_ _08497_ _08530_ _08581_ VGND VGND VPWR VPWR _08584_ sky130_fd_sc_hd__and3_1
X_15264_ _05339_ _05472_ VGND VGND VPWR VPWR _05554_ sky130_fd_sc_hd__and2b_1
X_12476_ _02510_ _02512_ VGND VGND VPWR VPWR _02569_ sky130_fd_sc_hd__xnor2_1
X_17003_ _07438_ _07440_ VGND VGND VPWR VPWR _07441_ sky130_fd_sc_hd__nand2_1
X_14215_ _02963_ _04404_ _04409_ VGND VGND VPWR VPWR _04410_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_124_678 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11427_ _03509_ VGND VGND VPWR VPWR _01520_ sky130_fd_sc_hd__buf_4
XANTENNA_5 _00206_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15195_ _05461_ _05462_ _05477_ VGND VGND VPWR VPWR _05479_ sky130_fd_sc_hd__or3_1
XFILLER_0_22_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14146_ _04332_ _04333_ VGND VGND VPWR VPWR _04334_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_6_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11358_ _01337_ _01377_ _01440_ _01441_ VGND VGND VPWR VPWR _01451_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_22_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10309_ _00204_ _00166_ _00260_ VGND VGND VPWR VPWR _00402_ sky130_fd_sc_hd__and3_1
XTAP_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18954_ clknet_4_1_0_clk _09415_ VGND VGND VPWR VPWR salida\[7\] sky130_fd_sc_hd__dfxtp_1
X_14077_ _03576_ _03579_ _03060_ VGND VGND VPWR VPWR _04258_ sky130_fd_sc_hd__mux2_1
X_11289_ _01279_ net140 _00794_ _01381_ VGND VGND VPWR VPWR _01382_ sky130_fd_sc_hd__o211ai_4
XTAP_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13028_ _03120_ VGND VGND VPWR VPWR _03121_ sky130_fd_sc_hd__buf_4
X_17905_ _02173_ _08423_ VGND VGND VPWR VPWR _08424_ sky130_fd_sc_hd__nor2_1
X_18885_ clknet_4_13_0_clk _00039_ VGND VGND VPWR VPWR ApproximateM_inst.lob_16.lob1.genblk1\[3\].genblk1.mux.sel
+ sky130_fd_sc_hd__dfxtp_1
X_17836_ _08294_ _08312_ VGND VGND VPWR VPWR _08348_ sky130_fd_sc_hd__nor2_1
XFILLER_0_89_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xrebuffer17 _01858_ VGND VGND VPWR VPWR net180 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer28 net337 VGND VGND VPWR VPWR net191 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17767_ _08271_ _08272_ VGND VGND VPWR VPWR _08273_ sky130_fd_sc_hd__nand2_1
Xrebuffer39 _04882_ VGND VGND VPWR VPWR net202 sky130_fd_sc_hd__clkbuf_1
X_14979_ _05240_ _05242_ VGND VGND VPWR VPWR _05243_ sky130_fd_sc_hd__xor2_2
X_16718_ _07035_ VGND VGND VPWR VPWR _07130_ sky130_fd_sc_hd__clkbuf_4
X_17698_ _08074_ _08076_ _08197_ VGND VGND VPWR VPWR _08198_ sky130_fd_sc_hd__o21a_1
XFILLER_0_76_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16649_ _07053_ _07054_ VGND VGND VPWR VPWR _07055_ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18319_ _08840_ _08841_ _08872_ VGND VGND VPWR VPWR _08873_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_5_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_114_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_144 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_142_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_130_615 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_142_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09954_ _08681_ _08973_ _08984_ _08995_ VGND VGND VPWR VPWR _09005_ sky130_fd_sc_hd__nand4_4
XFILLER_0_110_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09885_ _08148_ _08246_ VGND VGND VPWR VPWR _08256_ sky130_fd_sc_hd__xor2_4
XTAP_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_137_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10660_ _00750_ _00751_ _00585_ _00599_ VGND VGND VPWR VPWR _00753_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_82_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_153_707 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10591_ _00682_ _00683_ VGND VGND VPWR VPWR _00684_ sky130_fd_sc_hd__or2_1
XFILLER_0_146_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_152_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_340 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12330_ _00992_ _05638_ _00196_ _00871_ VGND VGND VPWR VPWR _02423_ sky130_fd_sc_hd__and4_1
XFILLER_0_51_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12261_ _07973_ _04220_ _00774_ _07984_ VGND VGND VPWR VPWR _02354_ sky130_fd_sc_hd__a22o_1
XFILLER_0_105_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14000_ _04014_ _04013_ VGND VGND VPWR VPWR _04174_ sky130_fd_sc_hd__or2b_1
X_11212_ _01293_ _01294_ _01303_ VGND VGND VPWR VPWR _01305_ sky130_fd_sc_hd__nand3_1
X_12192_ _02195_ _02198_ _02284_ VGND VGND VPWR VPWR _02285_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_120_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11143_ _01204_ _01233_ _01234_ _01235_ VGND VGND VPWR VPWR _01236_ sky130_fd_sc_hd__or4_4
Xoutput75 net75 VGND VGND VPWR VPWR leds[3] sky130_fd_sc_hd__buf_2
Xoutput86 net86 VGND VGND VPWR VPWR o_wb_data[12] sky130_fd_sc_hd__clkbuf_4
Xoutput97 net97 VGND VGND VPWR VPWR o_wb_data[22] sky130_fd_sc_hd__clkbuf_4
X_11074_ _03728_ _00218_ _01153_ _01152_ VGND VGND VPWR VPWR _01167_ sky130_fd_sc_hd__a31o_1
X_15951_ _06287_ VGND VGND VPWR VPWR _06297_ sky130_fd_sc_hd__inv_2
X_14902_ _05141_ _05142_ _05157_ VGND VGND VPWR VPWR _05160_ sky130_fd_sc_hd__nor3_1
X_10025_ _00105_ _00117_ VGND VGND VPWR VPWR _00118_ sky130_fd_sc_hd__and2_1
X_18670_ _09209_ _09210_ VGND VGND VPWR VPWR _09211_ sky130_fd_sc_hd__and2_1
X_15882_ _06221_ _06223_ VGND VGND VPWR VPWR _06225_ sky130_fd_sc_hd__xnor2_1
X_17621_ _08001_ _08002_ _08004_ VGND VGND VPWR VPWR _08114_ sky130_fd_sc_hd__a21o_1
X_14833_ _05082_ _05084_ _03081_ VGND VGND VPWR VPWR _05085_ sky130_fd_sc_hd__mux2_1
X_14764_ _05001_ _05008_ VGND VGND VPWR VPWR _05009_ sky130_fd_sc_hd__or2_1
X_17552_ _06421_ _08030_ _08031_ _08033_ _08038_ VGND VGND VPWR VPWR _08040_ sky130_fd_sc_hd__a311o_1
X_11976_ _02056_ _02066_ VGND VGND VPWR VPWR _02069_ sky130_fd_sc_hd__xor2_1
X_13715_ _09353_ _00398_ _03705_ _03704_ VGND VGND VPWR VPWR _03863_ sky130_fd_sc_hd__a31o_1
X_16503_ _06888_ _06896_ VGND VGND VPWR VPWR _06897_ sky130_fd_sc_hd__xor2_2
X_10927_ _00980_ _01018_ _01019_ VGND VGND VPWR VPWR _01020_ sky130_fd_sc_hd__nor3_2
X_17483_ _07955_ _07963_ VGND VGND VPWR VPWR _07964_ sky130_fd_sc_hd__xnor2_1
X_14695_ _04932_ _04933_ VGND VGND VPWR VPWR _04934_ sky130_fd_sc_hd__nor2_2
X_13646_ _03784_ _03785_ _03606_ net324 VGND VGND VPWR VPWR _03787_ sky130_fd_sc_hd__a211oi_4
X_16434_ _06769_ _06821_ VGND VGND VPWR VPWR _06822_ sky130_fd_sc_hd__or2_1
X_10858_ _04493_ _04416_ _03388_ _00949_ VGND VGND VPWR VPWR _00951_ sky130_fd_sc_hd__and4_1
XFILLER_0_54_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16365_ _04241_ _06739_ _06746_ _03117_ VGND VGND VPWR VPWR _06747_ sky130_fd_sc_hd__a211o_1
X_13577_ _03700_ _03711_ VGND VGND VPWR VPWR _03712_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10789_ _00877_ _00881_ VGND VGND VPWR VPWR _00882_ sky130_fd_sc_hd__nand2_1
XPHY_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15316_ _05607_ _05610_ VGND VGND VPWR VPWR _05611_ sky130_fd_sc_hd__xor2_1
XFILLER_0_5_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18104_ _07604_ _07623_ _08638_ VGND VGND VPWR VPWR _08640_ sky130_fd_sc_hd__a21o_1
XFILLER_0_143_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12528_ _02540_ _02620_ VGND VGND VPWR VPWR _02621_ sky130_fd_sc_hd__and2_1
XFILLER_0_54_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16296_ _00494_ _06509_ _06427_ VGND VGND VPWR VPWR _06672_ sky130_fd_sc_hd__a21o_1
XFILLER_0_140_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15247_ _05532_ _05533_ VGND VGND VPWR VPWR _05535_ sky130_fd_sc_hd__and2_1
XFILLER_0_2_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_124_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18035_ _08563_ _08564_ VGND VGND VPWR VPWR _08565_ sky130_fd_sc_hd__xor2_1
XFILLER_0_1_301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12459_ _07243_ _00145_ _00129_ _07221_ VGND VGND VPWR VPWR _02552_ sky130_fd_sc_hd__a22o_1
X_15178_ _05364_ VGND VGND VPWR VPWR _05460_ sky130_fd_sc_hd__inv_2
XFILLER_0_111_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14129_ _04123_ _04145_ _04313_ _04314_ VGND VGND VPWR VPWR _04315_ sky130_fd_sc_hd__o211a_2
X_18937_ clknet_4_3_0_clk _00091_ VGND VGND VPWR VPWR cla_inst.in2\[23\] sky130_fd_sc_hd__dfxtp_1
X_09670_ _04591_ VGND VGND VPWR VPWR _05921_ sky130_fd_sc_hd__buf_6
X_18868_ clknet_4_5_0_clk _00034_ VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__dfxtp_1
X_17819_ _03041_ _06511_ _02985_ VGND VGND VPWR VPWR _08330_ sky130_fd_sc_hd__and3b_1
X_18799_ _09308_ VGND VGND VPWR VPWR _00090_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_135_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_128_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_142_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09937_ _08800_ _08811_ VGND VGND VPWR VPWR _08822_ sky130_fd_sc_hd__xor2_1
XTAP_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09868_ _08039_ _06613_ _08049_ _06019_ VGND VGND VPWR VPWR _08071_ sky130_fd_sc_hd__a22o_1
XFILLER_0_99_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09799_ _07210_ _07297_ _07308_ VGND VGND VPWR VPWR _07319_ sky130_fd_sc_hd__nand3_4
XTAP_2502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11830_ _06591_ _00774_ _00909_ _00806_ VGND VGND VPWR VPWR _01923_ sky130_fd_sc_hd__a22o_1
XTAP_2524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11761_ _01657_ _01656_ VGND VGND VPWR VPWR _01854_ sky130_fd_sc_hd__and2b_1
XTAP_1834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13500_ _03625_ _03626_ VGND VGND VPWR VPWR _03627_ sky130_fd_sc_hd__nor2_1
XFILLER_0_67_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10712_ _00803_ _00804_ VGND VGND VPWR VPWR _00805_ sky130_fd_sc_hd__xor2_2
XFILLER_0_49_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14480_ _04628_ _04629_ _04674_ _04675_ VGND VGND VPWR VPWR _04698_ sky130_fd_sc_hd__and4bb_1
XTAP_1878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11692_ _01742_ _01753_ VGND VGND VPWR VPWR _01785_ sky130_fd_sc_hd__and2_1
XTAP_1889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_392 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13431_ _03105_ _03110_ _03048_ VGND VGND VPWR VPWR _03552_ sky130_fd_sc_hd__mux2_1
X_10643_ _00733_ _00734_ _00721_ _00722_ VGND VGND VPWR VPWR _00736_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_153_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16150_ _01113_ _06509_ _09354_ VGND VGND VPWR VPWR _06513_ sky130_fd_sc_hd__a21o_1
XFILLER_0_23_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13362_ _01504_ _00716_ VGND VGND VPWR VPWR _03477_ sky130_fd_sc_hd__nand2_1
XFILLER_0_36_598 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10574_ _06711_ _07384_ _00478_ _00319_ _08158_ VGND VGND VPWR VPWR _00667_ sky130_fd_sc_hd__a32o_1
Xrebuffer8 _03781_ VGND VGND VPWR VPWR net171 sky130_fd_sc_hd__clkbuf_1
X_15101_ _01745_ _03067_ VGND VGND VPWR VPWR _05376_ sky130_fd_sc_hd__nand2_1
XFILLER_0_140_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12313_ _02402_ _02404_ VGND VGND VPWR VPWR _02406_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_106_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16081_ _00558_ _06437_ VGND VGND VPWR VPWR _06438_ sky130_fd_sc_hd__and2_1
X_13293_ _04558_ _07962_ _03397_ _03398_ VGND VGND VPWR VPWR _03401_ sky130_fd_sc_hd__a22o_1
X_15032_ _05299_ _05300_ VGND VGND VPWR VPWR _05302_ sky130_fd_sc_hd__or2_1
X_12244_ _02244_ VGND VGND VPWR VPWR _02337_ sky130_fd_sc_hd__inv_2
XFILLER_0_31_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12175_ _02265_ _02267_ VGND VGND VPWR VPWR _02268_ sky130_fd_sc_hd__or2_4
X_11126_ _01132_ _01205_ _01216_ VGND VGND VPWR VPWR _01219_ sky130_fd_sc_hd__a21oi_2
X_16983_ _07416_ _07418_ VGND VGND VPWR VPWR _07419_ sky130_fd_sc_hd__nand2_1
X_18722_ _09247_ VGND VGND VPWR VPWR _00066_ sky130_fd_sc_hd__clkbuf_1
X_11057_ _01037_ _01036_ _01028_ VGND VGND VPWR VPWR _01150_ sky130_fd_sc_hd__a21o_1
X_15934_ _06278_ _06279_ VGND VGND VPWR VPWR _06280_ sky130_fd_sc_hd__nand2_1
X_10008_ _09350_ VGND VGND VPWR VPWR _09351_ sky130_fd_sc_hd__clkbuf_4
X_18653_ _09198_ VGND VGND VPWR VPWR _00040_ sky130_fd_sc_hd__buf_1
X_15865_ _06037_ _06163_ _02992_ _05652_ VGND VGND VPWR VPWR _06206_ sky130_fd_sc_hd__o211a_1
X_17604_ _08087_ _08095_ VGND VGND VPWR VPWR _08096_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_99_771 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14816_ _05063_ _05064_ _04967_ _04928_ VGND VGND VPWR VPWR _05066_ sky130_fd_sc_hd__a211o_1
X_18584_ net293 _09140_ _09147_ _09144_ VGND VGND VPWR VPWR _00015_ sky130_fd_sc_hd__o211a_1
X_15796_ _06086_ _06130_ VGND VGND VPWR VPWR _06132_ sky130_fd_sc_hd__nand2_1
XFILLER_0_148_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17535_ _02846_ _02847_ _04238_ VGND VGND VPWR VPWR _08021_ sky130_fd_sc_hd__a21oi_1
X_14747_ _04845_ _04988_ _04986_ _04987_ VGND VGND VPWR VPWR _04990_ sky130_fd_sc_hd__o211ai_4
X_11959_ _02042_ _02050_ _02027_ _02051_ VGND VGND VPWR VPWR _02052_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_129_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14678_ _04906_ _04914_ VGND VGND VPWR VPWR _04915_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_80_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17466_ _07943_ _07944_ VGND VGND VPWR VPWR _07945_ sky130_fd_sc_hd__xor2_1
XFILLER_0_13_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13629_ _03761_ _03762_ _03767_ VGND VGND VPWR VPWR _03768_ sky130_fd_sc_hd__nand3_1
X_16417_ _04340_ _04362_ VGND VGND VPWR VPWR _06803_ sky130_fd_sc_hd__or2_1
XFILLER_0_117_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17397_ _06875_ _07314_ VGND VGND VPWR VPWR _07870_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16348_ _02982_ _06619_ VGND VGND VPWR VPWR _06728_ sky130_fd_sc_hd__or2_1
XFILLER_0_54_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_152_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16279_ _06652_ VGND VGND VPWR VPWR _06653_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_120_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18018_ _08464_ _08532_ _08545_ VGND VGND VPWR VPWR _08546_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_23_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_687 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09722_ _06471_ VGND VGND VPWR VPWR _06482_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_129_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09653_ _05682_ VGND VGND VPWR VPWR _05736_ sky130_fd_sc_hd__buf_4
XFILLER_0_96_218 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09584_ _03717_ VGND VGND VPWR VPWR _04984_ sky130_fd_sc_hd__buf_6
XFILLER_0_89_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_708 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10290_ _07624_ _00240_ _00382_ VGND VGND VPWR VPWR _00383_ sky130_fd_sc_hd__a21o_1
XFILLER_0_131_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13980_ _09166_ _09172_ _04154_ _00563_ VGND VGND VPWR VPWR _04152_ sky130_fd_sc_hd__and4_1
X_12931_ _03023_ VGND VGND VPWR VPWR _03024_ sky130_fd_sc_hd__buf_2
X_15650_ _03015_ _03142_ _05884_ _05883_ VGND VGND VPWR VPWR _05973_ sky130_fd_sc_hd__a31o_1
X_12862_ _00904_ _02953_ _02952_ _02945_ VGND VGND VPWR VPWR _02955_ sky130_fd_sc_hd__o211ai_1
XTAP_2310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_730 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14601_ _04822_ _04824_ _04830_ VGND VGND VPWR VPWR _09356_ sky130_fd_sc_hd__a21bo_1
X_11813_ _01823_ _01821_ VGND VGND VPWR VPWR _01906_ sky130_fd_sc_hd__or2_1
X_15581_ _09351_ _07744_ _05896_ VGND VGND VPWR VPWR _05898_ sky130_fd_sc_hd__and3_1
XTAP_2354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12793_ _02873_ _02877_ _02885_ VGND VGND VPWR VPWR _02886_ sky130_fd_sc_hd__a21oi_1
XTAP_2365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14532_ _04741_ _04742_ _04753_ VGND VGND VPWR VPWR _04756_ sky130_fd_sc_hd__nand3_2
XTAP_1653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17320_ _07654_ _07658_ _07785_ VGND VGND VPWR VPWR _07786_ sky130_fd_sc_hd__o21ba_1
XTAP_1664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11744_ _01835_ _01832_ VGND VGND VPWR VPWR _01837_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_95_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14463_ _04533_ _04535_ _04678_ _04680_ VGND VGND VPWR VPWR _04681_ sky130_fd_sc_hd__a211oi_2
X_17251_ _07707_ _07709_ VGND VGND VPWR VPWR _07710_ sky130_fd_sc_hd__nand2_1
X_11675_ _01766_ _01767_ VGND VGND VPWR VPWR _01768_ sky130_fd_sc_hd__xnor2_1
X_16202_ _06532_ _06568_ VGND VGND VPWR VPWR _06570_ sky130_fd_sc_hd__nor2_2
X_13414_ _02977_ _00494_ _03533_ VGND VGND VPWR VPWR _03534_ sky130_fd_sc_hd__or3_2
XFILLER_0_153_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10626_ _00543_ _00552_ VGND VGND VPWR VPWR _00719_ sky130_fd_sc_hd__and2_1
X_17182_ _07630_ _07332_ _07632_ _07633_ VGND VGND VPWR VPWR _07636_ sky130_fd_sc_hd__o22ai_1
X_14394_ _04603_ _04604_ VGND VGND VPWR VPWR _04605_ sky130_fd_sc_hd__and2_1
XFILLER_0_52_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16133_ _01863_ _03186_ VGND VGND VPWR VPWR _06495_ sky130_fd_sc_hd__or2_1
XFILLER_0_24_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13345_ _02972_ _03456_ _03457_ VGND VGND VPWR VPWR _03458_ sky130_fd_sc_hd__and3_1
X_10557_ _05834_ _07123_ _00647_ _00648_ VGND VGND VPWR VPWR _00650_ sky130_fd_sc_hd__a22o_1
XFILLER_0_134_592 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16064_ _02965_ _06418_ _06419_ VGND VGND VPWR VPWR _06420_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_11_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13276_ _03379_ _03380_ _03381_ VGND VGND VPWR VPWR _03382_ sky130_fd_sc_hd__nand3_1
XFILLER_0_110_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10488_ _00578_ _00579_ _00396_ _00538_ VGND VGND VPWR VPWR _00581_ sky130_fd_sc_hd__o211a_1
X_15015_ _05262_ _05282_ VGND VGND VPWR VPWR _05283_ sky130_fd_sc_hd__nand2_1
XFILLER_0_121_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12227_ _02313_ _02319_ VGND VGND VPWR VPWR _02320_ sky130_fd_sc_hd__xnor2_1
X_12158_ _02247_ _02250_ VGND VGND VPWR VPWR _02251_ sky130_fd_sc_hd__xor2_1
X_11109_ _01051_ _01052_ _01039_ _01050_ VGND VGND VPWR VPWR _01202_ sky130_fd_sc_hd__a211oi_1
X_12089_ _02178_ _02181_ VGND VGND VPWR VPWR _02182_ sky130_fd_sc_hd__or2_1
X_16966_ _06766_ _07106_ _07398_ VGND VGND VPWR VPWR _07400_ sky130_fd_sc_hd__o21ai_1
X_18705_ _09209_ _09234_ VGND VGND VPWR VPWR _09235_ sky130_fd_sc_hd__and2_1
X_15917_ _06219_ _06261_ VGND VGND VPWR VPWR _06262_ sky130_fd_sc_hd__nand2_1
X_16897_ _07215_ _07223_ VGND VGND VPWR VPWR _07325_ sky130_fd_sc_hd__or2_1
X_18636_ net35 _03029_ _09183_ VGND VGND VPWR VPWR _09184_ sky130_fd_sc_hd__mux2_1
X_15848_ _06183_ _06187_ _03202_ VGND VGND VPWR VPWR _06188_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_59_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18567_ net252 _09098_ _09134_ _09126_ VGND VGND VPWR VPWR _00009_ sky130_fd_sc_hd__o211a_1
XFILLER_0_24_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15779_ _06111_ _06112_ VGND VGND VPWR VPWR _06113_ sky130_fd_sc_hd__nor2_1
XFILLER_0_148_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_129_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17518_ _07860_ _07865_ _07862_ VGND VGND VPWR VPWR _08002_ sky130_fd_sc_hd__a21bo_1
X_18498_ _06413_ _07274_ _09065_ _06720_ VGND VGND VPWR VPWR _09066_ sky130_fd_sc_hd__o211a_1
XFILLER_0_74_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17449_ _06426_ _06441_ _07916_ _07924_ _07926_ VGND VGND VPWR VPWR _07927_ sky130_fd_sc_hd__o311a_1
XFILLER_0_62_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09705_ _04088_ _03892_ _04395_ _04886_ VGND VGND VPWR VPWR _06298_ sky130_fd_sc_hd__and4_1
XFILLER_0_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09636_ _05442_ _05540_ VGND VGND VPWR VPWR _05551_ sky130_fd_sc_hd__xnor2_2
X_09567_ _03509_ _03914_ _03476_ _03531_ VGND VGND VPWR VPWR _04799_ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09498_ _03837_ VGND VGND VPWR VPWR _04045_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_81_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11460_ _04088_ _04121_ _00180_ _00130_ VGND VGND VPWR VPWR _01553_ sky130_fd_sc_hd__nand4_1
XFILLER_0_18_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10411_ _00501_ _00503_ VGND VGND VPWR VPWR _00504_ sky130_fd_sc_hd__xnor2_2
X_11391_ _01473_ _01482_ VGND VGND VPWR VPWR _01484_ sky130_fd_sc_hd__nor2_1
XFILLER_0_61_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13130_ _00625_ _00626_ VGND VGND VPWR VPWR _03226_ sky130_fd_sc_hd__nand2_1
X_10342_ _00432_ _00433_ _00434_ VGND VGND VPWR VPWR _00435_ sky130_fd_sc_hd__nand3_1
XFILLER_0_104_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13061_ _00665_ VGND VGND VPWR VPWR _03153_ sky130_fd_sc_hd__clkbuf_4
X_10273_ _00355_ _00356_ _00364_ VGND VGND VPWR VPWR _00366_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_29_18 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12012_ _02103_ _02104_ VGND VGND VPWR VPWR _02105_ sky130_fd_sc_hd__and2b_1
X_16820_ _07103_ _07138_ VGND VGND VPWR VPWR _07241_ sky130_fd_sc_hd__or2_1
X_16751_ _00214_ _06673_ _02533_ VGND VGND VPWR VPWR _07166_ sky130_fd_sc_hd__or3b_1
X_13963_ _04131_ _04133_ VGND VGND VPWR VPWR _04134_ sky130_fd_sc_hd__nor2_1
X_15702_ _06024_ _06027_ VGND VGND VPWR VPWR _06030_ sky130_fd_sc_hd__nor2_1
Xmax_cap6 _03753_ VGND VGND VPWR VPWR net324 sky130_fd_sc_hd__buf_1
X_12914_ _03006_ VGND VGND VPWR VPWR _03007_ sky130_fd_sc_hd__buf_2
X_13894_ net119 _03893_ VGND VGND VPWR VPWR _04059_ sky130_fd_sc_hd__nor2_2
X_16682_ _03921_ _07090_ VGND VGND VPWR VPWR _07092_ sky130_fd_sc_hd__nor2_1
XFILLER_0_69_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18421_ _08981_ _08982_ VGND VGND VPWR VPWR _08983_ sky130_fd_sc_hd__xnor2_1
X_15633_ _05924_ VGND VGND VPWR VPWR _05955_ sky130_fd_sc_hd__inv_2
X_12845_ _02936_ _02937_ VGND VGND VPWR VPWR _02938_ sky130_fd_sc_hd__or2b_1
XTAP_2140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18352_ _08906_ _08907_ VGND VGND VPWR VPWR _08909_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_424 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12776_ _02866_ _02868_ VGND VGND VPWR VPWR _02869_ sky130_fd_sc_hd__or2_1
XTAP_2195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15564_ _05804_ _05623_ _05807_ _03125_ _05880_ VGND VGND VPWR VPWR _09367_ sky130_fd_sc_hd__a221o_1
XTAP_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17303_ _07735_ _07765_ VGND VGND VPWR VPWR _07768_ sky130_fd_sc_hd__and2_1
X_14515_ _04584_ _04704_ _04735_ _04736_ VGND VGND VPWR VPWR _04737_ sky130_fd_sc_hd__o211a_4
X_11727_ _01816_ _01819_ VGND VGND VPWR VPWR _01820_ sky130_fd_sc_hd__or2b_1
XFILLER_0_126_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18283_ _03143_ _08428_ _01417_ VGND VGND VPWR VPWR _08834_ sky130_fd_sc_hd__or3b_1
X_15495_ _05084_ _05088_ _03081_ VGND VGND VPWR VPWR _05805_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17234_ _06484_ _07688_ _07689_ _07692_ _06462_ VGND VGND VPWR VPWR _07693_ sky130_fd_sc_hd__a311o_1
XFILLER_0_25_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14446_ _04653_ _04661_ VGND VGND VPWR VPWR _04662_ sky130_fd_sc_hd__xnor2_1
X_11658_ _01702_ _01704_ _01750_ VGND VGND VPWR VPWR _01751_ sky130_fd_sc_hd__o21a_1
XFILLER_0_126_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10609_ _00183_ VGND VGND VPWR VPWR _00702_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_25_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14377_ _04451_ _04452_ VGND VGND VPWR VPWR _04586_ sky130_fd_sc_hd__or2_1
XFILLER_0_4_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17165_ _07494_ _07588_ _07616_ VGND VGND VPWR VPWR _07617_ sky130_fd_sc_hd__o21a_1
XFILLER_0_142_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11589_ _05682_ _08409_ _01578_ _01577_ VGND VGND VPWR VPWR _01682_ sky130_fd_sc_hd__a31o_1
XFILLER_0_10_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13328_ _03005_ _01264_ VGND VGND VPWR VPWR _03439_ sky130_fd_sc_hd__nand2_1
XFILLER_0_51_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16116_ _03050_ _02607_ _03170_ _06470_ _06475_ VGND VGND VPWR VPWR _06476_ sky130_fd_sc_hd__o311a_1
X_17096_ _07539_ _07426_ _07540_ VGND VGND VPWR VPWR _07542_ sky130_fd_sc_hd__or3b_1
XFILLER_0_40_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_150_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13259_ _03202_ _03362_ _03363_ VGND VGND VPWR VPWR _03364_ sky130_fd_sc_hd__and3_1
X_16047_ _01359_ _03056_ VGND VGND VPWR VPWR _06401_ sky130_fd_sc_hd__or2_1
XFILLER_0_110_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17998_ _06915_ _08141_ _08524_ _06721_ VGND VGND VPWR VPWR _08525_ sky130_fd_sc_hd__o211a_1
X_16949_ _07333_ _07334_ VGND VGND VPWR VPWR _07381_ sky130_fd_sc_hd__or2b_1
XFILLER_0_79_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09421_ _03195_ VGND VGND VPWR VPWR _03206_ sky130_fd_sc_hd__buf_4
XFILLER_0_126_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18619_ net269 _09157_ _09170_ _09162_ VGND VGND VPWR VPWR _00030_ sky130_fd_sc_hd__o211a_1
XFILLER_0_149_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_251 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_142_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_632 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_162 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_132_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10960_ _01039_ _01050_ _01051_ _01052_ VGND VGND VPWR VPWR _01053_ sky130_fd_sc_hd__o211a_1
XFILLER_0_98_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09619_ _05355_ VGND VGND VPWR VPWR _05366_ sky130_fd_sc_hd__buf_6
X_10891_ _00982_ _00983_ VGND VGND VPWR VPWR _00984_ sky130_fd_sc_hd__and2b_1
XFILLER_0_66_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12630_ _07711_ _00193_ _02685_ VGND VGND VPWR VPWR _02723_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_66_733 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12561_ _02643_ _02652_ _02613_ _02653_ VGND VGND VPWR VPWR _02654_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_109_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14300_ _04500_ _04499_ VGND VGND VPWR VPWR _04502_ sky130_fd_sc_hd__or2b_1
X_11512_ _01551_ _01560_ VGND VGND VPWR VPWR _01605_ sky130_fd_sc_hd__nand2_1
XFILLER_0_108_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15280_ _05554_ _05555_ _05570_ VGND VGND VPWR VPWR _05571_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_124_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12492_ _02460_ _02472_ VGND VGND VPWR VPWR _02585_ sky130_fd_sc_hd__nand2_1
XFILLER_0_81_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14231_ _04332_ _04333_ VGND VGND VPWR VPWR _04426_ sky130_fd_sc_hd__or2b_1
X_11443_ _04362_ _00176_ _00145_ _04635_ VGND VGND VPWR VPWR _01536_ sky130_fd_sc_hd__a22o_1
XFILLER_0_124_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire145 _07389_ VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__buf_2
XFILLER_0_22_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_279 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_123_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14162_ _04338_ _04183_ _04349_ VGND VGND VPWR VPWR _04352_ sky130_fd_sc_hd__nand3_1
X_11374_ _01465_ _01464_ _01462_ VGND VGND VPWR VPWR _01467_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_33_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_195 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_150_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13113_ _03629_ _03596_ _05039_ _04460_ VGND VGND VPWR VPWR _03208_ sky130_fd_sc_hd__nand4_2
X_10325_ _00379_ _09342_ _00416_ _00417_ VGND VGND VPWR VPWR _00418_ sky130_fd_sc_hd__a211o_2
XFILLER_0_132_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14093_ _04273_ _04275_ VGND VGND VPWR VPWR _04276_ sky130_fd_sc_hd__or2b_1
X_18970_ clknet_4_4_0_clk _09401_ VGND VGND VPWR VPWR salida\[23\] sky130_fd_sc_hd__dfxtp_1
XTAP_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17921_ _06390_ _06790_ _08440_ _04336_ VGND VGND VPWR VPWR _08441_ sky130_fd_sc_hd__a22o_1
X_13044_ _03028_ _01136_ VGND VGND VPWR VPWR _03136_ sky130_fd_sc_hd__nor2_1
X_10256_ _00337_ _00338_ _00348_ VGND VGND VPWR VPWR _00349_ sky130_fd_sc_hd__a21o_2
XFILLER_0_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17852_ _08363_ _08364_ VGND VGND VPWR VPWR _08366_ sky130_fd_sc_hd__nand2_1
X_10187_ _08344_ _08354_ _08333_ VGND VGND VPWR VPWR _00280_ sky130_fd_sc_hd__a21bo_1
X_16803_ _07220_ _07222_ VGND VGND VPWR VPWR _07223_ sky130_fd_sc_hd__xnor2_1
X_17783_ _08277_ _08290_ VGND VGND VPWR VPWR _08291_ sky130_fd_sc_hd__xnor2_1
X_14995_ _05244_ _05245_ _05259_ VGND VGND VPWR VPWR _05261_ sky130_fd_sc_hd__or3_1
Xclkbuf_4_11_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_11_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_88_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16734_ _07146_ _07147_ VGND VGND VPWR VPWR _07148_ sky130_fd_sc_hd__and2_1
X_13946_ _04113_ _04114_ VGND VGND VPWR VPWR _04115_ sky130_fd_sc_hd__or2_1
XFILLER_0_72_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16665_ _02798_ _02830_ VGND VGND VPWR VPWR _07073_ sky130_fd_sc_hd__or2b_1
X_13877_ _04028_ _04039_ VGND VGND VPWR VPWR _04040_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_57_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18404_ _08964_ VGND VGND VPWR VPWR _08965_ sky130_fd_sc_hd__buf_1
X_15616_ _05934_ _05936_ VGND VGND VPWR VPWR _05937_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_57_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12828_ _00592_ _00214_ _00886_ VGND VGND VPWR VPWR _02921_ sky130_fd_sc_hd__and3_1
X_16596_ _06703_ _06707_ _06709_ _06715_ _03062_ _03081_ VGND VGND VPWR VPWR _06998_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_118_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18335_ _08880_ _08886_ _08890_ VGND VGND VPWR VPWR _08891_ sky130_fd_sc_hd__and3b_1
X_15547_ _05859_ _05860_ _05771_ _05808_ VGND VGND VPWR VPWR _05862_ sky130_fd_sc_hd__o211a_1
XTAP_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12759_ _01239_ _01246_ VGND VGND VPWR VPWR _02852_ sky130_fd_sc_hd__and2_1
XFILLER_0_72_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_122_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18266_ _08752_ _08754_ _08751_ VGND VGND VPWR VPWR _08816_ sky130_fd_sc_hd__a21o_1
X_15478_ _05703_ _05706_ VGND VGND VPWR VPWR _05787_ sky130_fd_sc_hd__and2b_1
XFILLER_0_4_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17217_ _07669_ _07670_ _07672_ VGND VGND VPWR VPWR _07674_ sky130_fd_sc_hd__or3_1
XFILLER_0_142_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14429_ _04641_ _04642_ VGND VGND VPWR VPWR _04643_ sky130_fd_sc_hd__or2_2
XFILLER_0_126_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18197_ _08739_ _08740_ VGND VGND VPWR VPWR _08741_ sky130_fd_sc_hd__or2_1
XFILLER_0_142_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17148_ _07594_ _07597_ VGND VGND VPWR VPWR _07598_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09970_ _09145_ _09037_ _09048_ VGND VGND VPWR VPWR _09158_ sky130_fd_sc_hd__and3_1
X_17079_ _07521_ _07522_ VGND VGND VPWR VPWR _07523_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_122_392 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_703 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_118_632 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_838 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_132_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_120_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10110_ cla_inst.in2\[21\] VGND VGND VPWR VPWR _00203_ sky130_fd_sc_hd__clkbuf_4
X_11090_ _05213_ _04864_ VGND VGND VPWR VPWR _01183_ sky130_fd_sc_hd__and2_1
X_10041_ _00132_ VGND VGND VPWR VPWR _00134_ sky130_fd_sc_hd__buf_4
Xsplit9 _03366_ VGND VGND VPWR VPWR net172 sky130_fd_sc_hd__buf_8
X_13800_ _03953_ _03954_ _04548_ _07374_ VGND VGND VPWR VPWR _03955_ sky130_fd_sc_hd__and4bb_1
Xhold86 salida\[0\] VGND VGND VPWR VPWR net249 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold97 _00007_ VGND VGND VPWR VPWR net260 sky130_fd_sc_hd__dlygate4sd3_1
X_14780_ _05023_ _05024_ _05019_ VGND VGND VPWR VPWR _05026_ sky130_fd_sc_hd__a21oi_1
X_11992_ _04690_ _00127_ VGND VGND VPWR VPWR _02085_ sky130_fd_sc_hd__nand2_1
X_13731_ _03877_ _03878_ _03667_ _03838_ VGND VGND VPWR VPWR _03880_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_58_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10943_ _01029_ _01030_ _01035_ VGND VGND VPWR VPWR _01036_ sky130_fd_sc_hd__a21o_1
XFILLER_0_85_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16450_ _02972_ _06837_ _06838_ VGND VGND VPWR VPWR _06839_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_38_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13662_ _03789_ _03802_ _03803_ VGND VGND VPWR VPWR _03805_ sky130_fd_sc_hd__nand3_2
XFILLER_0_42_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10874_ _00918_ net190 _00966_ VGND VGND VPWR VPWR _00967_ sky130_fd_sc_hd__o21a_1
XFILLER_0_66_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15401_ _05700_ _05702_ VGND VGND VPWR VPWR _05703_ sky130_fd_sc_hd__xnor2_1
X_12613_ _02664_ _02663_ _02658_ VGND VGND VPWR VPWR _02706_ sky130_fd_sc_hd__a21oi_1
X_13593_ _03727_ _03729_ VGND VGND VPWR VPWR _03730_ sky130_fd_sc_hd__nand2_1
X_16381_ _06758_ _06761_ _00132_ VGND VGND VPWR VPWR _06764_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_94_872 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18120_ _08655_ _08656_ VGND VGND VPWR VPWR _08657_ sky130_fd_sc_hd__or2_1
X_15332_ _05604_ _05605_ _05610_ VGND VGND VPWR VPWR _05628_ sky130_fd_sc_hd__or3b_1
X_12544_ _07243_ _01031_ _09179_ _07221_ VGND VGND VPWR VPWR _02637_ sky130_fd_sc_hd__a22o_1
XFILLER_0_108_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18051_ _08497_ _08530_ _08581_ VGND VGND VPWR VPWR _08582_ sky130_fd_sc_hd__a21oi_2
X_15263_ _05480_ _05496_ VGND VGND VPWR VPWR _05553_ sky130_fd_sc_hd__or2_1
X_12475_ _02482_ _02532_ _02567_ VGND VGND VPWR VPWR _02568_ sky130_fd_sc_hd__or3b_1
XFILLER_0_41_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17002_ _06749_ _07216_ _07437_ VGND VGND VPWR VPWR _07440_ sky130_fd_sc_hd__a21o_1
X_11426_ _03574_ _03662_ _09188_ _07591_ VGND VGND VPWR VPWR _01519_ sky130_fd_sc_hd__and4_1
X_14214_ _04068_ _04070_ _04236_ _04405_ _04408_ VGND VGND VPWR VPWR _04409_ sky130_fd_sc_hd__o311a_1
X_15194_ _05461_ _05462_ _05477_ VGND VGND VPWR VPWR _05478_ sky130_fd_sc_hd__o21ai_2
XANTENNA_6 _00309_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14145_ _04146_ _04167_ VGND VGND VPWR VPWR _04333_ sky130_fd_sc_hd__or2b_1
X_11357_ _01448_ _01446_ _01449_ VGND VGND VPWR VPWR _01450_ sky130_fd_sc_hd__or3_4
XFILLER_0_67_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_26 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10308_ _00258_ _00259_ VGND VGND VPWR VPWR _00401_ sky130_fd_sc_hd__and2_1
X_18953_ clknet_4_1_0_clk _09414_ VGND VGND VPWR VPWR salida\[6\] sky130_fd_sc_hd__dfxtp_1
X_14076_ _03537_ _04256_ VGND VGND VPWR VPWR _04257_ sky130_fd_sc_hd__and2_1
XTAP_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11288_ _00779_ _00793_ _00792_ VGND VGND VPWR VPWR _01381_ sky130_fd_sc_hd__a21o_1
XTAP_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13027_ _03119_ VGND VGND VPWR VPWR _03120_ sky130_fd_sc_hd__buf_2
X_17904_ _02846_ _02850_ _02469_ VGND VGND VPWR VPWR _08423_ sky130_fd_sc_hd__a21oi_2
X_10239_ _00303_ _00304_ _08529_ _08659_ VGND VGND VPWR VPWR _00332_ sky130_fd_sc_hd__a211o_1
X_18884_ clknet_4_8_0_clk _00038_ VGND VGND VPWR VPWR ApproximateM_inst.lob_16.lob1.genblk1\[2\].genblk1.mux.sel
+ sky130_fd_sc_hd__dfxtp_4
X_17835_ _08316_ _08317_ VGND VGND VPWR VPWR _08347_ sky130_fd_sc_hd__nand2_1
Xrebuffer18 net332 VGND VGND VPWR VPWR net181 sky130_fd_sc_hd__buf_1
XFILLER_0_83_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17766_ _08266_ _08270_ VGND VGND VPWR VPWR _08272_ sky130_fd_sc_hd__nand2_1
X_14978_ _05121_ _05122_ _05241_ VGND VGND VPWR VPWR _05242_ sky130_fd_sc_hd__o21ai_2
Xrebuffer29 net216 VGND VGND VPWR VPWR net192 sky130_fd_sc_hd__clkbuf_1
X_16717_ _07127_ _07128_ VGND VGND VPWR VPWR _07129_ sky130_fd_sc_hd__and2b_1
X_13929_ _03574_ _08757_ _04093_ _04094_ VGND VGND VPWR VPWR _04096_ sky130_fd_sc_hd__o2bb2a_1
X_17697_ _08188_ _08196_ VGND VGND VPWR VPWR _08197_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_76_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16648_ _07050_ _07052_ VGND VGND VPWR VPWR _07054_ sky130_fd_sc_hd__nor2_1
XFILLER_0_119_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16579_ _06976_ _06978_ VGND VGND VPWR VPWR _06979_ sky130_fd_sc_hd__xor2_1
XFILLER_0_85_883 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18318_ _08870_ _08871_ VGND VGND VPWR VPWR _08872_ sky130_fd_sc_hd__xor2_1
XFILLER_0_17_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18249_ _08716_ _08722_ _08720_ VGND VGND VPWR VPWR _08797_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_114_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_114_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09953_ _08659_ _08670_ _06373_ _08322_ VGND VGND VPWR VPWR _08995_ sky130_fd_sc_hd__o211ai_4
XTAP_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09884_ _08202_ _08213_ _08235_ VGND VGND VPWR VPWR _08246_ sky130_fd_sc_hd__or3_2
XTAP_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_817 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10590_ _00362_ _00223_ _00680_ _00681_ VGND VGND VPWR VPWR _00683_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_63_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12260_ _02243_ _02251_ VGND VGND VPWR VPWR _02353_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_31_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11211_ _01293_ _01294_ _01303_ VGND VGND VPWR VPWR _01304_ sky130_fd_sc_hd__a21o_1
X_12191_ _02132_ _02283_ VGND VGND VPWR VPWR _02284_ sky130_fd_sc_hd__nand2_1
XFILLER_0_120_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11142_ _01077_ _01203_ _01181_ _01201_ VGND VGND VPWR VPWR _01235_ sky130_fd_sc_hd__o211a_1
XFILLER_0_101_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput76 net76 VGND VGND VPWR VPWR leds[4] sky130_fd_sc_hd__clkbuf_4
Xoutput87 net87 VGND VGND VPWR VPWR o_wb_data[13] sky130_fd_sc_hd__clkbuf_4
X_11073_ _01149_ _01150_ _01165_ VGND VGND VPWR VPWR _01166_ sky130_fd_sc_hd__and3_2
X_15950_ _04823_ _06289_ _06290_ _06291_ _06296_ VGND VGND VPWR VPWR _09375_ sky130_fd_sc_hd__a32o_1
Xoutput98 net98 VGND VGND VPWR VPWR o_wb_data[23] sky130_fd_sc_hd__clkbuf_4
X_14901_ _05141_ _05142_ _05157_ VGND VGND VPWR VPWR _05158_ sky130_fd_sc_hd__o21a_1
X_10024_ _00114_ _00116_ VGND VGND VPWR VPWR _00117_ sky130_fd_sc_hd__nor2_1
X_15881_ _06178_ _06222_ VGND VGND VPWR VPWR _06223_ sky130_fd_sc_hd__or2_1
X_17620_ _08111_ _08112_ VGND VGND VPWR VPWR _08113_ sky130_fd_sc_hd__xor2_1
X_14832_ _03097_ _03106_ _03062_ VGND VGND VPWR VPWR _05084_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17551_ _06462_ _08035_ _08037_ VGND VGND VPWR VPWR _08038_ sky130_fd_sc_hd__or3b_1
X_14763_ _05004_ _05007_ VGND VGND VPWR VPWR _05008_ sky130_fd_sc_hd__or2_1
X_11975_ _02027_ _02051_ _02042_ _02050_ VGND VGND VPWR VPWR _02068_ sky130_fd_sc_hd__o211a_1
XFILLER_0_59_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16502_ _06893_ _06894_ VGND VGND VPWR VPWR _06896_ sky130_fd_sc_hd__xnor2_2
X_13714_ _03653_ _03659_ VGND VGND VPWR VPWR _03862_ sky130_fd_sc_hd__or2_1
X_10926_ _00978_ _00979_ net195 _00955_ VGND VGND VPWR VPWR _01019_ sky130_fd_sc_hd__a211oi_2
X_17482_ _07956_ _07961_ VGND VGND VPWR VPWR _07963_ sky130_fd_sc_hd__xnor2_1
X_14694_ _04758_ _04803_ _04931_ VGND VGND VPWR VPWR _04933_ sky130_fd_sc_hd__and3_1
X_16433_ _06800_ _06820_ VGND VGND VPWR VPWR _06821_ sky130_fd_sc_hd__xor2_1
X_13645_ _03606_ _03753_ _03784_ _03785_ VGND VGND VPWR VPWR _03786_ sky130_fd_sc_hd__o211a_2
XFILLER_0_73_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10857_ _04416_ _03399_ _00949_ _04493_ VGND VGND VPWR VPWR _00950_ sky130_fd_sc_hd__a22o_1
XFILLER_0_66_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16364_ _03916_ _06745_ VGND VGND VPWR VPWR _06746_ sky130_fd_sc_hd__nor2_1
X_13576_ _03447_ _03710_ VGND VGND VPWR VPWR _03711_ sky130_fd_sc_hd__xor2_1
X_10788_ _00207_ VGND VGND VPWR VPWR _00881_ sky130_fd_sc_hd__buf_4
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18103_ _07604_ _07623_ _08638_ VGND VGND VPWR VPWR _08639_ sky130_fd_sc_hd__and3_1
X_15315_ _05608_ _05609_ VGND VGND VPWR VPWR _05610_ sky130_fd_sc_hd__nand2_1
X_12527_ _02538_ _02539_ VGND VGND VPWR VPWR _02620_ sky130_fd_sc_hd__nand2_1
XFILLER_0_124_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16295_ _06649_ _06669_ _06670_ VGND VGND VPWR VPWR _06671_ sky130_fd_sc_hd__and3_1
XFILLER_0_41_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18034_ _08469_ _08480_ _08468_ VGND VGND VPWR VPWR _08564_ sky130_fd_sc_hd__a21o_1
XFILLER_0_151_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15246_ _05532_ _05533_ VGND VGND VPWR VPWR _05534_ sky130_fd_sc_hd__nor2_1
X_12458_ _07984_ _07973_ _00145_ _00196_ VGND VGND VPWR VPWR _02551_ sky130_fd_sc_hd__nand4_2
XFILLER_0_2_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11409_ _01501_ VGND VGND VPWR VPWR _01502_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15177_ _05457_ _05458_ VGND VGND VPWR VPWR _05459_ sky130_fd_sc_hd__nor2_1
X_12389_ _02479_ _02481_ VGND VGND VPWR VPWR _02482_ sky130_fd_sc_hd__and2_1
X_14128_ _04299_ _04300_ _04312_ VGND VGND VPWR VPWR _04314_ sky130_fd_sc_hd__o21ai_2
X_18936_ clknet_4_2_0_clk _00090_ VGND VGND VPWR VPWR cla_inst.in2\[22\] sky130_fd_sc_hd__dfxtp_1
X_14059_ _04065_ _04072_ _04236_ _04238_ VGND VGND VPWR VPWR _04239_ sky130_fd_sc_hd__a31o_1
X_18867_ clknet_4_7_0_clk net304 VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__dfxtp_1
X_17818_ _02985_ _06511_ _01695_ VGND VGND VPWR VPWR _08329_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_118_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18798_ _09298_ _09307_ VGND VGND VPWR VPWR _09308_ sky130_fd_sc_hd__and2_1
XFILLER_0_118_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17749_ _08212_ _08211_ VGND VGND VPWR VPWR _08253_ sky130_fd_sc_hd__or2b_1
XFILLER_0_49_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_134_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_791 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_143_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_162 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_772 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09936_ _05834_ _06094_ _06624_ _06602_ VGND VGND VPWR VPWR _08811_ sky130_fd_sc_hd__a31o_1
XFILLER_0_110_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09867_ _06019_ _08039_ _06613_ _08049_ VGND VGND VPWR VPWR _08060_ sky130_fd_sc_hd__and4_1
XTAP_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09798_ _07178_ _07199_ _07189_ VGND VGND VPWR VPWR _07308_ sky130_fd_sc_hd__a21o_1
XTAP_2503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11760_ _06971_ _04460_ VGND VGND VPWR VPWR _01853_ sky130_fd_sc_hd__nand2_1
XTAP_2558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10711_ _08452_ _05910_ _05899_ VGND VGND VPWR VPWR _00804_ sky130_fd_sc_hd__a21bo_1
XTAP_1857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11691_ _01783_ VGND VGND VPWR VPWR _01784_ sky130_fd_sc_hd__inv_2
XTAP_1868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_628 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_680 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10642_ _00721_ _00722_ _00733_ _00734_ VGND VGND VPWR VPWR _00735_ sky130_fd_sc_hd__a211o_2
X_13430_ _03549_ _03550_ _02489_ VGND VGND VPWR VPWR _03551_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_270 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13361_ _03473_ _03474_ VGND VGND VPWR VPWR _03475_ sky130_fd_sc_hd__nor2_1
XFILLER_0_106_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10573_ _06993_ _00665_ _00501_ _00500_ VGND VGND VPWR VPWR _00666_ sky130_fd_sc_hd__a31o_1
XFILLER_0_63_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15100_ _05373_ _05374_ VGND VGND VPWR VPWR _05375_ sky130_fd_sc_hd__xor2_1
Xrebuffer9 _03810_ VGND VGND VPWR VPWR net326 sky130_fd_sc_hd__dlymetal6s2s_1
X_12312_ _02402_ _02404_ VGND VGND VPWR VPWR _02405_ sky130_fd_sc_hd__nand2_1
X_13292_ _04558_ _06732_ _03397_ _03398_ VGND VGND VPWR VPWR _03400_ sky130_fd_sc_hd__nand4_1
X_16080_ _00593_ _00248_ _06436_ VGND VGND VPWR VPWR _06437_ sky130_fd_sc_hd__and3_1
X_15031_ _05188_ _05206_ _05298_ VGND VGND VPWR VPWR _05300_ sky130_fd_sc_hd__a21oi_1
X_12243_ _02208_ _02331_ _02335_ VGND VGND VPWR VPWR _02336_ sky130_fd_sc_hd__or3_1
XFILLER_0_31_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12174_ _02234_ _02239_ _02266_ VGND VGND VPWR VPWR _02267_ sky130_fd_sc_hd__a21oi_2
X_11125_ _01217_ VGND VGND VPWR VPWR _01218_ sky130_fd_sc_hd__inv_2
X_16982_ _06968_ _06946_ _07026_ _06890_ VGND VGND VPWR VPWR _07418_ sky130_fd_sc_hd__a22o_1
X_18721_ _09245_ _09246_ VGND VGND VPWR VPWR _09247_ sky130_fd_sc_hd__and2_1
X_11056_ _01037_ _01028_ _01036_ VGND VGND VPWR VPWR _01149_ sky130_fd_sc_hd__nand3_1
X_15933_ _06273_ _06276_ VGND VGND VPWR VPWR _06279_ sky130_fd_sc_hd__nand2_1
X_10007_ _09349_ VGND VGND VPWR VPWR _09350_ sky130_fd_sc_hd__clkbuf_4
X_18652_ _09176_ _09196_ VGND VGND VPWR VPWR _09198_ sky130_fd_sc_hd__and2_1
X_15864_ _06155_ _06204_ VGND VGND VPWR VPWR _06205_ sky130_fd_sc_hd__xnor2_1
X_17603_ _08092_ _08094_ VGND VGND VPWR VPWR _08095_ sky130_fd_sc_hd__xnor2_1
X_14815_ _04967_ _04928_ _05063_ _05064_ VGND VGND VPWR VPWR _05065_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_59_603 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18583_ salida\[11\] _09141_ _09142_ salida\[43\] _09146_ VGND VGND VPWR VPWR _09147_
+ sky130_fd_sc_hd__a221o_1
X_15795_ _06086_ _06130_ VGND VGND VPWR VPWR _06131_ sky130_fd_sc_hd__or2_1
XFILLER_0_99_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17534_ _08016_ _08018_ _08019_ VGND VGND VPWR VPWR _08020_ sky130_fd_sc_hd__a21oi_1
X_14746_ _04986_ _04987_ _04845_ _04988_ VGND VGND VPWR VPWR _04989_ sky130_fd_sc_hd__a211o_1
X_11958_ _02009_ _02024_ _02026_ VGND VGND VPWR VPWR _02051_ sky130_fd_sc_hd__and3_1
XFILLER_0_47_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10909_ _05355_ _04384_ _04471_ _05399_ VGND VGND VPWR VPWR _01002_ sky130_fd_sc_hd__a22o_1
X_17465_ _02347_ _06891_ VGND VGND VPWR VPWR _07944_ sky130_fd_sc_hd__nand2_1
X_14677_ _04907_ _04913_ VGND VGND VPWR VPWR _04914_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_74_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11889_ _01868_ _01981_ VGND VGND VPWR VPWR _01982_ sky130_fd_sc_hd__xor2_1
X_16416_ _05213_ _03003_ _03004_ _06523_ VGND VGND VPWR VPWR _06802_ sky130_fd_sc_hd__or4_1
XFILLER_0_13_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13628_ _03765_ _03766_ VGND VGND VPWR VPWR _03767_ sky130_fd_sc_hd__xor2_2
XFILLER_0_73_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17396_ _07867_ _07868_ VGND VGND VPWR VPWR _07869_ sky130_fd_sc_hd__nand2_1
XFILLER_0_104_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16347_ _06724_ _06726_ _03061_ VGND VGND VPWR VPWR _06727_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13559_ _03689_ _03691_ VGND VGND VPWR VPWR _03692_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_125_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_227 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16278_ _06427_ _06651_ VGND VGND VPWR VPWR _06652_ sky130_fd_sc_hd__or2_1
XFILLER_0_125_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18017_ _08537_ _08544_ VGND VGND VPWR VPWR _08545_ sky130_fd_sc_hd__xor2_1
X_15229_ _05426_ _05427_ _05515_ VGND VGND VPWR VPWR _05516_ sky130_fd_sc_hd__o21a_1
XFILLER_0_140_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09721_ _05497_ VGND VGND VPWR VPWR _06471_ sky130_fd_sc_hd__buf_6
X_18919_ clknet_4_8_0_clk _00073_ VGND VGND VPWR VPWR ApproximateM_inst.lob_16.lob2.genblk1\[5\].genblk1.mux.sel
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_0_38_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09652_ _05627_ _05660_ _05682_ _05715_ VGND VGND VPWR VPWR _05725_ sky130_fd_sc_hd__and4b_1
XFILLER_0_78_901 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_145_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09583_ _04941_ _04952_ _04962_ VGND VGND VPWR VPWR _04973_ sky130_fd_sc_hd__nand3_2
XFILLER_0_145_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_145_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_130_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold150 salida\[3\] VGND VGND VPWR VPWR net313 sky130_fd_sc_hd__buf_1
XFILLER_0_130_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09919_ _08615_ _05888_ _06417_ _06406_ VGND VGND VPWR VPWR _08626_ sky130_fd_sc_hd__a31o_1
X_12930_ _03022_ VGND VGND VPWR VPWR _03023_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_87_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12861_ _02945_ _02952_ _02953_ _00904_ VGND VGND VPWR VPWR _02954_ sky130_fd_sc_hd__a211o_1
XTAP_2311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14600_ _02976_ _03038_ _04826_ _04829_ _03121_ VGND VGND VPWR VPWR _04830_ sky130_fd_sc_hd__o32a_1
XTAP_2333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11812_ _04132_ _04984_ _07559_ _07602_ VGND VGND VPWR VPWR _01905_ sky130_fd_sc_hd__nand4_4
XTAP_2344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15580_ _09351_ _07744_ _05896_ VGND VGND VPWR VPWR _05897_ sky130_fd_sc_hd__a21oi_1
XTAP_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12792_ _02876_ _02875_ VGND VGND VPWR VPWR _02885_ sky130_fd_sc_hd__and2b_1
XTAP_2366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14531_ _04741_ _04742_ _04753_ VGND VGND VPWR VPWR _04754_ sky130_fd_sc_hd__a21oi_1
XTAP_1643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11743_ _01832_ _01835_ VGND VGND VPWR VPWR _01836_ sky130_fd_sc_hd__and2b_1
XTAP_2399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17250_ _06756_ _07410_ _07708_ _06542_ VGND VGND VPWR VPWR _07709_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_138_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14462_ _04676_ _04677_ _04566_ _04538_ VGND VGND VPWR VPWR _04680_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_50_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11674_ _01722_ _01723_ _01724_ _01732_ VGND VGND VPWR VPWR _01767_ sky130_fd_sc_hd__a31o_1
X_16201_ _00210_ _06528_ _06530_ _06533_ VGND VGND VPWR VPWR _06568_ sky130_fd_sc_hd__or4_4
X_13413_ _03032_ _03085_ _03089_ VGND VGND VPWR VPWR _03533_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10625_ _00714_ _00717_ VGND VGND VPWR VPWR _00718_ sky130_fd_sc_hd__xor2_2
X_17181_ _07630_ _07126_ _07632_ _07633_ VGND VGND VPWR VPWR _07634_ sky130_fd_sc_hd__or4_1
XFILLER_0_37_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14393_ _04304_ _04600_ _04601_ VGND VGND VPWR VPWR _04604_ sky130_fd_sc_hd__or3_1
XFILLER_0_51_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_153_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16132_ _06488_ _06492_ _03061_ VGND VGND VPWR VPWR _06494_ sky130_fd_sc_hd__mux2_1
X_10556_ _05834_ _08876_ _00647_ _00648_ VGND VGND VPWR VPWR _00649_ sky130_fd_sc_hd__nand4_2
X_13344_ _07091_ _00513_ VGND VGND VPWR VPWR _03457_ sky130_fd_sc_hd__nand2_1
XFILLER_0_106_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16063_ _03292_ _03217_ VGND VGND VPWR VPWR _06419_ sky130_fd_sc_hd__or2_1
XFILLER_0_121_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10487_ _00396_ _00538_ _00578_ _00579_ VGND VGND VPWR VPWR _00580_ sky130_fd_sc_hd__a211oi_2
X_13275_ _03207_ _03209_ _03208_ VGND VGND VPWR VPWR _03381_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_122_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15014_ _05281_ VGND VGND VPWR VPWR _05282_ sky130_fd_sc_hd__inv_2
X_12226_ _02317_ _02318_ VGND VGND VPWR VPWR _02319_ sky130_fd_sc_hd__nor2_1
X_12157_ _02248_ _02249_ VGND VGND VPWR VPWR _02250_ sky130_fd_sc_hd__xnor2_2
X_11108_ _01181_ _01198_ _01199_ _01200_ VGND VGND VPWR VPWR _01201_ sky130_fd_sc_hd__nand4_2
X_12088_ _08713_ _00147_ _02179_ _02180_ VGND VGND VPWR VPWR _02181_ sky130_fd_sc_hd__and4_1
X_16965_ _06766_ _07106_ _07398_ VGND VGND VPWR VPWR _07399_ sky130_fd_sc_hd__or3_1
X_11039_ _01126_ _01130_ _01131_ VGND VGND VPWR VPWR _01132_ sky130_fd_sc_hd__nand3_1
X_18704_ net52 _03056_ _09182_ VGND VGND VPWR VPWR _09234_ sky130_fd_sc_hd__mux2_1
X_15916_ _06178_ _06221_ VGND VGND VPWR VPWR _06261_ sky130_fd_sc_hd__nand2_1
X_16896_ _07322_ _07323_ VGND VGND VPWR VPWR _07324_ sky130_fd_sc_hd__nand2_1
X_18635_ _09182_ VGND VGND VPWR VPWR _09183_ sky130_fd_sc_hd__buf_2
X_15847_ _06184_ _06186_ VGND VGND VPWR VPWR _06187_ sky130_fd_sc_hd__and2_1
XFILLER_0_152_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18566_ salida\[5\] _09114_ _09118_ salida\[37\] _09128_ VGND VGND VPWR VPWR _09134_
+ sky130_fd_sc_hd__a221o_1
X_15778_ _06032_ _06110_ VGND VGND VPWR VPWR _06112_ sky130_fd_sc_hd__nor2_1
XFILLER_0_87_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17517_ _07855_ _07876_ _08000_ VGND VGND VPWR VPWR _08001_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_24_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14729_ _01520_ _07722_ _07406_ _03651_ VGND VGND VPWR VPWR _04970_ sky130_fd_sc_hd__a22o_1
XFILLER_0_74_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18497_ _03155_ _09064_ VGND VGND VPWR VPWR _09065_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17448_ _06376_ _06372_ _06375_ _06598_ _07925_ VGND VGND VPWR VPWR _07926_ sky130_fd_sc_hd__a311o_1
X_17379_ _07840_ _07849_ VGND VGND VPWR VPWR _07850_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_40_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_880 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09704_ _04121_ _04395_ _04657_ _04088_ VGND VGND VPWR VPWR _06288_ sky130_fd_sc_hd__a22oi_2
X_09635_ _05475_ _05529_ VGND VGND VPWR VPWR _05540_ sky130_fd_sc_hd__and2_1
XFILLER_0_97_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09566_ _03465_ _03410_ VGND VGND VPWR VPWR _04788_ sky130_fd_sc_hd__and2_1
XFILLER_0_139_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09497_ _03793_ VGND VGND VPWR VPWR _04034_ sky130_fd_sc_hd__buf_8
XFILLER_0_93_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_135_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10410_ _07363_ _00502_ VGND VGND VPWR VPWR _00503_ sky130_fd_sc_hd__nand2_1
XFILLER_0_151_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11390_ _01473_ _01482_ VGND VGND VPWR VPWR _01483_ sky130_fd_sc_hd__and2_1
XFILLER_0_60_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10341_ _03377_ _04384_ _04886_ _03356_ VGND VGND VPWR VPWR _00434_ sky130_fd_sc_hd__a22o_1
X_13060_ _01677_ VGND VGND VPWR VPWR _03152_ sky130_fd_sc_hd__clkbuf_4
X_10272_ _00355_ _00356_ _00364_ VGND VGND VPWR VPWR _00365_ sky130_fd_sc_hd__and3_1
XFILLER_0_131_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12011_ _02088_ _02089_ VGND VGND VPWR VPWR _02104_ sky130_fd_sc_hd__xor2_1
X_16750_ _02533_ _06510_ _00214_ VGND VGND VPWR VPWR _07165_ sky130_fd_sc_hd__a21bo_1
X_13962_ _05453_ _00645_ _00502_ _09248_ VGND VGND VPWR VPWR _04133_ sky130_fd_sc_hd__and4_1
XFILLER_0_45_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15701_ _06024_ _06027_ VGND VGND VPWR VPWR _06028_ sky130_fd_sc_hd__and2_1
X_12913_ _03005_ VGND VGND VPWR VPWR _03006_ sky130_fd_sc_hd__clkbuf_4
Xmax_cap7 _01329_ VGND VGND VPWR VPWR net325 sky130_fd_sc_hd__buf_1
X_16681_ _06741_ _06736_ _06738_ _06731_ _03912_ _03077_ VGND VGND VPWR VPWR _07090_
+ sky130_fd_sc_hd__mux4_2
X_13893_ _04055_ _04057_ VGND VGND VPWR VPWR _04058_ sky130_fd_sc_hd__nand2_2
X_18420_ _08926_ _08928_ _08925_ VGND VGND VPWR VPWR _08982_ sky130_fd_sc_hd__a21o_1
XTAP_2130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15632_ _04080_ _05623_ _05881_ _03125_ _05953_ VGND VGND VPWR VPWR _09368_ sky130_fd_sc_hd__a221o_1
X_12844_ _02913_ _02935_ _02934_ _02933_ VGND VGND VPWR VPWR _02937_ sky130_fd_sc_hd__a211o_1
XFILLER_0_69_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18351_ _08903_ _08905_ VGND VGND VPWR VPWR _08907_ sky130_fd_sc_hd__nand2_1
XTAP_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15563_ _05875_ _05877_ _05879_ VGND VGND VPWR VPWR _05880_ sky130_fd_sc_hd__a21oi_2
XTAP_2185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12775_ _02867_ _01808_ VGND VGND VPWR VPWR _02868_ sky130_fd_sc_hd__nor2_1
XTAP_2196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17302_ _07735_ _07765_ VGND VGND VPWR VPWR _07767_ sky130_fd_sc_hd__nor2_1
X_14514_ _04723_ _04724_ _04734_ VGND VGND VPWR VPWR _04736_ sky130_fd_sc_hd__or3_4
XTAP_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18282_ _01417_ _06512_ _03143_ VGND VGND VPWR VPWR _08833_ sky130_fd_sc_hd__a21bo_1
X_11726_ _01817_ _01818_ VGND VGND VPWR VPWR _01819_ sky130_fd_sc_hd__xor2_1
XTAP_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15494_ _05803_ _03918_ _03547_ VGND VGND VPWR VPWR _05804_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17233_ _06369_ _06790_ _07691_ _06368_ VGND VGND VPWR VPWR _07692_ sky130_fd_sc_hd__a22o_1
X_14445_ _04654_ _04660_ VGND VGND VPWR VPWR _04661_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_83_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11657_ _01748_ _01749_ VGND VGND VPWR VPWR _01750_ sky130_fd_sc_hd__and2_1
XFILLER_0_154_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10608_ _00562_ _00570_ VGND VGND VPWR VPWR _00701_ sky130_fd_sc_hd__or2b_1
X_17164_ _07603_ net238 VGND VGND VPWR VPWR _07616_ sky130_fd_sc_hd__xor2_1
X_14376_ _04581_ _04582_ _04583_ VGND VGND VPWR VPWR _04585_ sky130_fd_sc_hd__a21oi_1
X_11588_ _01670_ _01676_ _01679_ _01680_ VGND VGND VPWR VPWR _01681_ sky130_fd_sc_hd__or4_1
XFILLER_0_141_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16115_ _03027_ _03166_ _02685_ _02983_ VGND VGND VPWR VPWR _06475_ sky130_fd_sc_hd__a211o_1
X_13327_ _03258_ _03261_ VGND VGND VPWR VPWR _03438_ sky130_fd_sc_hd__and2b_1
XFILLER_0_122_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10539_ _00620_ _00621_ _00631_ VGND VGND VPWR VPWR _00632_ sky130_fd_sc_hd__o21ai_2
X_17095_ _07539_ _07426_ _07540_ VGND VGND VPWR VPWR _07541_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_150_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16046_ _06398_ _06399_ _05368_ VGND VGND VPWR VPWR _06400_ sky130_fd_sc_hd__a21o_1
X_13258_ _03358_ _03361_ VGND VGND VPWR VPWR _03363_ sky130_fd_sc_hd__or2_1
XFILLER_0_110_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12209_ _02290_ net322 _02151_ _02301_ VGND VGND VPWR VPWR _02302_ sky130_fd_sc_hd__o211a_4
XFILLER_0_110_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13189_ _03278_ _03288_ VGND VGND VPWR VPWR _03289_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_19_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17997_ _06392_ _06546_ _08523_ _00813_ VGND VGND VPWR VPWR _08524_ sky130_fd_sc_hd__o2bb2a_1
X_16948_ _07342_ _07343_ VGND VGND VPWR VPWR _07380_ sky130_fd_sc_hd__or2b_1
X_16879_ _07301_ _07304_ VGND VGND VPWR VPWR _07305_ sky130_fd_sc_hd__nor2_1
X_09420_ op_code\[2\] op_code\[3\] VGND VGND VPWR VPWR _03195_ sky130_fd_sc_hd__nand2_4
X_18618_ salida\[26\] _09159_ _09160_ salida\[58\] _09163_ VGND VGND VPWR VPWR _09170_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_126_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_149_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18549_ _09115_ net27 net1 VGND VGND VPWR VPWR _09120_ sky130_fd_sc_hd__or3b_1
XFILLER_0_118_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_145_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_644 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_118_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_480 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_530 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09618_ _05290_ VGND VGND VPWR VPWR _05355_ sky130_fd_sc_hd__buf_8
XFILLER_0_97_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10890_ _05290_ ApproximateM_inst.lob_16.lob1.genblk1\[14\].genblk1.mux.sel _03739_
+ ApproximateM_inst.lob_16.lob2.genblk1\[10\].genblk1.mux.sel VGND VGND VPWR VPWR
+ _00983_ sky130_fd_sc_hd__a22o_1
XFILLER_0_66_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09549_ _04558_ _04591_ VGND VGND VPWR VPWR _04602_ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12560_ _02605_ _02606_ _02612_ VGND VGND VPWR VPWR _02653_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_108_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11511_ _01564_ _01601_ _01602_ _01603_ VGND VGND VPWR VPWR _01604_ sky130_fd_sc_hd__nand4_2
XFILLER_0_108_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12491_ _02531_ _02583_ VGND VGND VPWR VPWR _02584_ sky130_fd_sc_hd__nor2_1
X_14230_ _04161_ _04335_ _04378_ _04379_ VGND VGND VPWR VPWR _04425_ sky130_fd_sc_hd__a211o_1
XFILLER_0_151_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11442_ _01533_ _01534_ VGND VGND VPWR VPWR _01535_ sky130_fd_sc_hd__or2_1
Xwire146 _07216_ VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__buf_2
XFILLER_0_123_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11373_ _01462_ _01464_ _01465_ VGND VGND VPWR VPWR _01466_ sky130_fd_sc_hd__nand3b_4
X_14161_ _04338_ _04183_ _04349_ VGND VGND VPWR VPWR _04350_ sky130_fd_sc_hd__a21o_1
XFILLER_0_132_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13112_ _03377_ _05039_ _04384_ _03356_ VGND VGND VPWR VPWR _03207_ sky130_fd_sc_hd__a22o_1
X_10324_ _00396_ _00397_ _00415_ VGND VGND VPWR VPWR _00417_ sky130_fd_sc_hd__and3_1
X_14092_ _04271_ _04272_ net174 _04095_ VGND VGND VPWR VPWR _04275_ sky130_fd_sc_hd__a211o_1
X_10255_ _00340_ _00347_ VGND VGND VPWR VPWR _00348_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_30_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17920_ _03368_ _06920_ _06921_ VGND VGND VPWR VPWR _08440_ sky130_fd_sc_hd__a21o_1
X_13043_ _01672_ _03134_ _03040_ VGND VGND VPWR VPWR _03135_ sky130_fd_sc_hd__o21a_1
X_17851_ _08349_ _08350_ _08362_ VGND VGND VPWR VPWR _08364_ sky130_fd_sc_hd__nand3_1
X_10186_ _00275_ _00277_ _00276_ VGND VGND VPWR VPWR _00279_ sky130_fd_sc_hd__a21o_1
X_16802_ _06579_ _07126_ VGND VGND VPWR VPWR _07222_ sky130_fd_sc_hd__or2_1
X_17782_ _08287_ _08288_ VGND VGND VPWR VPWR _08290_ sky130_fd_sc_hd__nor2_1
X_14994_ _05244_ _05245_ _05259_ VGND VGND VPWR VPWR _05260_ sky130_fd_sc_hd__o21ai_1
X_16733_ _07142_ _07144_ VGND VGND VPWR VPWR _07147_ sky130_fd_sc_hd__nand2_1
X_13945_ _04690_ _07722_ _04111_ _04112_ VGND VGND VPWR VPWR _04114_ sky130_fd_sc_hd__o2bb2a_1
X_16664_ _03206_ _07071_ VGND VGND VPWR VPWR _07072_ sky130_fd_sc_hd__nor2_1
X_13876_ _03823_ _04038_ VGND VGND VPWR VPWR _04039_ sky130_fd_sc_hd__xor2_1
X_15615_ _05935_ _05860_ VGND VGND VPWR VPWR _05936_ sky130_fd_sc_hd__nor2_1
X_18403_ _08961_ _08963_ VGND VGND VPWR VPWR _08964_ sky130_fd_sc_hd__or2_1
XFILLER_0_9_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12827_ _02918_ _02919_ VGND VGND VPWR VPWR _02920_ sky130_fd_sc_hd__nand2_1
X_16595_ _06343_ _06345_ _06995_ VGND VGND VPWR VPWR _06997_ sky130_fd_sc_hd__nand3_1
X_18334_ _08888_ _06402_ _06403_ _07084_ _08889_ VGND VGND VPWR VPWR _08890_ sky130_fd_sc_hd__a311o_1
XFILLER_0_84_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15546_ _05771_ _05808_ _05859_ _05860_ VGND VGND VPWR VPWR _05861_ sky130_fd_sc_hd__a211oi_2
XTAP_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12758_ _02176_ _02846_ _02850_ VGND VGND VPWR VPWR _02851_ sky130_fd_sc_hd__and3_1
XTAP_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18265_ _08813_ _08814_ VGND VGND VPWR VPWR _08815_ sky130_fd_sc_hd__nor2_1
X_11709_ _01771_ _01781_ _01800_ _01801_ VGND VGND VPWR VPWR _01802_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_84_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_20 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15477_ _05784_ _05785_ VGND VGND VPWR VPWR _05786_ sky130_fd_sc_hd__nand2_2
XFILLER_0_72_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_452 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12689_ _02713_ _02781_ VGND VGND VPWR VPWR _02782_ sky130_fd_sc_hd__nor2_1
X_17216_ _07669_ _07670_ _07672_ VGND VGND VPWR VPWR _07673_ sky130_fd_sc_hd__o21a_1
X_14428_ _04630_ _04640_ VGND VGND VPWR VPWR _04642_ sky130_fd_sc_hd__and2_1
X_18196_ _08696_ _08738_ VGND VGND VPWR VPWR _08740_ sky130_fd_sc_hd__and2_1
XFILLER_0_141_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17147_ _06542_ _07113_ _07489_ _07596_ VGND VGND VPWR VPWR _07597_ sky130_fd_sc_hd__and4_1
XFILLER_0_142_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14359_ _04315_ _04331_ _04487_ _04488_ VGND VGND VPWR VPWR _04566_ sky130_fd_sc_hd__o211a_1
XFILLER_0_24_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17078_ _06875_ _07035_ VGND VGND VPWR VPWR _07522_ sky130_fd_sc_hd__or2_1
XFILLER_0_97_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16029_ _02988_ _03111_ VGND VGND VPWR VPWR _06381_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_244 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_90 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10040_ _00126_ _00128_ _00106_ _00132_ VGND VGND VPWR VPWR _00133_ sky130_fd_sc_hd__and4b_1
Xhold87 net109 VGND VGND VPWR VPWR net250 sky130_fd_sc_hd__dlygate4sd3_1
X_11991_ _04438_ _09188_ _07591_ _04646_ VGND VGND VPWR VPWR _02084_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_97_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold98 net111 VGND VGND VPWR VPWR net261 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13730_ _03667_ _03838_ _03877_ _03878_ VGND VGND VPWR VPWR _03879_ sky130_fd_sc_hd__o211a_1
X_10942_ _01032_ _01033_ _01034_ VGND VGND VPWR VPWR _01035_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_98_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_129_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13661_ _03800_ _03801_ _03794_ VGND VGND VPWR VPWR _03803_ sky130_fd_sc_hd__a21o_1
XFILLER_0_97_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10873_ _00961_ _00965_ VGND VGND VPWR VPWR _00966_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_66_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15400_ _05600_ _05601_ _05701_ VGND VGND VPWR VPWR _05702_ sky130_fd_sc_hd__o21a_1
XFILLER_0_94_851 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12612_ _02664_ _02658_ _02663_ VGND VGND VPWR VPWR _02705_ sky130_fd_sc_hd__and3_1
X_16380_ net237 _06579_ _06657_ _06762_ VGND VGND VPWR VPWR _06763_ sky130_fd_sc_hd__and4bb_1
X_13592_ _03724_ _03725_ _03726_ VGND VGND VPWR VPWR _03729_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_94_884 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_108_110 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15331_ _05503_ _05506_ _05603_ VGND VGND VPWR VPWR _05626_ sky130_fd_sc_hd__a21o_1
XFILLER_0_54_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12543_ ApproximateM_inst.lob_16.lob2.genblk1\[2\].genblk1.mux.sel _00196_ VGND VGND
+ VPWR VPWR _02636_ sky130_fd_sc_hd__and2_1
X_18050_ _08578_ _08580_ VGND VGND VPWR VPWR _08581_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_151_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15262_ _05549_ _05550_ VGND VGND VPWR VPWR _05552_ sky130_fd_sc_hd__nand2_1
XFILLER_0_81_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12474_ _02542_ _02566_ VGND VGND VPWR VPWR _02567_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_123_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17001_ _06665_ _07318_ _07437_ VGND VGND VPWR VPWR _07438_ sky130_fd_sc_hd__or3b_1
X_14213_ _04233_ _04235_ _04407_ VGND VGND VPWR VPWR _04408_ sky130_fd_sc_hd__a21boi_1
X_11425_ _01516_ _01517_ VGND VGND VPWR VPWR _01518_ sky130_fd_sc_hd__xor2_1
XFILLER_0_124_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15193_ _05473_ _05476_ VGND VGND VPWR VPWR _05477_ sky130_fd_sc_hd__xnor2_1
XANTENNA_7 _00443_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_656 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_151_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14144_ _04330_ _04331_ VGND VGND VPWR VPWR _04332_ sky130_fd_sc_hd__or2_1
XFILLER_0_6_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11356_ _01444_ _01445_ _01370_ _01374_ VGND VGND VPWR VPWR _01449_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_22_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10307_ _00164_ _00399_ VGND VGND VPWR VPWR _00400_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18952_ clknet_4_1_0_clk _09413_ VGND VGND VPWR VPWR salida\[5\] sky130_fd_sc_hd__dfxtp_1
X_14075_ _03912_ _04254_ _04255_ VGND VGND VPWR VPWR _04256_ sky130_fd_sc_hd__o21ai_1
XTAP_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11287_ _01279_ _01286_ _01287_ VGND VGND VPWR VPWR _01380_ sky130_fd_sc_hd__nor3_1
XTAP_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17903_ _08413_ _08418_ _08421_ VGND VGND VPWR VPWR _08422_ sky130_fd_sc_hd__a21oi_1
XTAP_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13026_ _06765_ _03037_ VGND VGND VPWR VPWR _03119_ sky130_fd_sc_hd__nand2_2
X_10238_ _00326_ _00327_ _00329_ VGND VGND VPWR VPWR _00331_ sky130_fd_sc_hd__nand3_4
X_18883_ clknet_4_9_0_clk _00037_ VGND VGND VPWR VPWR ApproximateM_inst.lob_16.lob1.genblk1\[1\].genblk1.mux.sel
+ sky130_fd_sc_hd__dfxtp_4
X_10169_ _00250_ _00251_ _00261_ VGND VGND VPWR VPWR _00262_ sky130_fd_sc_hd__o21ai_1
X_17834_ _03041_ _06464_ net116 _08346_ VGND VGND VPWR VPWR _09396_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_89_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14977_ _05123_ _05134_ VGND VGND VPWR VPWR _05241_ sky130_fd_sc_hd__or2b_1
X_17765_ _08266_ _08270_ VGND VGND VPWR VPWR _08271_ sky130_fd_sc_hd__or2_1
Xrebuffer19 _01849_ VGND VGND VPWR VPWR net182 sky130_fd_sc_hd__clkbuf_1
X_13928_ _04093_ _04094_ _03574_ _08757_ VGND VGND VPWR VPWR _04095_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_89_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16716_ _06560_ _06951_ _06816_ _07125_ VGND VGND VPWR VPWR _07128_ sky130_fd_sc_hd__or4_4
X_17696_ _08194_ _08195_ VGND VGND VPWR VPWR _08196_ sky130_fd_sc_hd__xor2_1
XFILLER_0_16_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16647_ _07050_ _07052_ VGND VGND VPWR VPWR _07053_ sky130_fd_sc_hd__and2_1
X_13859_ _04019_ _03847_ VGND VGND VPWR VPWR _04020_ sky130_fd_sc_hd__nand2_1
XFILLER_0_85_862 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16578_ _06888_ _06896_ _06977_ VGND VGND VPWR VPWR _06978_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_32_63 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15529_ _05831_ _05749_ _05840_ VGND VGND VPWR VPWR _05842_ sky130_fd_sc_hd__and3_1
XFILLER_0_85_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18317_ _08802_ _08807_ VGND VGND VPWR VPWR _08871_ sky130_fd_sc_hd__nand2_1
XFILLER_0_123_87 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_127_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18248_ _08794_ _08795_ VGND VGND VPWR VPWR _08796_ sky130_fd_sc_hd__and2_1
XFILLER_0_25_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18179_ _08620_ _08622_ _08719_ VGND VGND VPWR VPWR _08721_ sky130_fd_sc_hd__and3_1
XFILLER_0_5_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09952_ _08951_ _08962_ _08930_ _08941_ VGND VGND VPWR VPWR _08984_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_0_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09883_ _07853_ _08224_ _07810_ VGND VGND VPWR VPWR _08235_ sky130_fd_sc_hd__a21oi_1
XTAP_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_4_10_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_10_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_31_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11210_ _01299_ _01302_ VGND VGND VPWR VPWR _01303_ sky130_fd_sc_hd__xnor2_1
X_12190_ _02129_ _02130_ _02131_ _02123_ VGND VGND VPWR VPWR _02283_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_102_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11141_ _01231_ _01232_ _01218_ _01228_ VGND VGND VPWR VPWR _01234_ sky130_fd_sc_hd__o211a_1
XFILLER_0_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11072_ _01156_ _01163_ _01164_ VGND VGND VPWR VPWR _01165_ sky130_fd_sc_hd__a21bo_1
Xoutput77 net77 VGND VGND VPWR VPWR leds[5] sky130_fd_sc_hd__buf_2
XFILLER_0_37_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput88 net88 VGND VGND VPWR VPWR o_wb_data[14] sky130_fd_sc_hd__clkbuf_4
Xoutput99 net99 VGND VGND VPWR VPWR o_wb_data[24] sky130_fd_sc_hd__clkbuf_4
X_14900_ _05155_ _05156_ VGND VGND VPWR VPWR _05157_ sky130_fd_sc_hd__xnor2_1
X_10023_ _00115_ _00108_ _00111_ _00113_ VGND VGND VPWR VPWR _00116_ sky130_fd_sc_hd__a22oi_1
X_15880_ _06128_ _06180_ VGND VGND VPWR VPWR _06222_ sky130_fd_sc_hd__nor2_1
X_14831_ _03033_ _03091_ _03062_ VGND VGND VPWR VPWR _05082_ sky130_fd_sc_hd__mux2_1
X_17550_ _03119_ _05423_ _06505_ _08036_ VGND VGND VPWR VPWR _08037_ sky130_fd_sc_hd__o22a_1
X_14762_ _07635_ _01866_ _05005_ _05002_ VGND VGND VPWR VPWR _05007_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_86_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11974_ _02056_ _02066_ VGND VGND VPWR VPWR _02067_ sky130_fd_sc_hd__or2b_1
X_16501_ _06749_ _06762_ VGND VGND VPWR VPWR _06894_ sky130_fd_sc_hd__nand2_1
X_13713_ _03701_ _03709_ _03860_ VGND VGND VPWR VPWR _03861_ sky130_fd_sc_hd__a21bo_1
X_10925_ _01016_ _01017_ VGND VGND VPWR VPWR _01018_ sky130_fd_sc_hd__nand2_1
X_17481_ _07959_ _07960_ VGND VGND VPWR VPWR _07961_ sky130_fd_sc_hd__xnor2_1
X_14693_ _04758_ _04803_ _04931_ VGND VGND VPWR VPWR _04932_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_86_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16432_ _06801_ _06818_ VGND VGND VPWR VPWR _06820_ sky130_fd_sc_hd__xnor2_1
X_13644_ _03772_ _03773_ _03783_ VGND VGND VPWR VPWR _03785_ sky130_fd_sc_hd__or3_4
X_10856_ ApproximateM_inst.lob_16.lob1.genblk1\[9\].genblk1.mux.sel VGND VGND VPWR
+ VPWR _00949_ sky130_fd_sc_hd__buf_4
XFILLER_0_94_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16363_ _03077_ _06741_ _06744_ _06487_ VGND VGND VPWR VPWR _06745_ sky130_fd_sc_hd__o2bb2a_1
X_13575_ _03701_ _03709_ VGND VGND VPWR VPWR _03710_ sky130_fd_sc_hd__xnor2_1
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10787_ _00877_ _00878_ _00879_ VGND VGND VPWR VPWR _00880_ sky130_fd_sc_hd__and3_1
XFILLER_0_93_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18102_ _07195_ _07741_ VGND VGND VPWR VPWR _08638_ sky130_fd_sc_hd__nor2_1
X_15314_ _03368_ _03072_ _05494_ VGND VGND VPWR VPWR _05609_ sky130_fd_sc_hd__nand3_1
XPHY_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_567 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12526_ net137 _02614_ _02604_ _02613_ VGND VGND VPWR VPWR _02619_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_124_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16294_ _06659_ _06668_ VGND VGND VPWR VPWR _06670_ sky130_fd_sc_hd__or2_1
XFILLER_0_82_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18033_ _08548_ _08562_ VGND VGND VPWR VPWR _08563_ sky130_fd_sc_hd__xor2_1
X_15245_ _05324_ _05439_ VGND VGND VPWR VPWR _05533_ sky130_fd_sc_hd__nand2_1
X_12457_ _02545_ _02548_ _02549_ VGND VGND VPWR VPWR _02550_ sky130_fd_sc_hd__nand3_1
XFILLER_0_112_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_442 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11408_ _01447_ _01450_ _01499_ _01500_ VGND VGND VPWR VPWR _01501_ sky130_fd_sc_hd__a211o_1
X_15176_ _05430_ _05342_ _05456_ VGND VGND VPWR VPWR _05458_ sky130_fd_sc_hd__and3_1
X_12388_ _02409_ _02480_ VGND VGND VPWR VPWR _02481_ sky130_fd_sc_hd__and2_1
XFILLER_0_1_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14127_ _04299_ _04300_ _04312_ VGND VGND VPWR VPWR _04313_ sky130_fd_sc_hd__or3_4
XFILLER_0_50_795 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11339_ _01430_ _01431_ VGND VGND VPWR VPWR _01432_ sky130_fd_sc_hd__and2_1
XFILLER_0_120_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18935_ clknet_4_2_0_clk _00089_ VGND VGND VPWR VPWR cla_inst.in2\[21\] sky130_fd_sc_hd__dfxtp_2
X_14058_ _02968_ VGND VGND VPWR VPWR _04238_ sky130_fd_sc_hd__clkbuf_8
X_13009_ _00593_ _03101_ _02505_ VGND VGND VPWR VPWR _03102_ sky130_fd_sc_hd__mux2_1
X_18866_ clknet_4_5_0_clk net309 VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__dfxtp_1
X_17817_ _08252_ _08223_ _08326_ VGND VGND VPWR VPWR _08328_ sky130_fd_sc_hd__nand3_1
X_18797_ _02998_ net49 _09301_ VGND VGND VPWR VPWR _09307_ sky130_fd_sc_hd__mux2_1
X_17748_ _08216_ _08217_ VGND VGND VPWR VPWR _08252_ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_475 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17679_ _07109_ _07665_ VGND VGND VPWR VPWR _08177_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_692 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_219 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_127_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_876 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_143_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_131_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09935_ _08735_ _08789_ VGND VGND VPWR VPWR _08800_ sky130_fd_sc_hd__xnor2_1
XTAP_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09866_ cla_inst.in1\[19\] VGND VGND VPWR VPWR _08049_ sky130_fd_sc_hd__clkbuf_4
XTAP_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09797_ _07265_ _07286_ VGND VGND VPWR VPWR _07297_ sky130_fd_sc_hd__nand2_2
XTAP_2504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10710_ _05235_ _05878_ VGND VGND VPWR VPWR _00803_ sky130_fd_sc_hd__nand2_1
XTAP_1847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11690_ _01741_ _01756_ _01781_ _01782_ VGND VGND VPWR VPWR _01783_ sky130_fd_sc_hd__a211o_1
XTAP_1869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_512 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10641_ _00723_ _00524_ _00732_ VGND VGND VPWR VPWR _00734_ sky130_fd_sc_hd__and3_1
XFILLER_0_76_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13360_ _00184_ _00174_ _03815_ _03914_ VGND VGND VPWR VPWR _03474_ sky130_fd_sc_hd__and4_1
XFILLER_0_106_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10572_ _00513_ VGND VGND VPWR VPWR _00665_ sky130_fd_sc_hd__buf_4
XFILLER_0_8_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_282 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12311_ _02334_ _02403_ VGND VGND VPWR VPWR _02404_ sky130_fd_sc_hd__nor2_1
XFILLER_0_23_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13291_ _04515_ _04438_ _00308_ _06689_ VGND VGND VPWR VPWR _03398_ sky130_fd_sc_hd__nand4_2
XFILLER_0_133_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15030_ _05188_ _05206_ _05298_ VGND VGND VPWR VPWR _05299_ sky130_fd_sc_hd__and3_1
XFILLER_0_133_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12242_ _07613_ _02205_ _02334_ VGND VGND VPWR VPWR _02335_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_20_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_121_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12173_ _02235_ _02238_ VGND VGND VPWR VPWR _02266_ sky130_fd_sc_hd__and2b_1
XFILLER_0_102_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11124_ _01132_ _01205_ _01216_ VGND VGND VPWR VPWR _01217_ sky130_fd_sc_hd__and3_1
X_16981_ _06816_ _06880_ _06944_ _07115_ VGND VGND VPWR VPWR _07416_ sky130_fd_sc_hd__or4_1
X_18720_ net58 _03155_ _09182_ VGND VGND VPWR VPWR _09246_ sky130_fd_sc_hd__mux2_1
X_11055_ _01079_ _01146_ _01145_ VGND VGND VPWR VPWR _01148_ sky130_fd_sc_hd__a21o_1
X_15932_ _06273_ _06276_ VGND VGND VPWR VPWR _06278_ sky130_fd_sc_hd__or2_1
X_10006_ cla_inst.in2\[26\] VGND VGND VPWR VPWR _09349_ sky130_fd_sc_hd__buf_2
X_15863_ _06153_ _06157_ _06158_ VGND VGND VPWR VPWR _06204_ sky130_fd_sc_hd__or3_1
X_18651_ net61 _03166_ _09193_ VGND VGND VPWR VPWR _09196_ sky130_fd_sc_hd__mux2_1
X_14814_ _05014_ _05015_ _05062_ VGND VGND VPWR VPWR _05064_ sky130_fd_sc_hd__a21o_1
X_17602_ _07630_ _07516_ _07982_ _07980_ VGND VGND VPWR VPWR _08094_ sky130_fd_sc_hd__o31a_1
X_15794_ _06128_ _06129_ VGND VGND VPWR VPWR _06130_ sky130_fd_sc_hd__nand2_1
X_18582_ _09127_ VGND VGND VPWR VPWR _09146_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_98_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14745_ _02200_ _03153_ _04846_ VGND VGND VPWR VPWR _04988_ sky130_fd_sc_hd__and3_1
XFILLER_0_58_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17533_ _08016_ _08018_ _06649_ VGND VGND VPWR VPWR _08019_ sky130_fd_sc_hd__o21ai_1
X_11957_ _02043_ _02047_ _02048_ _02049_ VGND VGND VPWR VPWR _02050_ sky130_fd_sc_hd__or4_4
XFILLER_0_129_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10908_ _05399_ _05355_ _04449_ _04471_ VGND VGND VPWR VPWR _01001_ sky130_fd_sc_hd__and4_1
X_17464_ _06764_ _07593_ VGND VGND VPWR VPWR _07943_ sky130_fd_sc_hd__nor2_1
X_14676_ _04911_ _04912_ VGND VGND VPWR VPWR _04913_ sky130_fd_sc_hd__or2_1
XFILLER_0_46_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11888_ _01971_ _01973_ VGND VGND VPWR VPWR _01981_ sky130_fd_sc_hd__nor2_1
XFILLER_0_73_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16415_ _06578_ _06764_ VGND VGND VPWR VPWR _06801_ sky130_fd_sc_hd__or2_1
X_13627_ _03990_ _00308_ VGND VGND VPWR VPWR _03766_ sky130_fd_sc_hd__nand2_1
X_10839_ _00916_ _00914_ _00915_ VGND VGND VPWR VPWR _00932_ sky130_fd_sc_hd__nand3_1
X_17395_ _07207_ _07751_ net146 _06947_ VGND VGND VPWR VPWR _07868_ sky130_fd_sc_hd__a22o_1
XFILLER_0_6_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16346_ _03049_ _06609_ _06725_ _06467_ VGND VGND VPWR VPWR _06726_ sky130_fd_sc_hd__o211a_1
XFILLER_0_54_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13558_ _03690_ _03482_ VGND VGND VPWR VPWR _03691_ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12509_ _02553_ _02600_ _02599_ VGND VGND VPWR VPWR _02602_ sky130_fd_sc_hd__nand3_1
X_16277_ _00218_ _06568_ _06650_ _03313_ VGND VGND VPWR VPWR _06651_ sky130_fd_sc_hd__o22a_4
XFILLER_0_113_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13489_ _03610_ _03613_ _03614_ VGND VGND VPWR VPWR _03615_ sky130_fd_sc_hd__and3_1
XFILLER_0_2_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_112_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15228_ _05512_ _05514_ VGND VGND VPWR VPWR _05515_ sky130_fd_sc_hd__xnor2_1
X_18016_ _08541_ _08542_ _08543_ VGND VGND VPWR VPWR _08544_ sky130_fd_sc_hd__or3_1
XFILLER_0_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15159_ _05437_ _05438_ VGND VGND VPWR VPWR _05439_ sky130_fd_sc_hd__and2_1
XFILLER_0_22_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09720_ _05017_ VGND VGND VPWR VPWR _06460_ sky130_fd_sc_hd__buf_6
X_18918_ clknet_4_11_0_clk _00072_ VGND VGND VPWR VPWR ApproximateM_inst.lob_16.lob2.genblk1\[4\].genblk1.mux.sel
+ sky130_fd_sc_hd__dfxtp_2
X_09651_ _05704_ VGND VGND VPWR VPWR _05715_ sky130_fd_sc_hd__clkbuf_8
X_18849_ clknet_4_6_0_clk net294 VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__dfxtp_1
X_09582_ _03946_ _03957_ _03706_ VGND VGND VPWR VPWR _04962_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_96_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_355 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_712 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_740 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_130_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold140 net104 VGND VGND VPWR VPWR net303 sky130_fd_sc_hd__dlygate4sd3_1
Xhold151 net106 VGND VGND VPWR VPWR net314 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09918_ _06460_ VGND VGND VPWR VPWR _08615_ sky130_fd_sc_hd__buf_6
X_09849_ _07853_ _07744_ _07766_ VGND VGND VPWR VPWR _07864_ sky130_fd_sc_hd__a21o_1
X_12860_ _00900_ _00903_ _00902_ VGND VGND VPWR VPWR _02953_ sky130_fd_sc_hd__o21a_1
XTAP_2301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11811_ _01897_ _01898_ _01876_ VGND VGND VPWR VPWR _01904_ sky130_fd_sc_hd__a21oi_1
XTAP_2334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12791_ _01450_ _02883_ VGND VGND VPWR VPWR _02884_ sky130_fd_sc_hd__nand2_2
XTAP_2345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14530_ _04603_ _04752_ VGND VGND VPWR VPWR _04753_ sky130_fd_sc_hd__xnor2_1
XTAP_1633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11742_ _01833_ _01834_ VGND VGND VPWR VPWR _01835_ sky130_fd_sc_hd__xnor2_1
XTAP_2389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14461_ _04566_ _04538_ _04676_ _04677_ VGND VGND VPWR VPWR _04678_ sky130_fd_sc_hd__o211a_1
XTAP_1688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11673_ _01764_ _01765_ VGND VGND VPWR VPWR _01766_ sky130_fd_sc_hd__or2_1
XTAP_1699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_331 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16200_ _06564_ _06566_ _03313_ VGND VGND VPWR VPWR _06567_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_37_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13412_ _03355_ _03362_ _03529_ _03530_ _02969_ VGND VGND VPWR VPWR _03532_ sky130_fd_sc_hd__a311o_1
X_10624_ _00163_ _00716_ VGND VGND VPWR VPWR _00717_ sky130_fd_sc_hd__nand2_1
X_17180_ _07042_ _07303_ _07130_ _07302_ VGND VGND VPWR VPWR _07633_ sky130_fd_sc_hd__o22a_1
X_14392_ _04600_ _04601_ _04304_ VGND VGND VPWR VPWR _04603_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_70_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16131_ _06467_ _06491_ VGND VGND VPWR VPWR _06492_ sky130_fd_sc_hd__nand2_1
X_13343_ _03455_ VGND VGND VPWR VPWR _03456_ sky130_fd_sc_hd__buf_4
X_10555_ _05453_ _00645_ _06732_ _05715_ VGND VGND VPWR VPWR _00648_ sky130_fd_sc_hd__nand4_2
XFILLER_0_122_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16062_ op_code\[3\] op_code\[2\] VGND VGND VPWR VPWR _06418_ sky130_fd_sc_hd__nand2b_2
X_13274_ _01521_ _05050_ net240 _03378_ VGND VGND VPWR VPWR _03380_ sky130_fd_sc_hd__nand4_1
X_10486_ _00577_ _00576_ _00373_ _00370_ VGND VGND VPWR VPWR _00579_ sky130_fd_sc_hd__o211a_1
XFILLER_0_121_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15013_ _05278_ _05280_ VGND VGND VPWR VPWR _05281_ sky130_fd_sc_hd__xor2_2
X_12225_ _02315_ _02316_ _02302_ _02314_ VGND VGND VPWR VPWR _02318_ sky130_fd_sc_hd__a211oi_2
X_12156_ _02233_ _02232_ VGND VGND VPWR VPWR _02249_ sky130_fd_sc_hd__and2b_1
X_11107_ _01179_ _01180_ _01166_ _01178_ VGND VGND VPWR VPWR _01200_ sky130_fd_sc_hd__a211o_1
X_12087_ _05301_ _00130_ _09212_ _05279_ VGND VGND VPWR VPWR _02180_ sky130_fd_sc_hd__a22o_1
X_16964_ _07393_ _07397_ VGND VGND VPWR VPWR _07398_ sky130_fd_sc_hd__nand2_1
X_18703_ net51 _09190_ _09233_ VGND VGND VPWR VPWR _00060_ sky130_fd_sc_hd__o21a_1
X_11038_ _01096_ _01125_ _01124_ VGND VGND VPWR VPWR _01131_ sky130_fd_sc_hd__a21o_1
X_15915_ _06258_ _06259_ VGND VGND VPWR VPWR _06260_ sky130_fd_sc_hd__nand2_1
X_16895_ _07310_ _07321_ VGND VGND VPWR VPWR _07323_ sky130_fd_sc_hd__nand2_1
X_18634_ _09181_ VGND VGND VPWR VPWR _09182_ sky130_fd_sc_hd__clkbuf_4
X_15846_ _06076_ _06079_ _06185_ VGND VGND VPWR VPWR _06186_ sky130_fd_sc_hd__a21o_1
X_18565_ net250 _09098_ _09133_ _09126_ VGND VGND VPWR VPWR _00008_ sky130_fd_sc_hd__o211a_1
X_15777_ _06032_ _06110_ VGND VGND VPWR VPWR _06111_ sky130_fd_sc_hd__and2_1
X_12989_ _03063_ _03078_ _03081_ VGND VGND VPWR VPWR _03082_ sky130_fd_sc_hd__mux2_2
XFILLER_0_87_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17516_ _07856_ _07857_ _07874_ VGND VGND VPWR VPWR _08000_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_129_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14728_ _04730_ _04833_ _04862_ _04863_ VGND VGND VPWR VPWR _04969_ sky130_fd_sc_hd__a211oi_4
X_18496_ _03011_ _06920_ _06921_ VGND VGND VPWR VPWR _09064_ sky130_fd_sc_hd__a21o_1
X_14659_ _00877_ _01112_ VGND VGND VPWR VPWR _04894_ sky130_fd_sc_hd__nand2_1
X_17447_ _06376_ _06375_ _06372_ VGND VGND VPWR VPWR _07925_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_27_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17378_ _07841_ _07848_ VGND VGND VPWR VPWR _07849_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_42_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_632 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16329_ _01677_ _02370_ _03175_ VGND VGND VPWR VPWR _06708_ sky130_fd_sc_hd__or3_1
XFILLER_0_42_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_6 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09703_ _04984_ _04700_ VGND VGND VPWR VPWR _06277_ sky130_fd_sc_hd__nand2_4
XFILLER_0_4_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09634_ _05235_ _05486_ _05475_ _05519_ VGND VGND VPWR VPWR _05529_ sky130_fd_sc_hd__nand4_2
X_09565_ _03356_ _03377_ _03914_ _03476_ VGND VGND VPWR VPWR _04777_ sky130_fd_sc_hd__nand4_1
XFILLER_0_78_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09496_ _04001_ _04012_ VGND VGND VPWR VPWR _04023_ sky130_fd_sc_hd__nand2_8
XFILLER_0_148_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_147_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_147_185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_135_358 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_104_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_144_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10340_ _03465_ _04395_ VGND VGND VPWR VPWR _00433_ sky130_fd_sc_hd__and2_1
XFILLER_0_103_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_116_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10271_ _00361_ _00363_ VGND VGND VPWR VPWR _00364_ sky130_fd_sc_hd__xor2_1
XFILLER_0_103_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12010_ _02098_ _02101_ _02102_ VGND VGND VPWR VPWR _02103_ sky130_fd_sc_hd__a21boi_1
X_13961_ _05453_ _09248_ _04130_ VGND VGND VPWR VPWR _04131_ sky130_fd_sc_hd__a21boi_1
X_12912_ cla_inst.in2\[31\] VGND VGND VPWR VPWR _03005_ sky130_fd_sc_hd__clkbuf_4
X_15700_ _06025_ _06026_ VGND VGND VPWR VPWR _06027_ sky130_fd_sc_hd__nor2_1
X_16680_ _07086_ _07088_ _04247_ VGND VGND VPWR VPWR _07089_ sky130_fd_sc_hd__mux2_2
X_13892_ _04052_ _04053_ _04054_ VGND VGND VPWR VPWR _04057_ sky130_fd_sc_hd__o21ai_1
X_12843_ _02933_ _02934_ _02935_ _02913_ VGND VGND VPWR VPWR _02936_ sky130_fd_sc_hd__o211a_1
X_15631_ _05947_ _05951_ _05952_ VGND VGND VPWR VPWR _05953_ sky130_fd_sc_hd__a21oi_2
XTAP_2120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15562_ _05875_ _05877_ _03202_ VGND VGND VPWR VPWR _05879_ sky130_fd_sc_hd__o21ai_1
XTAP_2164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18350_ _08903_ _08905_ VGND VGND VPWR VPWR _08906_ sky130_fd_sc_hd__or2_1
XTAP_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12774_ _01806_ VGND VGND VPWR VPWR _02867_ sky130_fd_sc_hd__inv_2
XTAP_2175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14513_ _04723_ _04724_ _04734_ VGND VGND VPWR VPWR _04735_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_68_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17301_ _07738_ _07764_ VGND VGND VPWR VPWR _07765_ sky130_fd_sc_hd__xnor2_1
XTAP_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11725_ _00146_ _01537_ _01536_ VGND VGND VPWR VPWR _01818_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_138_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18281_ _03056_ _06463_ _08831_ VGND VGND VPWR VPWR _09403_ sky130_fd_sc_hd__a21oi_2
X_15493_ _05087_ VGND VGND VPWR VPWR _05803_ sky130_fd_sc_hd__inv_2
XFILLER_0_154_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14444_ _04658_ _04659_ VGND VGND VPWR VPWR _04660_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_71_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17232_ _04725_ _06920_ _06921_ VGND VGND VPWR VPWR _07691_ sky130_fd_sc_hd__a21o_1
XFILLER_0_154_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11656_ _01744_ _01747_ _01698_ VGND VGND VPWR VPWR _01749_ sky130_fd_sc_hd__o21ai_1
X_10607_ _00568_ _00569_ VGND VGND VPWR VPWR _00700_ sky130_fd_sc_hd__nand2_1
X_17163_ _07606_ _07614_ VGND VGND VPWR VPWR _07615_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_154_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14375_ _04581_ _04582_ _04583_ VGND VGND VPWR VPWR _04584_ sky130_fd_sc_hd__and3_4
XFILLER_0_107_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11587_ _01673_ _01675_ VGND VGND VPWR VPWR _01680_ sky130_fd_sc_hd__and2_1
X_16114_ _06469_ _06473_ _03099_ VGND VGND VPWR VPWR _06474_ sky130_fd_sc_hd__mux2_1
X_13326_ _03286_ _03287_ _03436_ VGND VGND VPWR VPWR _03437_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_12_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10538_ _00622_ _00630_ VGND VGND VPWR VPWR _00631_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_101_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17094_ _07411_ _07414_ _07412_ VGND VGND VPWR VPWR _07540_ sky130_fd_sc_hd__o21a_1
X_16045_ _02994_ _04900_ VGND VGND VPWR VPWR _06399_ sky130_fd_sc_hd__or2_1
X_13257_ _03358_ _03361_ VGND VGND VPWR VPWR _03362_ sky130_fd_sc_hd__nand2_1
X_10469_ _00203_ _00399_ VGND VGND VPWR VPWR _00562_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12208_ _02134_ _02149_ _02150_ _02300_ VGND VGND VPWR VPWR _02301_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_86_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13188_ _03286_ _03287_ VGND VGND VPWR VPWR _03288_ sky130_fd_sc_hd__xor2_2
XFILLER_0_19_20 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12139_ _07243_ _00949_ _03421_ _07221_ VGND VGND VPWR VPWR _02232_ sky130_fd_sc_hd__a22o_1
X_17996_ _03000_ _06593_ _06594_ VGND VGND VPWR VPWR _08523_ sky130_fd_sc_hd__a21oi_1
X_16947_ _07339_ _07340_ VGND VGND VPWR VPWR _07379_ sky130_fd_sc_hd__nand2_1
XFILLER_0_35_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16878_ _06816_ _07302_ _07303_ _06764_ VGND VGND VPWR VPWR _07304_ sky130_fd_sc_hd__o22a_1
X_18617_ net263 _09157_ _09169_ _09162_ VGND VGND VPWR VPWR _00029_ sky130_fd_sc_hd__o211a_1
X_15829_ _06104_ _06108_ _06166_ VGND VGND VPWR VPWR _06167_ sky130_fd_sc_hd__a21o_1
X_18548_ net28 _09109_ VGND VGND VPWR VPWR _09119_ sky130_fd_sc_hd__or2_1
X_18479_ _09036_ _09008_ _09043_ VGND VGND VPWR VPWR _09045_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_118_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_542 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_141_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09617_ _05279_ _05301_ _05322_ _05333_ VGND VGND VPWR VPWR _05344_ sky130_fd_sc_hd__and4_1
XFILLER_0_97_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09548_ _04580_ VGND VGND VPWR VPWR _04591_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_38_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09479_ _03826_ VGND VGND VPWR VPWR _03837_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_136_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_256 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_779 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11510_ _01562_ _01563_ _01525_ _01540_ VGND VGND VPWR VPWR _01603_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_93_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12490_ _02580_ _02582_ VGND VGND VPWR VPWR _02583_ sky130_fd_sc_hd__nor2_1
X_11441_ _01529_ _01532_ _01530_ VGND VGND VPWR VPWR _01534_ sky130_fd_sc_hd__and3_1
XFILLER_0_34_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire136 _03205_ VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__buf_1
XFILLER_0_80_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14160_ _04347_ _04348_ VGND VGND VPWR VPWR _04349_ sky130_fd_sc_hd__nand2_1
X_11372_ _01382_ _01392_ _00821_ _01463_ VGND VGND VPWR VPWR _01465_ sky130_fd_sc_hd__a211o_2
XFILLER_0_150_158 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13111_ _00620_ _00621_ _00631_ VGND VGND VPWR VPWR _03205_ sky130_fd_sc_hd__nor3_1
X_10323_ _00396_ _00397_ _00415_ VGND VGND VPWR VPWR _00416_ sky130_fd_sc_hd__a21oi_1
X_14091_ net173 _04095_ _04271_ _04272_ VGND VGND VPWR VPWR _04273_ sky130_fd_sc_hd__o211a_1
XFILLER_0_104_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13042_ _03028_ _01692_ VGND VGND VPWR VPWR _03134_ sky130_fd_sc_hd__nor2_1
X_10254_ _00341_ _00346_ VGND VGND VPWR VPWR _00347_ sky130_fd_sc_hd__xor2_1
XFILLER_0_30_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17850_ _08349_ _08350_ _08362_ VGND VGND VPWR VPWR _08363_ sky130_fd_sc_hd__a21o_1
X_10185_ _00275_ _00276_ _00277_ VGND VGND VPWR VPWR _00278_ sky130_fd_sc_hd__nand3_1
XFILLER_0_56_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16801_ _07217_ _07219_ VGND VGND VPWR VPWR _07220_ sky130_fd_sc_hd__nand2_1
X_17781_ _08279_ _08286_ VGND VGND VPWR VPWR _08288_ sky130_fd_sc_hd__nor2_1
X_14993_ _05256_ _05258_ VGND VGND VPWR VPWR _05259_ sky130_fd_sc_hd__xnor2_1
X_16732_ _07142_ _07144_ VGND VGND VPWR VPWR _07146_ sky130_fd_sc_hd__or2_1
X_13944_ _04111_ _04112_ _04548_ _07722_ VGND VGND VPWR VPWR _04113_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_89_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13875_ _04029_ _04037_ VGND VGND VPWR VPWR _04038_ sky130_fd_sc_hd__xnor2_2
X_16663_ _07068_ _07070_ VGND VGND VPWR VPWR _07071_ sky130_fd_sc_hd__xor2_1
X_18402_ _08907_ _08946_ _08960_ VGND VGND VPWR VPWR _08963_ sky130_fd_sc_hd__and3_1
X_15614_ _05846_ VGND VGND VPWR VPWR _05935_ sky130_fd_sc_hd__inv_2
X_12826_ _02916_ _02917_ VGND VGND VPWR VPWR _02919_ sky130_fd_sc_hd__nand2_1
X_16594_ _06343_ _06345_ _06995_ VGND VGND VPWR VPWR _06996_ sky130_fd_sc_hd__a21o_1
X_18333_ _08888_ _06403_ _06402_ VGND VGND VPWR VPWR _08889_ sky130_fd_sc_hd__a21oi_1
X_15545_ _05858_ _05846_ _05847_ VGND VGND VPWR VPWR _05860_ sky130_fd_sc_hd__and3_1
XTAP_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12757_ _02330_ _02849_ VGND VGND VPWR VPWR _02850_ sky130_fd_sc_hd__nor2_1
XTAP_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11708_ _01790_ _01799_ _01798_ VGND VGND VPWR VPWR _01801_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_16_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15476_ _05665_ _05668_ _05783_ VGND VGND VPWR VPWR _05785_ sky130_fd_sc_hd__or3_1
X_18264_ _03055_ _06511_ _01359_ VGND VGND VPWR VPWR _08814_ sky130_fd_sc_hd__and3b_1
X_12688_ _06993_ _07646_ _02779_ _02780_ VGND VGND VPWR VPWR _02781_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_154_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14427_ _04630_ _04640_ VGND VGND VPWR VPWR _04641_ sky130_fd_sc_hd__nor2_1
X_17215_ _07671_ _07558_ VGND VGND VPWR VPWR _07672_ sky130_fd_sc_hd__nor2_1
XFILLER_0_154_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11639_ _01730_ _01726_ _01725_ VGND VGND VPWR VPWR _01732_ sky130_fd_sc_hd__and3b_1
XFILLER_0_114_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_166 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_108_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18195_ _08696_ _08738_ VGND VGND VPWR VPWR _08739_ sky130_fd_sc_hd__nor2_1
XFILLER_0_141_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14358_ _04425_ _04382_ _04540_ _04541_ VGND VGND VPWR VPWR _04565_ sky130_fd_sc_hd__a211o_1
XFILLER_0_107_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17146_ _07595_ VGND VGND VPWR VPWR _07596_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_24_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13309_ _05410_ _05301_ _07004_ _07102_ VGND VGND VPWR VPWR _03418_ sky130_fd_sc_hd__nand4_2
XFILLER_0_141_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17077_ _07519_ _07520_ VGND VGND VPWR VPWR _07521_ sky130_fd_sc_hd__nand2_1
X_14289_ _04487_ _04488_ _04315_ _04331_ VGND VGND VPWR VPWR _04490_ sky130_fd_sc_hd__a211o_1
XFILLER_0_123_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16028_ _06377_ _06378_ _06379_ VGND VGND VPWR VPWR _06380_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_110_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17979_ _08502_ _08503_ VGND VGND VPWR VPWR _08504_ sky130_fd_sc_hd__and2_1
XFILLER_0_149_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold88 _00008_ VGND VGND VPWR VPWR net251 sky130_fd_sc_hd__dlygate4sd3_1
X_11990_ _02003_ _02082_ VGND VGND VPWR VPWR _02083_ sky130_fd_sc_hd__xor2_1
Xhold99 _00010_ VGND VGND VPWR VPWR net262 sky130_fd_sc_hd__dlygate4sd3_1
X_10941_ _03531_ _03509_ _00130_ _07548_ VGND VGND VPWR VPWR _01034_ sky130_fd_sc_hd__nand4_2
X_13660_ _03794_ _03800_ _03801_ VGND VGND VPWR VPWR _03802_ sky130_fd_sc_hd__nand3_1
XFILLER_0_97_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10872_ _00963_ _00964_ VGND VGND VPWR VPWR _00965_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_85_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12611_ _02701_ _02702_ _02703_ VGND VGND VPWR VPWR _02704_ sky130_fd_sc_hd__nand3_1
XFILLER_0_38_223 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13591_ _03724_ _03725_ _03726_ VGND VGND VPWR VPWR _03727_ sky130_fd_sc_hd__or3_1
XFILLER_0_94_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_623 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15330_ _05624_ VGND VGND VPWR VPWR _05625_ sky130_fd_sc_hd__inv_2
X_12542_ _02602_ _02598_ _02601_ VGND VGND VPWR VPWR _02635_ sky130_fd_sc_hd__nand3_1
XFILLER_0_94_896 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_108_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15261_ _05526_ _05527_ _05548_ VGND VGND VPWR VPWR _05550_ sky130_fd_sc_hd__or3_1
X_12473_ _02544_ _02557_ _02565_ VGND VGND VPWR VPWR _02566_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_136_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_151_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14212_ _04233_ _04235_ _04065_ VGND VGND VPWR VPWR _04407_ sky130_fd_sc_hd__o21bai_1
X_17000_ _07435_ _07436_ VGND VGND VPWR VPWR _07437_ sky130_fd_sc_hd__xnor2_1
X_11424_ _04984_ _00181_ VGND VGND VPWR VPWR _01517_ sky130_fd_sc_hd__nand2_1
XFILLER_0_151_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15192_ _05350_ _05358_ _05474_ VGND VGND VPWR VPWR _05476_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_123_136 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_151_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_8 _00461_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_61_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_123 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14143_ _04315_ _04316_ _04328_ VGND VGND VPWR VPWR _04331_ sky130_fd_sc_hd__nor3_2
X_11355_ _01352_ _01354_ _01351_ VGND VGND VPWR VPWR _01448_ sky130_fd_sc_hd__o21ba_2
XFILLER_0_104_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10306_ _00398_ VGND VGND VPWR VPWR _00399_ sky130_fd_sc_hd__clkbuf_8
X_18951_ clknet_4_1_0_clk _09412_ VGND VGND VPWR VPWR salida\[4\] sky130_fd_sc_hd__dfxtp_1
X_14074_ _03080_ _02981_ _03560_ VGND VGND VPWR VPWR _04255_ sky130_fd_sc_hd__or3_1
X_11286_ _01290_ _01308_ _01309_ VGND VGND VPWR VPWR _01379_ sky130_fd_sc_hd__nor3_1
XTAP_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17902_ _06559_ _08419_ VGND VGND VPWR VPWR _08421_ sky130_fd_sc_hd__or2_1
XTAP_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13025_ _03082_ _03116_ _03117_ VGND VGND VPWR VPWR _03118_ sky130_fd_sc_hd__mux2_1
X_10237_ _00326_ _00327_ _00329_ VGND VGND VPWR VPWR _00330_ sky130_fd_sc_hd__a21o_1
X_18882_ clknet_4_9_0_clk _00036_ VGND VGND VPWR VPWR ApproximateM_inst.lob_16.lob1.mux.sel
+ sky130_fd_sc_hd__dfxtp_1
X_17833_ _06649_ _08327_ _08328_ _08345_ VGND VGND VPWR VPWR _08346_ sky130_fd_sc_hd__a31o_1
X_10168_ _00252_ _00260_ VGND VGND VPWR VPWR _00261_ sky130_fd_sc_hd__xnor2_1
X_17764_ _08268_ _08269_ VGND VGND VPWR VPWR _08270_ sky130_fd_sc_hd__nand2_1
X_14976_ _05228_ _05239_ VGND VGND VPWR VPWR _05240_ sky130_fd_sc_hd__xnor2_2
X_10099_ _00191_ VGND VGND VPWR VPWR _00192_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_89_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16715_ _07124_ _06816_ _07126_ net237 VGND VGND VPWR VPWR _07127_ sky130_fd_sc_hd__o22a_1
X_13927_ _03345_ net172 cla_inst.in1\[22\] cla_inst.in1\[20\] VGND VGND VPWR VPWR
+ _04094_ sky130_fd_sc_hd__and4_1
X_17695_ _08090_ _08091_ _08088_ VGND VGND VPWR VPWR _08195_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_89_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16646_ _06952_ _06958_ _07051_ VGND VGND VPWR VPWR _07052_ sky130_fd_sc_hd__o21ai_1
X_13858_ _03843_ _03844_ VGND VGND VPWR VPWR _04019_ sky130_fd_sc_hd__or2b_1
XFILLER_0_29_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12809_ _01458_ _01460_ _02900_ VGND VGND VPWR VPWR _02902_ sky130_fd_sc_hd__nor3_1
X_16577_ _06867_ _06887_ VGND VGND VPWR VPWR _06977_ sky130_fd_sc_hd__or2b_1
X_13789_ _03728_ _07962_ VGND VGND VPWR VPWR _03943_ sky130_fd_sc_hd__nand2_1
XFILLER_0_45_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18316_ _08868_ _08869_ VGND VGND VPWR VPWR _08870_ sky130_fd_sc_hd__or2_1
XFILLER_0_17_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15528_ _05831_ _05749_ _05840_ VGND VGND VPWR VPWR _05841_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_32_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18247_ _08712_ _08726_ _08793_ VGND VGND VPWR VPWR _08795_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_142_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15459_ _05763_ _05765_ VGND VGND VPWR VPWR _05766_ sky130_fd_sc_hd__or2_1
XFILLER_0_4_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18178_ _08620_ _08622_ _08719_ VGND VGND VPWR VPWR _08720_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_12_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17129_ _07577_ _06845_ _02979_ VGND VGND VPWR VPWR _07578_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09951_ _08930_ _08941_ _08951_ _08962_ VGND VGND VPWR VPWR _08973_ sky130_fd_sc_hd__a211o_1
XFILLER_0_111_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09882_ _08169_ VGND VGND VPWR VPWR _08224_ sky130_fd_sc_hd__buf_6
XTAP_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_811 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_442 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11140_ _01218_ _01228_ _01231_ _01232_ VGND VGND VPWR VPWR _01233_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_101_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11071_ _01157_ _01158_ _01162_ VGND VGND VPWR VPWR _01164_ sky130_fd_sc_hd__nand3_1
XFILLER_0_101_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput78 net78 VGND VGND VPWR VPWR leds[6] sky130_fd_sc_hd__buf_2
Xoutput89 net89 VGND VGND VPWR VPWR o_wb_data[15] sky130_fd_sc_hd__clkbuf_4
X_10022_ _00107_ VGND VGND VPWR VPWR _00115_ sky130_fd_sc_hd__buf_4
X_14830_ _05077_ _05079_ _03202_ VGND VGND VPWR VPWR _05081_ sky130_fd_sc_hd__o21a_1
XFILLER_0_98_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14761_ _05003_ VGND VGND VPWR VPWR _05005_ sky130_fd_sc_hd__inv_2
X_11973_ _02061_ _02062_ _02065_ VGND VGND VPWR VPWR _02066_ sky130_fd_sc_hd__a21bo_1
X_16500_ _06527_ _06809_ _06891_ _06892_ VGND VGND VPWR VPWR _06893_ sky130_fd_sc_hd__a31o_1
X_13712_ _03702_ _03708_ VGND VGND VPWR VPWR _03860_ sky130_fd_sc_hd__nand2_1
X_10924_ _01014_ _01015_ _00989_ _00997_ VGND VGND VPWR VPWR _01017_ sky130_fd_sc_hd__a211o_1
X_14692_ _04928_ _04929_ VGND VGND VPWR VPWR _04931_ sky130_fd_sc_hd__or2_1
X_17480_ _07106_ _07332_ VGND VGND VPWR VPWR _07960_ sky130_fd_sc_hd__nor2_1
XFILLER_0_67_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16431_ _06809_ _06817_ VGND VGND VPWR VPWR _06818_ sky130_fd_sc_hd__xor2_1
XFILLER_0_129_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13643_ net329 _03773_ _03783_ VGND VGND VPWR VPWR _03784_ sky130_fd_sc_hd__o21ai_2
X_10855_ _00942_ _00947_ VGND VGND VPWR VPWR _00948_ sky130_fd_sc_hd__xor2_1
XFILLER_0_67_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13574_ _03702_ _03708_ VGND VGND VPWR VPWR _03709_ sky130_fd_sc_hd__xor2_1
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16362_ _03164_ _06742_ VGND VGND VPWR VPWR _06744_ sky130_fd_sc_hd__nand2_1
X_10786_ _00870_ _00875_ VGND VGND VPWR VPWR _00879_ sky130_fd_sc_hd__xnor2_1
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18101_ _07390_ _07650_ _08535_ _08534_ VGND VGND VPWR VPWR _08636_ sky130_fd_sc_hd__a31o_1
X_15313_ _05491_ _05493_ VGND VGND VPWR VPWR _05608_ sky130_fd_sc_hd__or2b_1
X_12525_ _02616_ _02617_ VGND VGND VPWR VPWR _02618_ sky130_fd_sc_hd__nand2_1
XFILLER_0_81_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16293_ _06659_ _06668_ VGND VGND VPWR VPWR _06669_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18032_ _08559_ _08560_ VGND VGND VPWR VPWR _08562_ sky130_fd_sc_hd__and2_1
X_15244_ _05528_ _05531_ VGND VGND VPWR VPWR _05532_ sky130_fd_sc_hd__xnor2_1
X_12456_ _00832_ _00171_ _02494_ _02493_ VGND VGND VPWR VPWR _02549_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11407_ _01430_ _01498_ _01496_ _01497_ VGND VGND VPWR VPWR _01500_ sky130_fd_sc_hd__a211oi_2
X_15175_ _05430_ _05342_ _05456_ VGND VGND VPWR VPWR _05457_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_111_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12387_ _02360_ _02408_ _02406_ VGND VGND VPWR VPWR _02480_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_105_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14126_ _04301_ _04311_ VGND VGND VPWR VPWR _04312_ sky130_fd_sc_hd__xnor2_1
X_11338_ _01429_ _01347_ _01423_ VGND VGND VPWR VPWR _01431_ sky130_fd_sc_hd__or3_1
X_18934_ clknet_4_8_0_clk _00088_ VGND VGND VPWR VPWR cla_inst.in2\[20\] sky130_fd_sc_hd__dfxtp_2
X_14057_ _04065_ _04072_ _04236_ VGND VGND VPWR VPWR _04237_ sky130_fd_sc_hd__a21oi_1
X_11269_ _01355_ _01361_ VGND VGND VPWR VPWR _01362_ sky130_fd_sc_hd__nor2_1
X_13008_ _00248_ VGND VGND VPWR VPWR _03101_ sky130_fd_sc_hd__clkbuf_4
X_18865_ clknet_4_4_0_clk net268 VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__dfxtp_1
X_17816_ _08252_ _08223_ _08326_ VGND VGND VPWR VPWR _08327_ sky130_fd_sc_hd__a21o_1
X_18796_ _09306_ VGND VGND VPWR VPWR _00089_ sky130_fd_sc_hd__clkbuf_1
X_17747_ _08249_ _02329_ _08227_ _08250_ _02969_ VGND VGND VPWR VPWR _08251_ sky130_fd_sc_hd__a311oi_2
X_14959_ _05219_ _05220_ VGND VGND VPWR VPWR _05221_ sky130_fd_sc_hd__xor2_1
XFILLER_0_89_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17678_ _08174_ _08175_ VGND VGND VPWR VPWR _08176_ sky130_fd_sc_hd__nand2_1
X_16629_ _00398_ _07032_ VGND VGND VPWR VPWR _07033_ sky130_fd_sc_hd__nor2_1
XFILLER_0_85_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_143_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09934_ _08768_ _08778_ VGND VGND VPWR VPWR _08789_ sky130_fd_sc_hd__and2b_1
XFILLER_0_110_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09865_ ApproximateM_inst.lob_16.lob2.genblk1\[6\].genblk1.mux.sel VGND VGND VPWR
+ VPWR _08039_ sky130_fd_sc_hd__clkbuf_4
XTAP_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09796_ _06982_ _07156_ _07265_ _07276_ VGND VGND VPWR VPWR _07286_ sky130_fd_sc_hd__nand4_2
XTAP_2505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10640_ _00723_ _00524_ _00732_ VGND VGND VPWR VPWR _00733_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_36_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10571_ _00496_ _00505_ VGND VGND VPWR VPWR _00664_ sky130_fd_sc_hd__nand2_1
XFILLER_0_63_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12310_ _05235_ _09219_ _02332_ _02333_ VGND VGND VPWR VPWR _02403_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_91_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_118_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13290_ _04438_ _05704_ _06689_ _04646_ VGND VGND VPWR VPWR _03397_ sky130_fd_sc_hd__a22o_1
XFILLER_0_51_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12241_ _08713_ _00127_ _02332_ _02333_ VGND VGND VPWR VPWR _02334_ sky130_fd_sc_hd__and4_1
XFILLER_0_121_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12172_ _02111_ _02119_ VGND VGND VPWR VPWR _02265_ sky130_fd_sc_hd__xnor2_1
X_11123_ _01209_ _01214_ _01215_ VGND VGND VPWR VPWR _01216_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_101_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16980_ _07413_ _07414_ VGND VGND VPWR VPWR _07415_ sky130_fd_sc_hd__xnor2_1
X_11054_ _01079_ _01145_ _01146_ VGND VGND VPWR VPWR _01147_ sky130_fd_sc_hd__nand3_2
X_15931_ _06274_ _06250_ _06275_ VGND VGND VPWR VPWR _06276_ sky130_fd_sc_hd__or3b_1
X_10005_ _06938_ _08311_ _09344_ _09347_ VGND VGND VPWR VPWR _09348_ sky130_fd_sc_hd__a211o_4
X_18650_ _09195_ VGND VGND VPWR VPWR _00039_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15862_ _06199_ _06201_ VGND VGND VPWR VPWR _06203_ sky130_fd_sc_hd__nor2_1
X_17601_ _08090_ _08091_ VGND VGND VPWR VPWR _08092_ sky130_fd_sc_hd__xor2_1
X_14813_ _05014_ _05015_ _05062_ VGND VGND VPWR VPWR _05063_ sky130_fd_sc_hd__nand3_2
XFILLER_0_99_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18581_ net306 _09140_ _09143_ _09144_ VGND VGND VPWR VPWR _00014_ sky130_fd_sc_hd__o211a_1
X_15793_ _06058_ _06087_ _06126_ VGND VGND VPWR VPWR _06129_ sky130_fd_sc_hd__nand3_1
XFILLER_0_99_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17532_ _07900_ _07903_ _07901_ VGND VGND VPWR VPWR _08018_ sky130_fd_sc_hd__o21ai_4
X_14744_ _04982_ _04983_ _04985_ VGND VGND VPWR VPWR _04987_ sky130_fd_sc_hd__a21o_1
XFILLER_0_99_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_284 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11956_ _01964_ _02046_ VGND VGND VPWR VPWR _02049_ sky130_fd_sc_hd__nor2_1
XFILLER_0_59_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10907_ _08713_ _04580_ VGND VGND VPWR VPWR _01000_ sky130_fd_sc_hd__nand2_1
X_17463_ _07938_ _07941_ VGND VGND VPWR VPWR _07942_ sky130_fd_sc_hd__xnor2_1
X_14675_ _00106_ _05486_ _04909_ _04910_ VGND VGND VPWR VPWR _04912_ sky130_fd_sc_hd__o2bb2a_1
X_11887_ _01979_ VGND VGND VPWR VPWR _01980_ sky130_fd_sc_hd__inv_2
XFILLER_0_39_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16414_ _06572_ _06756_ VGND VGND VPWR VPWR _06800_ sky130_fd_sc_hd__nor2_1
X_13626_ _06689_ _03763_ _03764_ VGND VGND VPWR VPWR _03765_ sky130_fd_sc_hd__a21bo_1
X_10838_ _00929_ _00930_ VGND VGND VPWR VPWR _00931_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_55_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17394_ _07302_ _07303_ _07126_ _07318_ VGND VGND VPWR VPWR _07867_ sky130_fd_sc_hd__or4_1
XFILLER_0_116_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16345_ _02982_ _06614_ VGND VGND VPWR VPWR _06725_ sky130_fd_sc_hd__or2_1
X_10769_ _07853_ _00318_ _00861_ VGND VGND VPWR VPWR _00862_ sky130_fd_sc_hd__and3_2
X_13557_ _03478_ _03479_ VGND VGND VPWR VPWR _03690_ sky130_fd_sc_hd__or2b_1
XFILLER_0_54_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12508_ _02553_ _02599_ _02600_ VGND VGND VPWR VPWR _02601_ sky130_fd_sc_hd__a21o_1
X_13488_ _04690_ _07112_ _03611_ _03612_ VGND VGND VPWR VPWR _03614_ sky130_fd_sc_hd__a22o_1
X_16276_ _03410_ _06528_ _06565_ _06539_ _06520_ VGND VGND VPWR VPWR _06650_ sky130_fd_sc_hd__o32a_1
XFILLER_0_125_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_124_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18015_ _08459_ _08460_ _08540_ VGND VGND VPWR VPWR _08543_ sky130_fd_sc_hd__and3_1
X_15227_ _05513_ _05381_ VGND VGND VPWR VPWR _05514_ sky130_fd_sc_hd__nand2_1
X_12439_ _02479_ _02481_ VGND VGND VPWR VPWR _02532_ sky130_fd_sc_hd__nor2_1
XFILLER_0_112_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15158_ _05316_ _05433_ _05436_ VGND VGND VPWR VPWR _05438_ sky130_fd_sc_hd__o21ai_2
X_14109_ _04291_ _04292_ VGND VGND VPWR VPWR _04293_ sky130_fd_sc_hd__nand2_1
X_15089_ _05360_ _05362_ VGND VGND VPWR VPWR _05363_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_38_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18917_ clknet_4_13_0_clk _00071_ VGND VGND VPWR VPWR ApproximateM_inst.lob_16.lob2.genblk1\[3\].genblk1.mux.sel
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_38_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09650_ _05693_ VGND VGND VPWR VPWR _05704_ sky130_fd_sc_hd__buf_6
X_18848_ clknet_4_6_0_clk net307 VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__dfxtp_1
X_09581_ _04842_ _04930_ _04919_ VGND VGND VPWR VPWR _04952_ sky130_fd_sc_hd__a21o_1
X_18779_ _09292_ VGND VGND VPWR VPWR _00084_ sky130_fd_sc_hd__buf_1
XFILLER_0_89_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_147_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_888 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_143_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_131_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold130 net85 VGND VGND VPWR VPWR net293 sky130_fd_sc_hd__dlygate4sd3_1
Xhold141 _00033_ VGND VGND VPWR VPWR net304 sky130_fd_sc_hd__dlygate4sd3_1
Xhold152 salida\[2\] VGND VGND VPWR VPWR net315 sky130_fd_sc_hd__buf_1
XFILLER_0_130_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09917_ _08539_ _08594_ VGND VGND VPWR VPWR _08605_ sky130_fd_sc_hd__xnor2_2
XTAP_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09848_ _07788_ VGND VGND VPWR VPWR _07853_ sky130_fd_sc_hd__clkbuf_8
X_09779_ cla_inst.in1\[25\] VGND VGND VPWR VPWR _07102_ sky130_fd_sc_hd__buf_4
XTAP_2302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11810_ _01747_ _01901_ _01902_ VGND VGND VPWR VPWR _01903_ sky130_fd_sc_hd__a21bo_2
XTAP_2324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12790_ _01446_ _01449_ _01448_ VGND VGND VPWR VPWR _02883_ sky130_fd_sc_hd__o21ai_1
XTAP_2335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11741_ _01591_ _01590_ VGND VGND VPWR VPWR _01834_ sky130_fd_sc_hd__and2b_1
XTAP_2368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14460_ _04628_ _04629_ _04674_ _04675_ VGND VGND VPWR VPWR _04677_ sky130_fd_sc_hd__a2bb2o_1
X_11672_ _01763_ _01762_ _01716_ _01713_ VGND VGND VPWR VPWR _01765_ sky130_fd_sc_hd__o211a_1
XTAP_1678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13411_ _03355_ _03362_ _03529_ VGND VGND VPWR VPWR _03530_ sky130_fd_sc_hd__a21oi_1
X_10623_ _00715_ VGND VGND VPWR VPWR _00716_ sky130_fd_sc_hd__buf_6
XFILLER_0_126_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14391_ _04447_ _04455_ VGND VGND VPWR VPWR _04601_ sky130_fd_sc_hd__and2_1
XFILLER_0_153_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13342_ _00509_ VGND VGND VPWR VPWR _03455_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_91_471 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16130_ _06489_ _06490_ _01677_ VGND VGND VPWR VPWR _06491_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10554_ _05464_ _07962_ _05715_ _05453_ VGND VGND VPWR VPWR _00647_ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13273_ _03574_ _05050_ net241 _03378_ VGND VGND VPWR VPWR _03379_ sky130_fd_sc_hd__a22o_1
X_16061_ _06200_ _06246_ VGND VGND VPWR VPWR _06416_ sky130_fd_sc_hd__or2_1
X_10485_ _00370_ _00373_ _00576_ _00577_ VGND VGND VPWR VPWR _00578_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_122_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15012_ _01873_ _03067_ VGND VGND VPWR VPWR _05280_ sky130_fd_sc_hd__nand2_1
X_12224_ _02302_ _02314_ _02315_ _02316_ VGND VGND VPWR VPWR _02317_ sky130_fd_sc_hd__o211a_1
XFILLER_0_20_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12155_ _07352_ _04056_ VGND VGND VPWR VPWR _02248_ sky130_fd_sc_hd__nand2_1
X_11106_ _01196_ _01197_ _01187_ _01192_ VGND VGND VPWR VPWR _01199_ sky130_fd_sc_hd__o211ai_2
X_12086_ _02178_ VGND VGND VPWR VPWR _02179_ sky130_fd_sc_hd__inv_2
X_16963_ _06655_ _07394_ _07396_ _07113_ VGND VGND VPWR VPWR _07397_ sky130_fd_sc_hd__a22o_1
X_18702_ _06776_ _09183_ net69 VGND VGND VPWR VPWR _09233_ sky130_fd_sc_hd__a21oi_1
X_11037_ _01127_ _01129_ VGND VGND VPWR VPWR _01130_ sky130_fd_sc_hd__nand2_1
X_15914_ _06257_ _06236_ VGND VGND VPWR VPWR _06259_ sky130_fd_sc_hd__or2b_1
X_16894_ _07310_ _07321_ VGND VGND VPWR VPWR _07322_ sky130_fd_sc_hd__or2_1
X_18633_ _09119_ _09180_ VGND VGND VPWR VPWR _09181_ sky130_fd_sc_hd__or2_1
X_15845_ _06074_ _06137_ VGND VGND VPWR VPWR _06185_ sky130_fd_sc_hd__nand2_1
XFILLER_0_87_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18564_ salida\[4\] _09114_ _09118_ salida\[36\] _09128_ VGND VGND VPWR VPWR _09133_
+ sky130_fd_sc_hd__a221o_1
X_15776_ _06108_ _06109_ VGND VGND VPWR VPWR _06110_ sky130_fd_sc_hd__nand2_1
X_12988_ _03080_ VGND VGND VPWR VPWR _03081_ sky130_fd_sc_hd__buf_4
X_17515_ _07997_ _07998_ VGND VGND VPWR VPWR _07999_ sky130_fd_sc_hd__nor2_1
X_14727_ _04867_ _04868_ _04879_ VGND VGND VPWR VPWR _04968_ sky130_fd_sc_hd__nand3_1
XFILLER_0_86_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11939_ _06008_ _05584_ _03421_ _04220_ VGND VGND VPWR VPWR _02032_ sky130_fd_sc_hd__and4_1
X_18495_ _03155_ _06451_ VGND VGND VPWR VPWR _09063_ sky130_fd_sc_hd__nor2_1
XFILLER_0_28_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17446_ _02974_ _03119_ _05306_ _07923_ VGND VGND VPWR VPWR _07924_ sky130_fd_sc_hd__o31a_1
X_14658_ _04891_ _04892_ VGND VGND VPWR VPWR _04893_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_46_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13609_ _03741_ _03746_ VGND VGND VPWR VPWR _03747_ sky130_fd_sc_hd__or2_1
X_17377_ _07843_ _07847_ VGND VGND VPWR VPWR _07848_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_15_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14589_ _04816_ _04817_ VGND VGND VPWR VPWR _04818_ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_600 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_131_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16328_ _03089_ _06495_ _06706_ _06626_ VGND VGND VPWR VPWR _06707_ sky130_fd_sc_hd__o211a_1
XFILLER_0_15_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_858 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_152_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16259_ _06470_ _06631_ VGND VGND VPWR VPWR _06632_ sky130_fd_sc_hd__and2_1
XFILLER_0_51_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09702_ _06234_ _06245_ _06256_ VGND VGND VPWR VPWR _06267_ sky130_fd_sc_hd__nand3_1
X_09633_ _05464_ _05388_ _05497_ _05508_ VGND VGND VPWR VPWR _05519_ sky130_fd_sc_hd__a22o_1
XFILLER_0_65_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09564_ _04318_ _04744_ _04755_ VGND VGND VPWR VPWR _04766_ sky130_fd_sc_hd__nand3_2
XFILLER_0_77_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_744 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09495_ _03815_ VGND VGND VPWR VPWR _04012_ sky130_fd_sc_hd__buf_8
XFILLER_0_77_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_147_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_104_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_104_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10270_ _00362_ _00134_ VGND VGND VPWR VPWR _00363_ sky130_fd_sc_hd__nand2_1
XFILLER_0_103_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13960_ _00645_ _09256_ VGND VGND VPWR VPWR _04130_ sky130_fd_sc_hd__nand2_1
X_12911_ _04493_ ApproximateM_inst.lob_16.lob2.genblk1\[12\].genblk1.mux.sel ApproximateM_inst.lob_16.lob2.genblk1\[11\].genblk1.mux.sel
+ VGND VGND VPWR VPWR _03004_ sky130_fd_sc_hd__or3_4
X_13891_ _04052_ _04053_ _04054_ VGND VGND VPWR VPWR _04055_ sky130_fd_sc_hd__or3_1
XFILLER_0_69_700 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15630_ _05947_ _05951_ _03202_ VGND VGND VPWR VPWR _05952_ sky130_fd_sc_hd__o21ai_1
XTAP_2110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12842_ _02895_ _02915_ VGND VGND VPWR VPWR _02935_ sky130_fd_sc_hd__nand2_1
XTAP_2121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15561_ _05789_ _05796_ _05876_ VGND VGND VPWR VPWR _05877_ sky130_fd_sc_hd__a21oi_1
XTAP_2165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12773_ _02853_ _02865_ VGND VGND VPWR VPWR _02866_ sky130_fd_sc_hd__xnor2_1
XTAP_2176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17300_ _07762_ _07763_ VGND VGND VPWR VPWR _07764_ sky130_fd_sc_hd__nor2_1
X_14512_ _04726_ _04732_ VGND VGND VPWR VPWR _04734_ sky130_fd_sc_hd__xnor2_2
XTAP_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11724_ _04690_ _00218_ VGND VGND VPWR VPWR _01817_ sky130_fd_sc_hd__nand2_1
X_18280_ _03206_ _08812_ _08818_ _08830_ VGND VGND VPWR VPWR _08831_ sky130_fd_sc_hd__o211a_1
XTAP_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15492_ _04823_ _05797_ _05798_ _05801_ VGND VGND VPWR VPWR _09365_ sky130_fd_sc_hd__a31o_1
XTAP_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17231_ _03913_ _06913_ _03920_ VGND VGND VPWR VPWR _07689_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_138_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14443_ _00107_ _06482_ VGND VGND VPWR VPWR _04659_ sky130_fd_sc_hd__nand2_1
X_11655_ _01698_ _01744_ _01747_ VGND VGND VPWR VPWR _01748_ sky130_fd_sc_hd__or3_1
XFILLER_0_71_419 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_138_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_154_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10606_ _00349_ _00531_ _00529_ _00530_ VGND VGND VPWR VPWR _00699_ sky130_fd_sc_hd__a211oi_2
X_17162_ _07488_ _07612_ VGND VGND VPWR VPWR _07614_ sky130_fd_sc_hd__xnor2_1
X_14374_ _04435_ _04441_ _04434_ VGND VGND VPWR VPWR _04583_ sky130_fd_sc_hd__a21bo_1
X_11586_ _01677_ _01678_ _01672_ VGND VGND VPWR VPWR _01679_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_153_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16113_ _02983_ _02563_ _03173_ _06470_ _06472_ VGND VGND VPWR VPWR _06473_ sky130_fd_sc_hd__o311a_1
X_13325_ _03278_ _03288_ VGND VGND VPWR VPWR _03436_ sky130_fd_sc_hd__nand2_1
X_10537_ _00628_ _00629_ VGND VGND VPWR VPWR _00630_ sky130_fd_sc_hd__and2b_1
X_17093_ _07409_ _07424_ VGND VGND VPWR VPWR _07539_ sky130_fd_sc_hd__and2_1
XFILLER_0_40_828 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_56 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16044_ _06396_ _06397_ _05162_ VGND VGND VPWR VPWR _06398_ sky130_fd_sc_hd__a21o_1
X_10468_ _00204_ _00248_ _00410_ VGND VGND VPWR VPWR _00561_ sky130_fd_sc_hd__and3_1
X_13256_ _02963_ _03359_ _03360_ VGND VGND VPWR VPWR _03361_ sky130_fd_sc_hd__a21o_1
XFILLER_0_10_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12207_ _02148_ VGND VGND VPWR VPWR _02300_ sky130_fd_sc_hd__inv_2
X_13187_ _00666_ _00674_ _00672_ VGND VGND VPWR VPWR _03287_ sky130_fd_sc_hd__a21oi_2
X_10399_ _00341_ _00346_ VGND VGND VPWR VPWR _00492_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12138_ _02203_ _02228_ _02229_ VGND VGND VPWR VPWR _02231_ sky130_fd_sc_hd__nor3_1
X_17995_ _06426_ _06445_ _08521_ VGND VGND VPWR VPWR _08522_ sky130_fd_sc_hd__or3_1
X_12069_ _02079_ _02078_ VGND VGND VPWR VPWR _02162_ sky130_fd_sc_hd__nor2_1
X_16946_ _03101_ _06464_ _07351_ _07378_ VGND VGND VPWR VPWR _09387_ sky130_fd_sc_hd__o2bb2a_1
X_16877_ _07115_ VGND VGND VPWR VPWR _07303_ sky130_fd_sc_hd__clkbuf_4
X_18616_ salida\[25\] _09159_ _09160_ salida\[57\] _09163_ VGND VGND VPWR VPWR _09169_
+ sky130_fd_sc_hd__a221o_1
X_15828_ _06095_ _06165_ VGND VGND VPWR VPWR _06166_ sky130_fd_sc_hd__xnor2_1
X_18547_ _09117_ VGND VGND VPWR VPWR _09118_ sky130_fd_sc_hd__buf_2
X_15759_ _06089_ _06090_ VGND VGND VPWR VPWR _06091_ sky130_fd_sc_hd__nor2_1
XFILLER_0_47_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_747 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18478_ _09036_ _09008_ _09043_ VGND VGND VPWR VPWR _09044_ sky130_fd_sc_hd__and3_1
XFILLER_0_47_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_706 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_118_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17429_ _07902_ _07903_ _07904_ VGND VGND VPWR VPWR _07905_ sky130_fd_sc_hd__a21o_1
XFILLER_0_117_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_144_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_110 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_132_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_132_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_141_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_384 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09616_ net234 VGND VGND VPWR VPWR _05333_ sky130_fd_sc_hd__buf_6
XFILLER_0_92_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09547_ _04569_ VGND VGND VPWR VPWR _04580_ sky130_fd_sc_hd__buf_6
X_09478_ ApproximateM_inst.lob_16.lob1.genblk1\[11\].genblk1.mux.sel VGND VGND VPWR
+ VPWR _03826_ sky130_fd_sc_hd__buf_6
XFILLER_0_93_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11440_ _01529_ _01530_ _01532_ VGND VGND VPWR VPWR _01533_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_135_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire148 net149 VGND VGND VPWR VPWR net148 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_123_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_638 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11371_ _00821_ _01463_ _01382_ _01392_ VGND VGND VPWR VPWR _01464_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_61_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13110_ _00696_ _00697_ _00743_ _00744_ VGND VGND VPWR VPWR _03204_ sky130_fd_sc_hd__nor4_2
X_10322_ _00400_ _00414_ VGND VGND VPWR VPWR _00415_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_104_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14090_ _01521_ _05964_ _04269_ _04270_ VGND VGND VPWR VPWR _04272_ sky130_fd_sc_hd__a22o_1
XFILLER_0_104_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13041_ _02976_ _03132_ VGND VGND VPWR VPWR _03133_ sky130_fd_sc_hd__nor2_1
X_10253_ _00342_ _00345_ VGND VGND VPWR VPWR _00346_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_30_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10184_ _03377_ _04471_ _03903_ _03356_ VGND VGND VPWR VPWR _00277_ sky130_fd_sc_hd__a22o_1
XFILLER_0_100_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16800_ net334 _06951_ _06961_ _07218_ VGND VGND VPWR VPWR _07219_ sky130_fd_sc_hd__or4_4
X_17780_ _08279_ _08286_ VGND VGND VPWR VPWR _08287_ sky130_fd_sc_hd__and2_1
X_14992_ _05143_ _05153_ _05151_ VGND VGND VPWR VPWR _05258_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_89_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16731_ _06665_ _07143_ VGND VGND VPWR VPWR _07144_ sky130_fd_sc_hd__or2_1
X_13943_ _04635_ _04427_ cla_inst.in1\[27\] _07004_ VGND VGND VPWR VPWR _04112_ sky130_fd_sc_hd__and4_1
XFILLER_0_72_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16662_ _06983_ _06985_ _06981_ VGND VGND VPWR VPWR _07070_ sky130_fd_sc_hd__a21o_1
X_13874_ _04030_ _04036_ VGND VGND VPWR VPWR _04037_ sky130_fd_sc_hd__xnor2_2
X_18401_ _08907_ _08946_ _08960_ VGND VGND VPWR VPWR _08961_ sky130_fd_sc_hd__a21oi_1
X_15613_ _05931_ _05933_ VGND VGND VPWR VPWR _05934_ sky130_fd_sc_hd__or2_1
X_12825_ _02916_ _02917_ VGND VGND VPWR VPWR _02918_ sky130_fd_sc_hd__or2_1
X_16593_ _06346_ _06926_ _02358_ VGND VGND VPWR VPWR _06995_ sky130_fd_sc_hd__a21o_1
X_18332_ _01417_ _03143_ VGND VGND VPWR VPWR _08888_ sky130_fd_sc_hd__nand2_1
XFILLER_0_139_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15544_ _05846_ _05847_ _05858_ VGND VGND VPWR VPWR _05859_ sky130_fd_sc_hd__a21oi_1
XTAP_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12756_ _02847_ _02848_ VGND VGND VPWR VPWR _02849_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11707_ _01790_ _01798_ _01799_ VGND VGND VPWR VPWR _01800_ sky130_fd_sc_hd__or3_4
X_18263_ _01359_ _06512_ _03056_ VGND VGND VPWR VPWR _08813_ sky130_fd_sc_hd__a21boi_1
X_15475_ _05665_ _05668_ _05783_ VGND VGND VPWR VPWR _05784_ sky130_fd_sc_hd__o21ai_1
X_12687_ _07091_ VGND VGND VPWR VPWR _02780_ sky130_fd_sc_hd__clkinv_4
XFILLER_0_127_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17214_ _07554_ _07555_ VGND VGND VPWR VPWR _07671_ sky130_fd_sc_hd__and2b_1
X_14426_ _04638_ _04639_ VGND VGND VPWR VPWR _04640_ sky130_fd_sc_hd__or2_1
X_11638_ _01725_ _01726_ _01730_ VGND VGND VPWR VPWR _01731_ sky130_fd_sc_hd__a21boi_1
X_18194_ _08736_ _08737_ VGND VGND VPWR VPWR _08738_ sky130_fd_sc_hd__or2b_1
XFILLER_0_126_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_108_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17145_ _04725_ _06889_ VGND VGND VPWR VPWR _07595_ sky130_fd_sc_hd__and2_1
X_14357_ _04540_ VGND VGND VPWR VPWR _04564_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11569_ _03399_ _01659_ _01661_ VGND VGND VPWR VPWR _01662_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_123_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_141_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13308_ _05301_ _07004_ _07102_ _05279_ VGND VGND VPWR VPWR _03417_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17076_ _06944_ _06957_ _07207_ _06969_ VGND VGND VPWR VPWR _07520_ sky130_fd_sc_hd__a2bb2o_1
X_14288_ _04315_ _04331_ _04487_ _04488_ VGND VGND VPWR VPWR _04489_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_40_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16027_ _02989_ _03693_ VGND VGND VPWR VPWR _06379_ sky130_fd_sc_hd__nand2_1
X_13239_ _03295_ _03296_ _03339_ _03340_ VGND VGND VPWR VPWR _03342_ sky130_fd_sc_hd__a22o_2
XFILLER_0_20_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17978_ _08403_ _08448_ _08501_ VGND VGND VPWR VPWR _08503_ sky130_fd_sc_hd__or3_1
XFILLER_0_34_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16929_ _07168_ _07170_ _07259_ _07359_ VGND VGND VPWR VPWR _07360_ sky130_fd_sc_hd__a31o_1
XFILLER_0_79_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_872 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_153_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_599 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_118_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_118_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_579 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold89 net110 VGND VGND VPWR VPWR net252 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10940_ net242 _00196_ _09179_ _03345_ VGND VGND VPWR VPWR _01033_ sky130_fd_sc_hd__a22o_1
XFILLER_0_98_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10871_ _00910_ _00912_ VGND VGND VPWR VPWR _00964_ sky130_fd_sc_hd__and2_1
XFILLER_0_78_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12610_ _02662_ _02695_ _02700_ VGND VGND VPWR VPWR _02703_ sky130_fd_sc_hd__o21bai_1
X_13590_ _03512_ _03514_ VGND VGND VPWR VPWR _03726_ sky130_fd_sc_hd__and2_1
XFILLER_0_38_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_270 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_109_635 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12541_ _02616_ _02629_ VGND VGND VPWR VPWR _02634_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_136_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_109_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_471 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15260_ _05526_ _05527_ _05548_ VGND VGND VPWR VPWR _05549_ sky130_fd_sc_hd__o21ai_1
X_12472_ _02558_ _02560_ _02562_ _02564_ VGND VGND VPWR VPWR _02565_ sky130_fd_sc_hd__nor4_1
XFILLER_0_46_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14211_ _03745_ _04402_ VGND VGND VPWR VPWR _04405_ sky130_fd_sc_hd__nand2_1
X_11423_ _00197_ _01509_ _01515_ VGND VGND VPWR VPWR _01516_ sky130_fd_sc_hd__a21bo_1
X_15191_ _05351_ _05357_ VGND VGND VPWR VPWR _05474_ sky130_fd_sc_hd__nor2_1
XFILLER_0_105_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_123_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_9 _00516_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14142_ _04315_ _04316_ _04328_ VGND VGND VPWR VPWR _04330_ sky130_fd_sc_hd__o21a_1
X_11354_ _01446_ VGND VGND VPWR VPWR _01447_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_135 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10305_ _04143_ VGND VGND VPWR VPWR _00398_ sky130_fd_sc_hd__buf_4
X_11285_ _01312_ _01332_ _01333_ _01334_ VGND VGND VPWR VPWR _01378_ sky130_fd_sc_hd__nand4_2
X_14073_ _03561_ _03575_ _03060_ VGND VGND VPWR VPWR _04254_ sky130_fd_sc_hd__mux2_1
X_18950_ clknet_4_5_0_clk _09411_ VGND VGND VPWR VPWR salida\[3\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_131_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17901_ _08413_ _08418_ VGND VGND VPWR VPWR _08419_ sky130_fd_sc_hd__nor2_1
X_10236_ _08800_ _08811_ _00328_ VGND VGND VPWR VPWR _00329_ sky130_fd_sc_hd__a21o_1
XTAP_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13024_ _02975_ VGND VGND VPWR VPWR _03117_ sky130_fd_sc_hd__buf_4
X_18881_ clknet_4_15_0_clk net318 VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__dfxtp_1
X_17832_ _06508_ _08332_ _08334_ _08343_ VGND VGND VPWR VPWR _08345_ sky130_fd_sc_hd__a31o_1
X_10167_ _00258_ _00259_ VGND VGND VPWR VPWR _00260_ sky130_fd_sc_hd__xor2_1
XFILLER_0_83_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17763_ _06957_ _07035_ _07487_ _07593_ VGND VGND VPWR VPWR _08269_ sky130_fd_sc_hd__or4_2
X_14975_ _05237_ _05238_ VGND VGND VPWR VPWR _05239_ sky130_fd_sc_hd__and2_1
X_10098_ _00175_ VGND VGND VPWR VPWR _00191_ sky130_fd_sc_hd__buf_2
XFILLER_0_83_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16714_ _07125_ VGND VGND VPWR VPWR _07126_ sky130_fd_sc_hd__buf_2
X_13926_ _03509_ _05606_ _05246_ _03531_ VGND VGND VPWR VPWR _04093_ sky130_fd_sc_hd__a22oi_2
X_17694_ _08192_ _08193_ VGND VGND VPWR VPWR _08194_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_107_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16645_ _06959_ _06962_ VGND VGND VPWR VPWR _07051_ sky130_fd_sc_hd__nand2_1
X_13857_ _04016_ _04017_ VGND VGND VPWR VPWR _04018_ sky130_fd_sc_hd__nand2_1
XFILLER_0_57_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12808_ _01458_ _01460_ _02900_ VGND VGND VPWR VPWR _02901_ sky130_fd_sc_hd__o21a_2
XFILLER_0_69_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16576_ _06967_ _06975_ VGND VGND VPWR VPWR _06976_ sky130_fd_sc_hd__xor2_1
X_13788_ _00308_ _03940_ _03941_ VGND VGND VPWR VPWR _03942_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_146_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18315_ _08795_ _08842_ _08867_ VGND VGND VPWR VPWR _08869_ sky130_fd_sc_hd__and3_1
XTAP_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15527_ _05838_ _05839_ VGND VGND VPWR VPWR _05840_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_84_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12739_ _02776_ _02778_ _02798_ _02800_ VGND VGND VPWR VPWR _02832_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_139_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_120_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18246_ _08712_ _08726_ _08793_ VGND VGND VPWR VPWR _08794_ sky130_fd_sc_hd__or3_1
X_15458_ _05449_ _01317_ _05764_ _05761_ VGND VGND VPWR VPWR _05765_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_127_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14409_ _04619_ _04620_ VGND VGND VPWR VPWR _04621_ sky130_fd_sc_hd__and2_1
X_18177_ _08717_ _08718_ VGND VGND VPWR VPWR _08719_ sky130_fd_sc_hd__nor2_1
X_15389_ _05688_ _05689_ VGND VGND VPWR VPWR _05690_ sky130_fd_sc_hd__nor2_1
XFILLER_0_40_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17128_ _06469_ _06498_ _02980_ VGND VGND VPWR VPWR _07577_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09950_ _06667_ _06798_ VGND VGND VPWR VPWR _08962_ sky130_fd_sc_hd__and2_1
XFILLER_0_110_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17059_ _07499_ _07500_ VGND VGND VPWR VPWR _07501_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_110_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09881_ _08191_ _07820_ VGND VGND VPWR VPWR _08213_ sky130_fd_sc_hd__and2b_1
XTAP_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_842 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_91 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11070_ _01157_ _01158_ _01162_ VGND VGND VPWR VPWR _01163_ sky130_fd_sc_hd__a21o_1
XFILLER_0_102_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput79 net79 VGND VGND VPWR VPWR leds[7] sky130_fd_sc_hd__buf_2
X_10021_ _00107_ _00108_ _00111_ _00113_ VGND VGND VPWR VPWR _00114_ sky130_fd_sc_hd__and4_1
X_14760_ _05002_ _06482_ _07635_ _05003_ VGND VGND VPWR VPWR _05004_ sky130_fd_sc_hd__and4b_1
XFILLER_0_98_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11972_ _02023_ _02063_ _02064_ VGND VGND VPWR VPWR _02065_ sky130_fd_sc_hd__or3_1
XFILLER_0_98_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13711_ _03700_ _03711_ VGND VGND VPWR VPWR _03858_ sky130_fd_sc_hd__nand2_1
X_10923_ _00989_ _00997_ _01014_ _01015_ VGND VGND VPWR VPWR _01016_ sky130_fd_sc_hd__o211ai_4
X_14691_ net202 _04883_ _04926_ _04927_ VGND VGND VPWR VPWR _04929_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_58_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_691 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16430_ _06522_ _06525_ _06816_ _01113_ VGND VGND VPWR VPWR _06817_ sky130_fd_sc_hd__a211o_1
X_13642_ _03774_ _03781_ VGND VGND VPWR VPWR _03783_ sky130_fd_sc_hd__xnor2_2
X_10854_ _00943_ _00946_ VGND VGND VPWR VPWR _00947_ sky130_fd_sc_hd__xnor2_2
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16361_ _03083_ _03166_ _03086_ _03169_ _06477_ _03161_ VGND VGND VPWR VPWR _06742_
+ sky130_fd_sc_hd__mux4_1
X_13573_ _03705_ _03707_ VGND VGND VPWR VPWR _03708_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_67_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10785_ _00172_ VGND VGND VPWR VPWR _00878_ sky130_fd_sc_hd__clkbuf_8
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18100_ _08553_ _08554_ _08552_ VGND VGND VPWR VPWR _08635_ sky130_fd_sc_hd__o21ai_2
X_15312_ _05604_ _05605_ VGND VGND VPWR VPWR _05607_ sky130_fd_sc_hd__or2_1
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12524_ _02561_ _02615_ VGND VGND VPWR VPWR _02617_ sky130_fd_sc_hd__nand2_1
XFILLER_0_81_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16292_ _06665_ _06666_ _06582_ VGND VGND VPWR VPWR _06668_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18031_ _08473_ _08475_ _08558_ VGND VGND VPWR VPWR _08560_ sky130_fd_sc_hd__or3_1
X_15243_ _05434_ _05438_ _05530_ VGND VGND VPWR VPWR _05531_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_152_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12455_ _05671_ _09212_ _02546_ _02547_ VGND VGND VPWR VPWR _02548_ sky130_fd_sc_hd__a31o_1
X_11406_ _01496_ _01497_ _01430_ _01498_ VGND VGND VPWR VPWR _01499_ sky130_fd_sc_hd__o211a_1
X_15174_ _05443_ _05455_ VGND VGND VPWR VPWR _05456_ sky130_fd_sc_hd__xnor2_1
X_12386_ _02475_ _02478_ VGND VGND VPWR VPWR _02479_ sky130_fd_sc_hd__and2_1
XFILLER_0_105_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14125_ _04309_ _04310_ VGND VGND VPWR VPWR _04311_ sky130_fd_sc_hd__nor2_1
XFILLER_0_120_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11337_ _01347_ _01423_ _01429_ VGND VGND VPWR VPWR _01430_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_132_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18933_ clknet_4_12_0_clk _00087_ VGND VGND VPWR VPWR cla_inst.in2\[19\] sky130_fd_sc_hd__dfxtp_2
X_14056_ _04233_ _04235_ VGND VGND VPWR VPWR _04236_ sky130_fd_sc_hd__xnor2_2
X_11268_ _01358_ _01360_ VGND VGND VPWR VPWR _01361_ sky130_fd_sc_hd__or2_1
XFILLER_0_94_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13007_ _03091_ _03097_ _03099_ VGND VGND VPWR VPWR _03100_ sky130_fd_sc_hd__mux2_1
X_10219_ _05464_ _06689_ _08757_ _05508_ VGND VGND VPWR VPWR _00312_ sky130_fd_sc_hd__a22o_1
X_11199_ _01007_ _01012_ VGND VGND VPWR VPWR _01292_ sky130_fd_sc_hd__and2_1
X_18864_ clknet_4_4_0_clk net270 VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__dfxtp_1
X_17815_ _08324_ _08325_ VGND VGND VPWR VPWR _08326_ sky130_fd_sc_hd__nand2_1
XFILLER_0_27_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18795_ _09298_ _09305_ VGND VGND VPWR VPWR _09306_ sky130_fd_sc_hd__and2_1
X_17746_ _08249_ _08227_ _02329_ VGND VGND VPWR VPWR _08250_ sky130_fd_sc_hd__a21oi_1
X_14958_ _05109_ _05110_ _05111_ _05108_ _05106_ VGND VGND VPWR VPWR _05220_ sky130_fd_sc_hd__o32ai_4
XFILLER_0_49_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13909_ _03130_ _03172_ _03060_ VGND VGND VPWR VPWR _04075_ sky130_fd_sc_hd__mux2_1
X_17677_ _07126_ _07195_ _07318_ _07608_ VGND VGND VPWR VPWR _08175_ sky130_fd_sc_hd__or4_1
X_14889_ _00125_ _00459_ _05322_ _00151_ VGND VGND VPWR VPWR _05145_ sky130_fd_sc_hd__a22o_1
XFILLER_0_89_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16628_ _04864_ _06812_ _06529_ VGND VGND VPWR VPWR _07032_ sky130_fd_sc_hd__or3_4
XFILLER_0_58_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_812 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16559_ _06954_ _06956_ _00172_ VGND VGND VPWR VPWR _06957_ sky130_fd_sc_hd__a21bo_4
XFILLER_0_17_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_84_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18229_ _00789_ _07743_ _07390_ _03311_ VGND VGND VPWR VPWR _08775_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_60_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09933_ _05366_ _08757_ _05246_ _05508_ VGND VGND VPWR VPWR _08778_ sky130_fd_sc_hd__a22o_1
XFILLER_0_110_162 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09864_ _07352_ _07112_ _07265_ _07276_ VGND VGND VPWR VPWR _08028_ sky130_fd_sc_hd__a22o_1
XTAP_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09795_ _07254_ cla_inst.in1\[24\] _05693_ _07232_ VGND VGND VPWR VPWR _07276_ sky130_fd_sc_hd__a22o_1
XFILLER_0_84_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10570_ _00497_ _00504_ VGND VGND VPWR VPWR _00663_ sky130_fd_sc_hd__nand2_1
XFILLER_0_64_856 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_119_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_720 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12240_ _05301_ _07548_ _07591_ _05279_ VGND VGND VPWR VPWR _02333_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12171_ _02256_ _02261_ _02262_ _02263_ VGND VGND VPWR VPWR _02264_ sky130_fd_sc_hd__or4_4
X_11122_ _01129_ _01213_ _01210_ VGND VGND VPWR VPWR _01215_ sky130_fd_sc_hd__nand3_2
XFILLER_0_102_674 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11053_ _01020_ _01021_ _01078_ VGND VGND VPWR VPWR _01146_ sky130_fd_sc_hd__o21ai_1
X_15930_ _06200_ _03072_ _06249_ VGND VGND VPWR VPWR _06275_ sky130_fd_sc_hd__a21o_1
X_10004_ _09341_ _09345_ _09343_ _09346_ VGND VGND VPWR VPWR _09347_ sky130_fd_sc_hd__a2bb2oi_2
X_15861_ _06200_ _03149_ _06198_ VGND VGND VPWR VPWR _06201_ sky130_fd_sc_hd__a21oi_1
X_17600_ _07630_ _07511_ VGND VGND VPWR VPWR _08091_ sky130_fd_sc_hd__or2_1
X_14812_ _05059_ _05060_ VGND VGND VPWR VPWR _05062_ sky130_fd_sc_hd__nor2_1
X_18580_ _09125_ VGND VGND VPWR VPWR _09144_ sky130_fd_sc_hd__buf_2
X_15792_ _06058_ _06087_ _06126_ VGND VGND VPWR VPWR _06128_ sky130_fd_sc_hd__a21o_1
XFILLER_0_98_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17531_ _08014_ _08015_ VGND VGND VPWR VPWR _08016_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_87_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14743_ _04982_ _04983_ _04985_ VGND VGND VPWR VPWR _04986_ sky130_fd_sc_hd__nand3_4
XFILLER_0_59_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwb_buttons_leds_160 VGND VGND VPWR VPWR wb_buttons_leds_160/HI led_enb[9] sky130_fd_sc_hd__conb_1
XFILLER_0_58_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11955_ _00845_ _01962_ _01963_ VGND VGND VPWR VPWR _02048_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_98_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10906_ _00948_ _00952_ VGND VGND VPWR VPWR _00999_ sky130_fd_sc_hd__nand2_1
X_17462_ _07829_ _07830_ _07939_ VGND VGND VPWR VPWR _07941_ sky130_fd_sc_hd__a21boi_2
X_14674_ _04909_ _04910_ cla_inst.in2\[25\] _05486_ VGND VGND VPWR VPWR _04911_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_86_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11886_ _01945_ _01976_ _01978_ VGND VGND VPWR VPWR _01979_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_67_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16413_ _03083_ _06464_ _06748_ _06799_ VGND VGND VPWR VPWR _09411_ sky130_fd_sc_hd__o2bb2a_1
X_13625_ _03782_ cla_inst.in1\[22\] _08746_ _03848_ VGND VGND VPWR VPWR _03764_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_363 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10837_ _03717_ _03432_ VGND VGND VPWR VPWR _00930_ sky130_fd_sc_hd__nand2_1
X_17393_ _07863_ _07865_ VGND VGND VPWR VPWR _07866_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16344_ _03049_ _03064_ _06626_ VGND VGND VPWR VPWR _06724_ sky130_fd_sc_hd__and3_1
X_13556_ _03687_ _03688_ VGND VGND VPWR VPWR _03689_ sky130_fd_sc_hd__nand2_1
X_10768_ _00120_ _07123_ VGND VGND VPWR VPWR _00861_ sky130_fd_sc_hd__and2_4
X_12507_ _05595_ ApproximateM_inst.lob_16.lob2.genblk1\[5\].genblk1.mux.sel _07548_
+ _07581_ VGND VGND VPWR VPWR _02600_ sky130_fd_sc_hd__and4_1
XFILLER_0_124_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16275_ _06516_ VGND VGND VPWR VPWR _06649_ sky130_fd_sc_hd__buf_4
X_13487_ _05017_ _07156_ _03611_ _03612_ VGND VGND VPWR VPWR _03613_ sky130_fd_sc_hd__nand4_2
X_10699_ _00785_ _00791_ VGND VGND VPWR VPWR _00792_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_125_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18014_ _07039_ _08150_ _08538_ VGND VGND VPWR VPWR _08542_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_152_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15226_ _05378_ _05379_ VGND VGND VPWR VPWR _05513_ sky130_fd_sc_hd__or2b_1
X_12438_ _02526_ _02530_ VGND VGND VPWR VPWR _02531_ sky130_fd_sc_hd__or2_1
XFILLER_0_140_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15157_ _05316_ _05433_ _05436_ VGND VGND VPWR VPWR _05437_ sky130_fd_sc_hd__or3_1
XFILLER_0_140_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12369_ _02400_ _02461_ VGND VGND VPWR VPWR _02462_ sky130_fd_sc_hd__nor2_1
X_14108_ _06460_ _09311_ _04288_ _04289_ VGND VGND VPWR VPWR _04292_ sky130_fd_sc_hd__a22o_1
X_15088_ _05247_ _05254_ _05361_ VGND VGND VPWR VPWR _05362_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_129_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14039_ _04214_ _04215_ _04171_ _04172_ VGND VGND VPWR VPWR _04217_ sky130_fd_sc_hd__o211a_1
X_18916_ clknet_4_9_0_clk _00070_ VGND VGND VPWR VPWR ApproximateM_inst.lob_16.lob2.genblk1\[2\].genblk1.mux.sel
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_0_129_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18847_ clknet_4_1_0_clk net278 VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__dfxtp_1
X_09580_ _04842_ _04919_ _04930_ VGND VGND VPWR VPWR _04941_ sky130_fd_sc_hd__nand3_1
X_18778_ _09273_ _09291_ VGND VGND VPWR VPWR _09292_ sky130_fd_sc_hd__and2_1
XFILLER_0_145_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17729_ _08023_ _08129_ _08130_ VGND VGND VPWR VPWR _08232_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_148_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold120 net97 VGND VGND VPWR VPWR net283 sky130_fd_sc_hd__dlygate4sd3_1
Xhold131 _00015_ VGND VGND VPWR VPWR net294 sky130_fd_sc_hd__dlygate4sd3_1
Xhold142 ApproximateM_inst.lob_16.lob1.genblk1\[2\].genblk1.mux.sel VGND VGND VPWR
+ VPWR net305 sky130_fd_sc_hd__buf_1
Xhold153 salida\[1\] VGND VGND VPWR VPWR net316 sky130_fd_sc_hd__buf_1
XFILLER_0_0_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09916_ _08550_ _08583_ VGND VGND VPWR VPWR _08594_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_95_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09847_ _07777_ _07820_ VGND VGND VPWR VPWR _07842_ sky130_fd_sc_hd__or2_1
XTAP_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09778_ _07080_ VGND VGND VPWR VPWR _07091_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_69_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11740_ _05224_ _03673_ VGND VGND VPWR VPWR _01833_ sky130_fd_sc_hd__nand2_1
XTAP_2369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11671_ _01713_ _01716_ _01762_ _01763_ VGND VGND VPWR VPWR _01764_ sky130_fd_sc_hd__a211oi_2
XTAP_1679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_828 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13410_ _03527_ _03528_ VGND VGND VPWR VPWR _03529_ sky130_fd_sc_hd__nand2_1
X_10622_ _03750_ VGND VGND VPWR VPWR _00715_ sky130_fd_sc_hd__buf_12
X_14390_ _04454_ _04448_ VGND VGND VPWR VPWR _04600_ sky130_fd_sc_hd__and2b_1
XFILLER_0_107_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13341_ _05736_ _09248_ _03244_ _03452_ VGND VGND VPWR VPWR _03453_ sky130_fd_sc_hd__a31o_1
X_10553_ _00644_ _00645_ _05758_ _05975_ VGND VGND VPWR VPWR _00646_ sky130_fd_sc_hd__and4_1
XFILLER_0_24_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16060_ _06200_ _06246_ _06248_ _06414_ VGND VGND VPWR VPWR _06415_ sky130_fd_sc_hd__a211o_1
X_13272_ _03531_ _03366_ net224 _04569_ VGND VGND VPWR VPWR _03378_ sky130_fd_sc_hd__nand4_2
XFILLER_0_122_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10484_ _00555_ _00556_ _00575_ VGND VGND VPWR VPWR _00577_ sky130_fd_sc_hd__and3_1
XFILLER_0_106_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15011_ _05276_ _05277_ VGND VGND VPWR VPWR _05278_ sky130_fd_sc_hd__nor2_1
X_12223_ _02154_ _02157_ _02156_ VGND VGND VPWR VPWR _02316_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_110_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12154_ _02244_ _02246_ VGND VGND VPWR VPWR _02247_ sky130_fd_sc_hd__or2_1
X_11105_ _01187_ _01192_ _01196_ _01197_ VGND VGND VPWR VPWR _01198_ sky130_fd_sc_hd__a211o_1
X_12085_ ApproximateM_inst.lob_16.lob2.genblk1\[10\].genblk1.mux.sel _05290_ _00129_
+ _01031_ VGND VGND VPWR VPWR _02178_ sky130_fd_sc_hd__and4_1
X_16962_ _03324_ _03003_ _06814_ _07289_ VGND VGND VPWR VPWR _07396_ sky130_fd_sc_hd__a211oi_4
X_18701_ _09231_ VGND VGND VPWR VPWR _00059_ sky130_fd_sc_hd__buf_1
X_11036_ _06982_ _05845_ _01127_ _01128_ VGND VGND VPWR VPWR _01129_ sky130_fd_sc_hd__nand4_2
X_15913_ _06236_ _06257_ VGND VGND VPWR VPWR _06258_ sky130_fd_sc_hd__or2b_1
X_16893_ _07317_ _07320_ VGND VGND VPWR VPWR _07321_ sky130_fd_sc_hd__xnor2_1
X_15844_ _06071_ _06134_ _06136_ VGND VGND VPWR VPWR _06184_ sky130_fd_sc_hd__a21o_1
X_18632_ net24 net27 _09111_ _09178_ VGND VGND VPWR VPWR _09180_ sky130_fd_sc_hd__or4_1
X_15775_ _06100_ _06107_ VGND VGND VPWR VPWR _06109_ sky130_fd_sc_hd__or2_1
X_18563_ net259 _09098_ _09132_ _09126_ VGND VGND VPWR VPWR _00007_ sky130_fd_sc_hd__o211a_1
X_12987_ _03079_ VGND VGND VPWR VPWR _03080_ sky130_fd_sc_hd__buf_4
X_17514_ _07851_ _07878_ _07996_ VGND VGND VPWR VPWR _07998_ sky130_fd_sc_hd__nor3_1
X_14726_ _04882_ VGND VGND VPWR VPWR _04967_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11938_ _06982_ _04012_ _02029_ _02030_ VGND VGND VPWR VPWR _02031_ sky130_fd_sc_hd__a31o_1
X_18494_ _02951_ _09060_ _09061_ _02968_ VGND VGND VPWR VPWR _09062_ sky130_fd_sc_hd__a211o_1
XFILLER_0_115_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17445_ _06680_ _07918_ _07922_ VGND VGND VPWR VPWR _07923_ sky130_fd_sc_hd__nor3_1
XFILLER_0_129_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14657_ _04760_ _04763_ _04761_ VGND VGND VPWR VPWR _04892_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_24_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11869_ _04700_ VGND VGND VPWR VPWR _01962_ sky130_fd_sc_hd__buf_6
XFILLER_0_67_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13608_ _02963_ _03742_ _03745_ VGND VGND VPWR VPWR _03746_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_28_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17376_ _07845_ _07846_ VGND VGND VPWR VPWR _07847_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_145_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14588_ net243 _04686_ _04815_ VGND VGND VPWR VPWR _04817_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_82_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16327_ _01677_ _02125_ _03179_ VGND VGND VPWR VPWR _06706_ sky130_fd_sc_hd__or3_1
X_13539_ _03652_ _03669_ VGND VGND VPWR VPWR _03670_ sky130_fd_sc_hd__xor2_2
XFILLER_0_70_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16258_ _03086_ _03169_ _00881_ _03094_ _06477_ _02983_ VGND VGND VPWR VPWR _06631_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_125_596 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15209_ _05491_ _05493_ VGND VGND VPWR VPWR _05494_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_101_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16189_ _06508_ _06514_ _06555_ _06462_ VGND VGND VPWR VPWR _06556_ sky130_fd_sc_hd__a211o_1
XFILLER_0_140_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09701_ _04788_ _04799_ _04777_ VGND VGND VPWR VPWR _06256_ sky130_fd_sc_hd__a21bo_1
X_09632_ _05399_ VGND VGND VPWR VPWR _05508_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_65_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09563_ _03968_ _03979_ _04307_ VGND VGND VPWR VPWR _04755_ sky130_fd_sc_hd__a21o_1
XFILLER_0_77_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09494_ _03990_ VGND VGND VPWR VPWR _04001_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_81_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_214 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_552 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_144_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12910_ _03771_ ApproximateM_inst.lob_16.lob2.genblk1\[14\].genblk1.mux.sel VGND
+ VGND VPWR VPWR _03003_ sky130_fd_sc_hd__or2_4
X_13890_ _03879_ _03882_ VGND VGND VPWR VPWR _04054_ sky130_fd_sc_hd__nor2_1
X_12841_ _00884_ _02921_ _02932_ VGND VGND VPWR VPWR _02934_ sky130_fd_sc_hd__nor3_1
XFILLER_0_69_712 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15560_ _05786_ _05788_ VGND VGND VPWR VPWR _05876_ sky130_fd_sc_hd__nor2_1
XFILLER_0_57_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12772_ _02863_ _02864_ VGND VGND VPWR VPWR _02865_ sky130_fd_sc_hd__and2_1
XTAP_2155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14511_ _04730_ _04731_ VGND VGND VPWR VPWR _04732_ sky130_fd_sc_hd__and2_1
XTAP_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11723_ _01813_ _01815_ VGND VGND VPWR VPWR _01816_ sky130_fd_sc_hd__nor2_1
XFILLER_0_96_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15491_ _03573_ _05307_ _05800_ _03124_ VGND VGND VPWR VPWR _05801_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_83_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_139_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17230_ _03081_ _07686_ _07687_ _02973_ VGND VGND VPWR VPWR _07688_ sky130_fd_sc_hd__a211o_1
X_14442_ _04655_ _04656_ VGND VGND VPWR VPWR _04658_ sky130_fd_sc_hd__nor2_1
XTAP_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11654_ _01745_ cla_inst.in2\[20\] _01746_ _01357_ VGND VGND VPWR VPWR _01747_ sky130_fd_sc_hd__and4_4
XFILLER_0_153_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10605_ _00555_ _00556_ _00575_ VGND VGND VPWR VPWR _00698_ sky130_fd_sc_hd__nand3_1
XFILLER_0_24_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17161_ _07607_ _07611_ VGND VGND VPWR VPWR _07612_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_24_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14373_ _04573_ _04574_ _04579_ VGND VGND VPWR VPWR _04582_ sky130_fd_sc_hd__a21o_1
X_11585_ _05888_ VGND VGND VPWR VPWR _01678_ sky130_fd_sc_hd__buf_4
XFILLER_0_51_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16112_ _03049_ _02370_ _03175_ VGND VGND VPWR VPWR _06472_ sky130_fd_sc_hd__or3_1
X_13324_ _03431_ _03433_ _03374_ _03264_ VGND VGND VPWR VPWR _03435_ sky130_fd_sc_hd__a211oi_4
X_10536_ _00626_ _00627_ _00623_ VGND VGND VPWR VPWR _00629_ sky130_fd_sc_hd__a21o_1
X_17092_ _07483_ _07430_ _07535_ VGND VGND VPWR VPWR _07538_ sky130_fd_sc_hd__nor3_1
XFILLER_0_12_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_596 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16043_ _02997_ _01112_ VGND VGND VPWR VPWR _06397_ sky130_fd_sc_hd__or2_1
XFILLER_0_122_544 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13255_ _00757_ _00906_ _00758_ VGND VGND VPWR VPWR _03360_ sky130_fd_sc_hd__o21ba_1
X_10467_ _00408_ _00409_ VGND VGND VPWR VPWR _00560_ sky130_fd_sc_hd__and2_1
X_12206_ _02295_ _02297_ _02298_ VGND VGND VPWR VPWR _02299_ sky130_fd_sc_hd__nor3_1
X_13186_ _03279_ _03285_ VGND VGND VPWR VPWR _03286_ sky130_fd_sc_hd__xnor2_2
X_10398_ net184 net340 _00489_ _00490_ VGND VGND VPWR VPWR _00491_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_102_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12137_ _02203_ _02228_ _02229_ VGND VGND VPWR VPWR _02230_ sky130_fd_sc_hd__or3_1
X_17994_ _03044_ _06444_ VGND VGND VPWR VPWR _08521_ sky130_fd_sc_hd__nor2_1
X_12068_ _02135_ _02159_ _02160_ VGND VGND VPWR VPWR _02161_ sky130_fd_sc_hd__o21ba_1
X_16945_ _07353_ _03202_ _07354_ _07377_ VGND VGND VPWR VPWR _07378_ sky130_fd_sc_hd__a31o_1
X_11019_ _05758_ VGND VGND VPWR VPWR _01112_ sky130_fd_sc_hd__buf_4
X_16876_ _06944_ VGND VGND VPWR VPWR _07302_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_126_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18615_ net287 _09157_ _09168_ _09162_ VGND VGND VPWR VPWR _00028_ sky130_fd_sc_hd__o211a_1
X_15827_ _06163_ _06164_ VGND VGND VPWR VPWR _06165_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_35_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_126_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15758_ _03010_ _03012_ _03149_ _03067_ VGND VGND VPWR VPWR _06090_ sky130_fd_sc_hd__and4_1
X_18546_ net27 _09115_ _09116_ VGND VGND VPWR VPWR _09117_ sky130_fd_sc_hd__nor3_2
XFILLER_0_47_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14709_ _04819_ _04816_ VGND VGND VPWR VPWR _04949_ sky130_fd_sc_hd__nand2_1
X_15689_ _05947_ _05951_ _05945_ VGND VGND VPWR VPWR _06016_ sky130_fd_sc_hd__o21a_1
X_18477_ _09041_ _09042_ VGND VGND VPWR VPWR _09043_ sky130_fd_sc_hd__xor2_1
XFILLER_0_51_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_759 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_117_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17428_ _07902_ _07903_ _06516_ VGND VGND VPWR VPWR _07904_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_90_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_145_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17359_ _02977_ _07657_ net168 _06753_ VGND VGND VPWR VPWR _07828_ sky130_fd_sc_hd__nand4_1
XFILLER_0_126_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_144_168 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_140_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_140_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09615_ _05311_ VGND VGND VPWR VPWR _05322_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_97_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09546_ cla_inst.in1\[16\] VGND VGND VPWR VPWR _04569_ sky130_fd_sc_hd__buf_6
XFILLER_0_66_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09477_ _03804_ VGND VGND VPWR VPWR _03815_ sky130_fd_sc_hd__buf_6
XFILLER_0_109_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_707 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_135_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire116 _08251_ VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_136_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire149 _09108_ VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_33_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11370_ _00797_ _00820_ _00819_ VGND VGND VPWR VPWR _01463_ sky130_fd_sc_hd__o21a_1
XFILLER_0_150_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10321_ _00412_ _00413_ VGND VGND VPWR VPWR _00414_ sky130_fd_sc_hd__and2b_1
XFILLER_0_131_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13040_ _02977_ _03131_ VGND VGND VPWR VPWR _03132_ sky130_fd_sc_hd__or2_1
X_10252_ _00343_ _00344_ VGND VGND VPWR VPWR _00345_ sky130_fd_sc_hd__and2b_1
X_10183_ _03465_ _04886_ VGND VGND VPWR VPWR _00276_ sky130_fd_sc_hd__and2_1
X_14991_ _05132_ _05255_ VGND VGND VPWR VPWR _05256_ sky130_fd_sc_hd__xnor2_1
X_13942_ _00294_ cla_inst.in1\[27\] _07004_ _04351_ VGND VGND VPWR VPWR _04111_ sky130_fd_sc_hd__a22oi_1
X_16730_ _07042_ VGND VGND VPWR VPWR _07143_ sky130_fd_sc_hd__clkbuf_4
X_16661_ _07066_ _07067_ VGND VGND VPWR VPWR _07068_ sky130_fd_sc_hd__or2b_1
X_13873_ _04033_ _04035_ VGND VGND VPWR VPWR _04036_ sky130_fd_sc_hd__xnor2_2
X_15612_ _05929_ _05930_ _05892_ VGND VGND VPWR VPWR _05933_ sky130_fd_sc_hd__a21oi_1
X_18400_ _08958_ _08959_ VGND VGND VPWR VPWR _08960_ sky130_fd_sc_hd__nand2_1
X_12824_ _01496_ _01500_ VGND VGND VPWR VPWR _02917_ sky130_fd_sc_hd__nor2_2
XFILLER_0_97_851 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16592_ _06990_ _06991_ _06836_ VGND VGND VPWR VPWR _06994_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_69_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_84_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15543_ _05855_ _05857_ VGND VGND VPWR VPWR _05858_ sky130_fd_sc_hd__and2_1
X_18331_ _06426_ _06448_ _08881_ _08882_ _08885_ VGND VGND VPWR VPWR _08886_ sky130_fd_sc_hd__o311a_1
XFILLER_0_97_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12755_ _02466_ _02398_ VGND VGND VPWR VPWR _02848_ sky130_fd_sc_hd__xnor2_1
XTAP_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_603 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_139_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11706_ _01236_ _01789_ _01760_ _01769_ VGND VGND VPWR VPWR _01799_ sky130_fd_sc_hd__a211oi_2
X_18262_ _08773_ _08810_ VGND VGND VPWR VPWR _08812_ sky130_fd_sc_hd__xnor2_2
X_15474_ _05781_ _05782_ VGND VGND VPWR VPWR _05783_ sky130_fd_sc_hd__xor2_1
XTAP_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12686_ _07613_ VGND VGND VPWR VPWR _02779_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14425_ _04496_ _04631_ _04637_ VGND VGND VPWR VPWR _04639_ sky130_fd_sc_hd__o21a_1
X_17213_ _07586_ _07587_ _07667_ VGND VGND VPWR VPWR _07670_ sky130_fd_sc_hd__o21a_1
X_11637_ _01727_ _01728_ _01729_ VGND VGND VPWR VPWR _01730_ sky130_fd_sc_hd__or3_1
X_18193_ _08660_ _08697_ _08734_ VGND VGND VPWR VPWR _08737_ sky130_fd_sc_hd__or3b_1
XFILLER_0_25_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17144_ _06572_ _07487_ _07593_ _06563_ VGND VGND VPWR VPWR _07594_ sky130_fd_sc_hd__o22a_1
X_14356_ _04560_ _04562_ _03539_ VGND VGND VPWR VPWR _04563_ sky130_fd_sc_hd__mux2_1
X_11568_ ApproximateM_inst.lob_16.lob2.genblk1\[6\].genblk1.mux.sel _03826_ _03388_
+ _06008_ VGND VGND VPWR VPWR _01661_ sky130_fd_sc_hd__a22o_1
XFILLER_0_52_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13307_ _03414_ _03415_ VGND VGND VPWR VPWR _03416_ sky130_fd_sc_hd__xor2_2
XFILLER_0_123_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10519_ _03881_ _03892_ _05028_ VGND VGND VPWR VPWR _00612_ sky130_fd_sc_hd__and3_1
X_17075_ _06880_ _06944_ _06957_ _07115_ VGND VGND VPWR VPWR _07519_ sky130_fd_sc_hd__or4_1
X_14287_ _04470_ _04472_ _04486_ VGND VGND VPWR VPWR _04488_ sky130_fd_sc_hd__nand3_2
XFILLER_0_0_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11499_ _08713_ _00165_ _01590_ _01591_ VGND VGND VPWR VPWR _01592_ sky130_fd_sc_hd__a31o_1
XFILLER_0_122_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16026_ _02989_ _03693_ VGND VGND VPWR VPWR _06378_ sky130_fd_sc_hd__or2_1
X_13238_ _03295_ _03296_ _03339_ _03340_ VGND VGND VPWR VPWR _03341_ sky130_fd_sc_hd__nand4_4
XFILLER_0_21_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13169_ _00655_ _00657_ VGND VGND VPWR VPWR _03268_ sky130_fd_sc_hd__nand2_2
X_17977_ _08403_ _08448_ _08501_ VGND VGND VPWR VPWR _08502_ sky130_fd_sc_hd__o21ai_2
X_16928_ _07165_ _07358_ _07258_ VGND VGND VPWR VPWR _07359_ sky130_fd_sc_hd__a21oi_1
X_16859_ _07240_ _07244_ VGND VGND VPWR VPWR _07283_ sky130_fd_sc_hd__nand2_1
XFILLER_0_153_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_149_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_52 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_884 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18529_ _09097_ VGND VGND VPWR VPWR _09098_ sky130_fd_sc_hd__buf_2
XFILLER_0_153_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_117_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_132_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10870_ _00775_ _00962_ VGND VGND VPWR VPWR _00963_ sky130_fd_sc_hd__nor2_2
XFILLER_0_79_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09529_ ApproximateM_inst.lob_16.lob1.genblk2.mux_final.sel VGND VGND VPWR VPWR _04384_
+ sky130_fd_sc_hd__buf_4
XFILLER_0_149_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12540_ _02590_ _02632_ VGND VGND VPWR VPWR _02633_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_93_364 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_148_282 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_109_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_483 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12471_ _00846_ _00214_ _02563_ VGND VGND VPWR VPWR _02564_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_124_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14210_ _04403_ VGND VGND VPWR VPWR _04404_ sky130_fd_sc_hd__inv_2
X_11422_ _01151_ _00196_ _00871_ _03848_ VGND VGND VPWR VPWR _01515_ sky130_fd_sc_hd__a22o_1
XFILLER_0_124_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15190_ _05339_ _05472_ VGND VGND VPWR VPWR _05473_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_50_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14141_ _04317_ _04327_ VGND VGND VPWR VPWR _04328_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_22_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11353_ _01370_ _01374_ _01444_ _01445_ VGND VGND VPWR VPWR _01446_ sky130_fd_sc_hd__o211a_1
XFILLER_0_105_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10304_ _00395_ _00380_ _00381_ VGND VGND VPWR VPWR _00397_ sky130_fd_sc_hd__nand3_1
X_14072_ _04240_ _04244_ _04252_ VGND VGND VPWR VPWR _09382_ sky130_fd_sc_hd__nand3_1
XFILLER_0_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11284_ _01337_ _01366_ _01367_ VGND VGND VPWR VPWR _01377_ sky130_fd_sc_hd__nor3_2
XFILLER_0_120_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13023_ _03100_ _03115_ _03080_ VGND VGND VPWR VPWR _03116_ sky130_fd_sc_hd__mux2_2
X_17900_ _08018_ _08415_ _08417_ VGND VGND VPWR VPWR _08418_ sky130_fd_sc_hd__o21a_1
X_10235_ _08822_ _08908_ VGND VGND VPWR VPWR _00328_ sky130_fd_sc_hd__and2_1
X_18880_ clknet_4_15_0_clk net317 VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__dfxtp_1
X_17831_ _06421_ _08335_ _08336_ _08342_ VGND VGND VPWR VPWR _08343_ sky130_fd_sc_hd__a31o_1
X_10166_ _00216_ _00220_ VGND VGND VPWR VPWR _00259_ sky130_fd_sc_hd__or2_1
X_17762_ _07130_ _07487_ _07593_ _07143_ VGND VGND VPWR VPWR _08268_ sky130_fd_sc_hd__o22ai_1
X_14974_ _05229_ _05236_ VGND VGND VPWR VPWR _05238_ sky130_fd_sc_hd__nand2_1
X_10097_ _00189_ VGND VGND VPWR VPWR _00190_ sky130_fd_sc_hd__clkbuf_4
X_16713_ _06871_ _07032_ _00213_ VGND VGND VPWR VPWR _07125_ sky130_fd_sc_hd__a21bo_2
X_13925_ _03934_ _03936_ _03937_ VGND VGND VPWR VPWR _04092_ sky130_fd_sc_hd__and3_1
X_17693_ _07630_ _07621_ VGND VGND VPWR VPWR _08193_ sky130_fd_sc_hd__nor2_1
X_13856_ _00204_ _01866_ _04015_ VGND VGND VPWR VPWR _04017_ sky130_fd_sc_hd__a21o_1
X_16644_ _06876_ _06885_ _06964_ VGND VGND VPWR VPWR _07050_ sky130_fd_sc_hd__and3_1
XFILLER_0_76_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12807_ _00887_ _00867_ VGND VGND VPWR VPWR _02900_ sky130_fd_sc_hd__xor2_2
XFILLER_0_147_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13787_ _03782_ _05693_ _05606_ _03848_ VGND VGND VPWR VPWR _03941_ sky130_fd_sc_hd__a22o_1
XFILLER_0_57_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16575_ _06973_ _06974_ VGND VGND VPWR VPWR _06975_ sky130_fd_sc_hd__or2_1
X_10999_ _01086_ _01091_ VGND VGND VPWR VPWR _01092_ sky130_fd_sc_hd__xnor2_2
X_18314_ _08795_ _08842_ _08867_ VGND VGND VPWR VPWR _08868_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_32_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15526_ _02998_ _03153_ _05743_ _05742_ VGND VGND VPWR VPWR _05839_ sky130_fd_sc_hd__a31o_1
X_12738_ _02830_ _02800_ VGND VGND VPWR VPWR _02831_ sky130_fd_sc_hd__and2b_1
XFILLER_0_123_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15457_ _05762_ VGND VGND VPWR VPWR _05764_ sky130_fd_sc_hd__inv_2
XFILLER_0_127_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18245_ _08791_ _08792_ VGND VGND VPWR VPWR _08793_ sky130_fd_sc_hd__and2_1
X_12669_ _02753_ _02761_ VGND VGND VPWR VPWR _02762_ sky130_fd_sc_hd__nor2_2
XFILLER_0_115_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14408_ _04616_ _04618_ _04612_ VGND VGND VPWR VPWR _04620_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_113_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15388_ _05530_ _05676_ _05687_ VGND VGND VPWR VPWR _05689_ sky130_fd_sc_hd__nor3_1
X_18176_ _07608_ _07741_ _07859_ _07394_ VGND VGND VPWR VPWR _08718_ sky130_fd_sc_hd__o211a_1
XFILLER_0_4_336 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_114_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14339_ _04542_ _04543_ _04423_ _04424_ VGND VGND VPWR VPWR _04545_ sky130_fd_sc_hd__o211a_2
X_17127_ _06331_ _06790_ _07575_ _00558_ VGND VGND VPWR VPWR _07576_ sky130_fd_sc_hd__a22o_1
XFILLER_0_12_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_171 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17058_ _07018_ _07106_ VGND VGND VPWR VPWR _07500_ sky130_fd_sc_hd__nor2_1
X_16009_ _06356_ _06357_ _06358_ VGND VGND VPWR VPWR _06359_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_148_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09880_ _07820_ _08191_ VGND VGND VPWR VPWR _08202_ sky130_fd_sc_hd__and2b_1
XFILLER_0_111_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10020_ _09350_ _07570_ _07602_ _00112_ VGND VGND VPWR VPWR _00113_ sky130_fd_sc_hd__a22o_1
X_11971_ _02061_ _02062_ VGND VGND VPWR VPWR _02064_ sky130_fd_sc_hd__xnor2_1
X_13710_ _03447_ _03710_ VGND VGND VPWR VPWR _03857_ sky130_fd_sc_hd__or2_1
X_10922_ _00998_ _00999_ _01013_ VGND VGND VPWR VPWR _01015_ sky130_fd_sc_hd__nand3_2
X_14690_ _04882_ _04883_ _04926_ _04927_ VGND VGND VPWR VPWR _04928_ sky130_fd_sc_hd__and4_1
XFILLER_0_58_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13641_ _03775_ _03780_ VGND VGND VPWR VPWR _03781_ sky130_fd_sc_hd__xor2_2
X_10853_ _00944_ _00945_ VGND VGND VPWR VPWR _00946_ sky130_fd_sc_hd__and2b_1
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16360_ _06470_ _06740_ VGND VGND VPWR VPWR _06741_ sky130_fd_sc_hd__and2_1
XFILLER_0_149_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13572_ _09352_ _00398_ VGND VGND VPWR VPWR _03707_ sky130_fd_sc_hd__nand2_1
X_10784_ _00203_ VGND VGND VPWR VPWR _00877_ sky130_fd_sc_hd__buf_4
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15311_ _05503_ _05506_ _05603_ VGND VGND VPWR VPWR _05605_ sky130_fd_sc_hd__and3_1
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_835 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_137_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12523_ _02561_ _02615_ VGND VGND VPWR VPWR _02616_ sky130_fd_sc_hd__or2_1
XFILLER_0_109_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16291_ _06563_ _06665_ VGND VGND VPWR VPWR _06666_ sky130_fd_sc_hd__nor2_1
XFILLER_0_125_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15242_ _05318_ _05438_ _05434_ VGND VGND VPWR VPWR _05530_ sky130_fd_sc_hd__a21oi_2
X_18030_ _08473_ _08475_ _08558_ VGND VGND VPWR VPWR _08559_ sky130_fd_sc_hd__o21ai_2
X_12454_ _05562_ _05584_ ApproximateM_inst.lob_16.lob1.genblk1\[1\].genblk1.mux.sel
+ ApproximateM_inst.lob_16.lob1.mux.sel VGND VGND VPWR VPWR _02547_ sky130_fd_sc_hd__and4_1
XFILLER_0_124_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11405_ _01422_ _01432_ VGND VGND VPWR VPWR _01498_ sky130_fd_sc_hd__or2b_2
XFILLER_0_90_890 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15173_ _05452_ _05454_ VGND VGND VPWR VPWR _05455_ sky130_fd_sc_hd__and2_1
XFILLER_0_78_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12385_ _02402_ _02477_ VGND VGND VPWR VPWR _02478_ sky130_fd_sc_hd__nor2_1
XFILLER_0_151_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14124_ _04302_ _04117_ _04308_ VGND VGND VPWR VPWR _04310_ sky130_fd_sc_hd__nor3_1
XFILLER_0_50_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11336_ _01424_ _01428_ VGND VGND VPWR VPWR _01429_ sky130_fd_sc_hd__xnor2_2
X_14055_ _04058_ _04059_ _04234_ VGND VGND VPWR VPWR _04235_ sky130_fd_sc_hd__o21ai_4
X_18932_ clknet_4_12_0_clk _00086_ VGND VGND VPWR VPWR cla_inst.in2\[18\] sky130_fd_sc_hd__dfxtp_1
X_11267_ _01359_ _01357_ _01110_ VGND VGND VPWR VPWR _01360_ sky130_fd_sc_hd__a21oi_1
X_13006_ _03098_ VGND VGND VPWR VPWR _03099_ sky130_fd_sc_hd__buf_4
X_10218_ _05508_ _05366_ _06689_ _08757_ VGND VGND VPWR VPWR _00311_ sky130_fd_sc_hd__and4_1
X_18863_ clknet_4_4_0_clk net264 VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__dfxtp_1
X_11198_ _01004_ _01006_ VGND VGND VPWR VPWR _01291_ sky130_fd_sc_hd__and2_1
X_17814_ _08253_ _08254_ _08323_ VGND VGND VPWR VPWR _08325_ sky130_fd_sc_hd__a21o_1
XFILLER_0_118_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10149_ _00235_ _00241_ VGND VGND VPWR VPWR _00242_ sky130_fd_sc_hd__xnor2_1
X_18794_ _03000_ net48 _09301_ VGND VGND VPWR VPWR _09305_ sky130_fd_sc_hd__mux2_1
X_17745_ _02321_ _02325_ VGND VGND VPWR VPWR _08249_ sky130_fd_sc_hd__nand2_1
X_14957_ _05210_ _05218_ VGND VGND VPWR VPWR _05219_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_89_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13908_ _03930_ _04072_ _04073_ VGND VGND VPWR VPWR _04074_ sky130_fd_sc_hd__and3_1
X_17676_ _07394_ net146 _07604_ _07751_ VGND VGND VPWR VPWR _08174_ sky130_fd_sc_hd__a22o_1
X_14888_ _00362_ _06482_ _05003_ _05002_ VGND VGND VPWR VPWR _05144_ sky130_fd_sc_hd__a31o_1
XFILLER_0_134_45 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16627_ _06945_ _07030_ VGND VGND VPWR VPWR _07031_ sky130_fd_sc_hd__xnor2_1
X_13839_ _03805_ _03807_ _03996_ VGND VGND VPWR VPWR _03998_ sky130_fd_sc_hd__and3_1
XFILLER_0_43_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16558_ sel_op\[0\] _06804_ _06955_ VGND VGND VPWR VPWR _06956_ sky130_fd_sc_hd__or3_1
XFILLER_0_85_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15509_ _05817_ _05818_ _05813_ VGND VGND VPWR VPWR _05820_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_127_241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16489_ _06522_ _06525_ _06880_ _00515_ VGND VGND VPWR VPWR _06881_ sky130_fd_sc_hd__a211o_1
XFILLER_0_94_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18228_ _02045_ _00789_ _07743_ _07387_ VGND VGND VPWR VPWR _08774_ sky130_fd_sc_hd__or4_1
XFILLER_0_150_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18159_ _06366_ _07650_ _07596_ VGND VGND VPWR VPWR _08699_ sky130_fd_sc_hd__and3_1
XFILLER_0_7_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09932_ _05410_ _05366_ _08757_ _05246_ VGND VGND VPWR VPWR _08768_ sky130_fd_sc_hd__and4_1
XFILLER_0_110_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09863_ _07951_ _08006_ VGND VGND VPWR VPWR _08017_ sky130_fd_sc_hd__nand2_1
XTAP_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09794_ _07232_ _07254_ _06722_ _05704_ VGND VGND VPWR VPWR _07265_ sky130_fd_sc_hd__nand4_2
XFILLER_0_84_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_450 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_119_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12170_ _02258_ _02260_ VGND VGND VPWR VPWR _02263_ sky130_fd_sc_hd__nor2_1
XFILLER_0_102_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11121_ _01129_ _01210_ _01213_ VGND VGND VPWR VPWR _01214_ sky130_fd_sc_hd__a21o_1
XFILLER_0_31_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_686 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11052_ _01120_ _01144_ VGND VGND VPWR VPWR _01145_ sky130_fd_sc_hd__xor2_1
X_10003_ net167 _06906_ _09005_ _09016_ VGND VGND VPWR VPWR _09346_ sky130_fd_sc_hd__o211ai_4
X_15860_ _03007_ VGND VGND VPWR VPWR _06200_ sky130_fd_sc_hd__clkbuf_4
X_14811_ _05056_ _05057_ _05058_ VGND VGND VPWR VPWR _05060_ sky130_fd_sc_hd__a21oi_1
X_15791_ _06124_ _06125_ VGND VGND VPWR VPWR _06126_ sky130_fd_sc_hd__nand2_1
X_17530_ _07931_ _07932_ _08013_ VGND VGND VPWR VPWR _08015_ sky130_fd_sc_hd__or3b_4
X_14742_ _04843_ _04848_ _04841_ VGND VGND VPWR VPWR _04985_ sky130_fd_sc_hd__a21bo_1
Xwb_buttons_leds_161 VGND VGND VPWR VPWR wb_buttons_leds_161/HI led_enb[10] sky130_fd_sc_hd__conb_1
X_11954_ _01964_ _02046_ VGND VGND VPWR VPWR _02047_ sky130_fd_sc_hd__and2_1
XFILLER_0_59_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10905_ _00942_ _00947_ VGND VGND VPWR VPWR _00998_ sky130_fd_sc_hd__nand2_1
X_14673_ _00109_ _09349_ _05388_ _05497_ VGND VGND VPWR VPWR _04910_ sky130_fd_sc_hd__and4_1
X_17461_ _07828_ _07827_ VGND VGND VPWR VPWR _07939_ sky130_fd_sc_hd__or2_1
X_11885_ _01890_ _01977_ VGND VGND VPWR VPWR _01978_ sky130_fd_sc_hd__nand2_1
X_13624_ _04078_ _01151_ _08746_ VGND VGND VPWR VPWR _03763_ sky130_fd_sc_hd__and3_1
X_16412_ _06649_ _06778_ _06779_ _06797_ VGND VGND VPWR VPWR _06799_ sky130_fd_sc_hd__a31o_1
X_10836_ _00927_ _00928_ VGND VGND VPWR VPWR _00929_ sky130_fd_sc_hd__and2b_1
XFILLER_0_67_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17392_ _06581_ _07741_ VGND VGND VPWR VPWR _07865_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13555_ _03685_ _03686_ VGND VGND VPWR VPWR _03688_ sky130_fd_sc_hd__nand2_1
X_16343_ _06671_ _06694_ _06719_ _06723_ _06427_ VGND VGND VPWR VPWR _09408_ sky130_fd_sc_hd__o32a_1
X_10767_ _00140_ _00139_ VGND VGND VPWR VPWR _00860_ sky130_fd_sc_hd__and2b_1
XFILLER_0_81_131 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12506_ _00832_ _00177_ _02551_ _02552_ VGND VGND VPWR VPWR _02599_ sky130_fd_sc_hd__a22o_1
X_16274_ _01746_ _06464_ _06648_ VGND VGND VPWR VPWR _09397_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_152_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13486_ _04351_ _04373_ cla_inst.in1\[24\] _05693_ VGND VGND VPWR VPWR _03612_ sky130_fd_sc_hd__nand4_2
X_10698_ _00786_ _00787_ _00789_ _00790_ VGND VGND VPWR VPWR _00791_ sky130_fd_sc_hd__o22ai_4
XFILLER_0_124_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15225_ _05510_ _05511_ VGND VGND VPWR VPWR _05512_ sky130_fd_sc_hd__or2_1
X_18013_ _08459_ _08460_ _08540_ VGND VGND VPWR VPWR _08541_ sky130_fd_sc_hd__a21oi_1
X_12437_ _02523_ _02525_ _02524_ VGND VGND VPWR VPWR _02530_ sky130_fd_sc_hd__o21a_1
XFILLER_0_152_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15156_ _05318_ _05434_ _05435_ VGND VGND VPWR VPWR _05436_ sky130_fd_sc_hd__o21a_1
XFILLER_0_10_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12368_ _02458_ _02460_ VGND VGND VPWR VPWR _02461_ sky130_fd_sc_hd__and2b_1
X_14107_ _04290_ VGND VGND VPWR VPWR _04291_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11319_ _01409_ _01411_ VGND VGND VPWR VPWR _01412_ sky130_fd_sc_hd__xor2_1
X_15087_ _05253_ _05248_ VGND VGND VPWR VPWR _05361_ sky130_fd_sc_hd__and2b_1
X_12299_ _02385_ net123 _02390_ _02391_ VGND VGND VPWR VPWR _02392_ sky130_fd_sc_hd__o211a_1
X_14038_ _04171_ _04172_ _04214_ _04215_ VGND VGND VPWR VPWR _04216_ sky130_fd_sc_hd__a211oi_2
X_18915_ clknet_4_8_0_clk _00069_ VGND VGND VPWR VPWR ApproximateM_inst.lob_16.lob2.genblk1\[1\].genblk1.mux.sel
+ sky130_fd_sc_hd__dfxtp_2
X_18846_ clknet_4_1_0_clk net272 VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__dfxtp_1
X_18777_ _02989_ net42 _09276_ VGND VGND VPWR VPWR _09291_ sky130_fd_sc_hd__mux2_1
X_15989_ _02977_ _01248_ VGND VGND VPWR VPWR _06337_ sky130_fd_sc_hd__nand2_1
XFILLER_0_54_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_145_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17728_ _01678_ _07355_ _02987_ VGND VGND VPWR VPWR _08231_ sky130_fd_sc_hd__or3b_1
X_17659_ _08153_ _08154_ VGND VGND VPWR VPWR _08155_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_148_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_194 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_890 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_116_789 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_130_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold110 net112 VGND VGND VPWR VPWR net273 sky130_fd_sc_hd__dlygate4sd3_1
Xhold121 _00026_ VGND VGND VPWR VPWR net284 sky130_fd_sc_hd__dlygate4sd3_1
Xhold132 net83 VGND VGND VPWR VPWR net295 sky130_fd_sc_hd__dlygate4sd3_1
Xhold143 net84 VGND VGND VPWR VPWR net306 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold154 op_code\[2\] VGND VGND VPWR VPWR net317 sky130_fd_sc_hd__clkbuf_2
X_09915_ _08561_ _08572_ VGND VGND VPWR VPWR _08583_ sky130_fd_sc_hd__and2b_1
XFILLER_0_95_60 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09846_ _07777_ _07820_ VGND VGND VPWR VPWR _07831_ sky130_fd_sc_hd__and2_1
XTAP_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09777_ _07069_ VGND VGND VPWR VPWR _07080_ sky130_fd_sc_hd__clkbuf_4
XTAP_2304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11670_ _01217_ _01219_ _01227_ VGND VGND VPWR VPWR _01763_ sky130_fd_sc_hd__nor3_1
XTAP_1669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10621_ _00712_ _00713_ VGND VGND VPWR VPWR _00714_ sky130_fd_sc_hd__nor2_1
XFILLER_0_107_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13340_ _06029_ _06051_ _00498_ _08169_ VGND VGND VPWR VPWR _03452_ sky130_fd_sc_hd__and4_1
X_10552_ _05366_ VGND VGND VPWR VPWR _00645_ sky130_fd_sc_hd__buf_6
XFILLER_0_134_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13271_ net172 net234 cla_inst.in1\[16\] _03345_ VGND VGND VPWR VPWR _03376_ sky130_fd_sc_hd__a22o_4
X_10483_ _00555_ _00556_ _00575_ VGND VGND VPWR VPWR _00576_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_51_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_121_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15010_ _05263_ _05171_ _05275_ VGND VGND VPWR VPWR _05277_ sky130_fd_sc_hd__and3_1
XFILLER_0_122_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12222_ _02154_ _02156_ _02157_ VGND VGND VPWR VPWR _02315_ sky130_fd_sc_hd__or3_1
XFILLER_0_121_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_735 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12153_ _02244_ _02245_ ApproximateM_inst.lob_16.lob2.genblk1\[5\].genblk1.mux.sel
+ _00217_ VGND VGND VPWR VPWR _02246_ sky130_fd_sc_hd__and4b_1
XFILLER_0_20_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_130_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11104_ _01193_ _01194_ _01195_ VGND VGND VPWR VPWR _01197_ sky130_fd_sc_hd__and3_1
X_12084_ _02093_ _02096_ VGND VGND VPWR VPWR _02177_ sky130_fd_sc_hd__xor2_1
X_16961_ _02476_ _07105_ VGND VGND VPWR VPWR _07394_ sky130_fd_sc_hd__and2_4
X_18700_ _09209_ _09230_ VGND VGND VPWR VPWR _09231_ sky130_fd_sc_hd__and2_1
X_11035_ _07254_ _05333_ _05039_ _07232_ VGND VGND VPWR VPWR _01128_ sky130_fd_sc_hd__a22o_1
X_15912_ _06254_ _06255_ VGND VGND VPWR VPWR _06257_ sky130_fd_sc_hd__and2_1
X_16892_ _06579_ _07318_ VGND VGND VPWR VPWR _07320_ sky130_fd_sc_hd__or2_1
X_18631_ net34 net67 net68 VGND VGND VPWR VPWR _09178_ sky130_fd_sc_hd__nand3_2
X_15843_ _06180_ _06182_ VGND VGND VPWR VPWR _06183_ sky130_fd_sc_hd__xor2_2
XFILLER_0_91_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18562_ salida\[3\] _09114_ _09118_ salida\[35\] _09128_ VGND VGND VPWR VPWR _09132_
+ sky130_fd_sc_hd__a221o_1
X_15774_ _06100_ _06107_ VGND VGND VPWR VPWR _06108_ sky130_fd_sc_hd__nand2_1
X_12986_ _02780_ VGND VGND VPWR VPWR _03079_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_99_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17513_ _07851_ _07878_ _07996_ VGND VGND VPWR VPWR _07997_ sky130_fd_sc_hd__o21a_1
XFILLER_0_115_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14725_ _04794_ _04796_ _04924_ _04925_ VGND VGND VPWR VPWR _04966_ sky130_fd_sc_hd__o211a_1
X_11937_ _01082_ _01081_ _03826_ _03388_ VGND VGND VPWR VPWR _02030_ sky130_fd_sc_hd__and4_1
X_18493_ _02951_ _09060_ VGND VGND VPWR VPWR _09061_ sky130_fd_sc_hd__nor2_1
X_17444_ _02973_ _07920_ _07921_ _06484_ VGND VGND VPWR VPWR _07922_ sky130_fd_sc_hd__o211a_1
XFILLER_0_28_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14656_ _04887_ _04890_ VGND VGND VPWR VPWR _04891_ sky130_fd_sc_hd__xnor2_2
X_11868_ _01946_ _01959_ VGND VGND VPWR VPWR _01961_ sky130_fd_sc_hd__xnor2_1
X_10819_ _03465_ _00909_ _00910_ _00911_ VGND VGND VPWR VPWR _00912_ sky130_fd_sc_hd__nand4_2
X_13607_ _03358_ _03360_ _03527_ _03528_ _03744_ VGND VGND VPWR VPWR _03745_ sky130_fd_sc_hd__a41o_1
XFILLER_0_7_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17375_ _07039_ _07108_ VGND VGND VPWR VPWR _07846_ sky130_fd_sc_hd__nand2_1
XFILLER_0_27_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14587_ net244 _04686_ _04815_ VGND VGND VPWR VPWR _04816_ sky130_fd_sc_hd__or3_1
X_11799_ _01887_ _01890_ _01707_ _01891_ VGND VGND VPWR VPWR _01892_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_138_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16326_ _06698_ _06704_ _03080_ VGND VGND VPWR VPWR _06705_ sky130_fd_sc_hd__mux2_1
X_13538_ _03667_ _03668_ VGND VGND VPWR VPWR _03669_ sky130_fd_sc_hd__or2b_1
XFILLER_0_131_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13469_ _03629_ _03596_ _05333_ _00439_ VGND VGND VPWR VPWR _03593_ sky130_fd_sc_hd__and4_1
X_16257_ _06617_ _06629_ _04247_ VGND VGND VPWR VPWR _06630_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_679 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_112_214 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15208_ _05375_ _05376_ _05492_ VGND VGND VPWR VPWR _05493_ sky130_fd_sc_hd__o21ai_2
X_16188_ _06516_ _06527_ _06542_ _06554_ VGND VGND VPWR VPWR _06555_ sky130_fd_sc_hd__a31o_1
XFILLER_0_23_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15139_ _05407_ _05416_ VGND VGND VPWR VPWR _05418_ sky130_fd_sc_hd__nand2_1
XFILLER_0_140_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09700_ _06202_ _06224_ _06213_ VGND VGND VPWR VPWR _06245_ sky130_fd_sc_hd__a21o_1
X_09631_ _05028_ VGND VGND VPWR VPWR _05497_ sky130_fd_sc_hd__buf_4
X_18829_ net69 _09116_ _09180_ VGND VGND VPWR VPWR _09331_ sky130_fd_sc_hd__or3_4
X_09562_ _04624_ _04733_ VGND VGND VPWR VPWR _04744_ sky130_fd_sc_hd__xnor2_2
X_09493_ _03717_ VGND VGND VPWR VPWR _03990_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_93_716 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_147_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_226 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_148_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_116_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_143_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_131_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09829_ _07570_ VGND VGND VPWR VPWR _07646_ sky130_fd_sc_hd__clkbuf_4
X_12840_ _00884_ _02921_ _02932_ VGND VGND VPWR VPWR _02933_ sky130_fd_sc_hd__o21a_1
XTAP_2101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12771_ _02860_ _02861_ _02862_ VGND VGND VPWR VPWR _02864_ sky130_fd_sc_hd__o21bai_1
XTAP_2145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14510_ _04576_ _04577_ _04729_ VGND VGND VPWR VPWR _04731_ sky130_fd_sc_hd__or3_1
XFILLER_0_56_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11722_ _01813_ _01814_ _03990_ _09212_ VGND VGND VPWR VPWR _01815_ sky130_fd_sc_hd__and4b_1
XFILLER_0_84_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15490_ _02973_ _03583_ _05799_ VGND VGND VPWR VPWR _05800_ sky130_fd_sc_hd__o21ai_1
XTAP_2189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14441_ _00148_ _00149_ _08452_ _04700_ VGND VGND VPWR VPWR _04656_ sky130_fd_sc_hd__and4_1
XTAP_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11653_ _07646_ VGND VGND VPWR VPWR _01746_ sky130_fd_sc_hd__clkbuf_4
XTAP_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10604_ _00694_ _00695_ _00491_ _00535_ VGND VGND VPWR VPWR _00697_ sky130_fd_sc_hd__o211a_1
X_14372_ _04573_ net178 _04579_ VGND VGND VPWR VPWR _04581_ sky130_fd_sc_hd__nand3_1
XFILLER_0_64_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17160_ _07609_ _07610_ VGND VGND VPWR VPWR _07611_ sky130_fd_sc_hd__and2b_1
X_11584_ _00845_ VGND VGND VPWR VPWR _01677_ sky130_fd_sc_hd__buf_4
XFILLER_0_36_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_326 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_153_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13323_ _03374_ _03264_ _03431_ _03433_ VGND VGND VPWR VPWR _03434_ sky130_fd_sc_hd__o211a_2
X_16111_ _06467_ VGND VGND VPWR VPWR _06470_ sky130_fd_sc_hd__buf_2
X_10535_ _00623_ _00626_ _00627_ VGND VGND VPWR VPWR _00628_ sky130_fd_sc_hd__and3_1
XFILLER_0_24_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17091_ _07483_ _07430_ _07535_ VGND VGND VPWR VPWR _07536_ sky130_fd_sc_hd__o21a_1
XFILLER_0_135_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13254_ _00759_ _00908_ VGND VGND VPWR VPWR _03359_ sky130_fd_sc_hd__and2_1
X_16042_ _06393_ _06394_ _04887_ VGND VGND VPWR VPWR _06396_ sky130_fd_sc_hd__a21bo_1
X_10466_ _00163_ _00558_ VGND VGND VPWR VPWR _00559_ sky130_fd_sc_hd__nand2_1
XFILLER_0_122_556 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12205_ net129 _02294_ _02230_ _02282_ VGND VGND VPWR VPWR _02298_ sky130_fd_sc_hd__o211a_1
XFILLER_0_110_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13185_ _03280_ _03284_ VGND VGND VPWR VPWR _03285_ sky130_fd_sc_hd__xor2_2
XFILLER_0_86_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10397_ _00486_ _00487_ _00488_ _00467_ VGND VGND VPWR VPWR _00490_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12136_ _02198_ _02199_ _02202_ VGND VGND VPWR VPWR _02229_ sky130_fd_sc_hd__a21oi_1
X_17993_ _07084_ _08517_ _08519_ VGND VGND VPWR VPWR _08520_ sky130_fd_sc_hd__or3_1
X_12067_ _02154_ _02158_ _02136_ _02137_ VGND VGND VPWR VPWR _02160_ sky130_fd_sc_hd__o211a_1
X_16944_ _06508_ _07361_ _07362_ _07376_ VGND VGND VPWR VPWR _07377_ sky130_fd_sc_hd__a31o_1
XFILLER_0_19_78 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11018_ _01107_ _01109_ VGND VGND VPWR VPWR _01111_ sky130_fd_sc_hd__nor2_1
X_16875_ _06762_ _06890_ _06947_ _07026_ VGND VGND VPWR VPWR _07301_ sky130_fd_sc_hd__and4_1
X_18614_ salida\[24\] _09159_ _09160_ salida\[56\] _09163_ VGND VGND VPWR VPWR _09168_
+ sky130_fd_sc_hd__a221o_1
X_15826_ _06037_ _05652_ _02992_ VGND VGND VPWR VPWR _06164_ sky130_fd_sc_hd__and3b_1
XFILLER_0_35_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18545_ net28 net148 VGND VGND VPWR VPWR _09116_ sky130_fd_sc_hd__nand2_1
X_15757_ _03012_ _03149_ _03067_ _03010_ VGND VGND VPWR VPWR _06089_ sky130_fd_sc_hd__a22oi_1
X_12969_ _03061_ VGND VGND VPWR VPWR _03062_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_143_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14708_ _04551_ _04691_ _04693_ _04818_ VGND VGND VPWR VPWR _04948_ sky130_fd_sc_hd__or4_4
X_18476_ _08961_ _09036_ _09004_ VGND VGND VPWR VPWR _09042_ sky130_fd_sc_hd__a21o_1
XFILLER_0_129_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15688_ _06013_ _06014_ VGND VGND VPWR VPWR _06015_ sky130_fd_sc_hd__or2_1
XTAP_2690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17427_ _07790_ _07794_ _07791_ VGND VGND VPWR VPWR _07903_ sky130_fd_sc_hd__o21a_4
XFILLER_0_145_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14639_ _04870_ _05921_ _03014_ _04871_ VGND VGND VPWR VPWR _04872_ sky130_fd_sc_hd__and4b_1
XFILLER_0_117_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17358_ _00557_ _07825_ VGND VGND VPWR VPWR _07827_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16309_ _06333_ _06334_ VGND VGND VPWR VPWR _06686_ sky130_fd_sc_hd__and2_1
XFILLER_0_153_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_808 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_141_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17289_ _07207_ _07039_ _07751_ _06947_ VGND VGND VPWR VPWR _07752_ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_141_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09614_ cla_inst.in1\[19\] VGND VGND VPWR VPWR _05311_ sky130_fd_sc_hd__buf_6
XFILLER_0_97_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09545_ _04548_ VGND VGND VPWR VPWR _04558_ sky130_fd_sc_hd__buf_4
XFILLER_0_78_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09476_ ApproximateM_inst.lob_16.lob1.genblk1\[12\].genblk1.mux.sel VGND VGND VPWR
+ VPWR _03804_ sky130_fd_sc_hd__buf_6
XFILLER_0_38_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_136 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire117 _05408_ VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__buf_2
XFILLER_0_18_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire139 _01406_ VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__buf_1
XFILLER_0_135_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10320_ _00411_ _00401_ _00402_ VGND VGND VPWR VPWR _00413_ sky130_fd_sc_hd__or3_1
XFILLER_0_61_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10251_ _07080_ cla_inst.in1\[28\] _07374_ _07047_ VGND VGND VPWR VPWR _00344_ sky130_fd_sc_hd__a22o_1
XFILLER_0_100_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10182_ _03629_ _03596_ _04482_ _03815_ VGND VGND VPWR VPWR _00275_ sky130_fd_sc_hd__nand4_2
X_14990_ _05247_ _05254_ VGND VGND VPWR VPWR _05255_ sky130_fd_sc_hd__xor2_1
X_13941_ _04001_ _07134_ _03941_ _03940_ _00309_ VGND VGND VPWR VPWR _04109_ sky130_fd_sc_hd__a32o_1
XFILLER_0_89_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16660_ _07065_ _07063_ VGND VGND VPWR VPWR _07067_ sky130_fd_sc_hd__or2b_1
X_13872_ cla_inst.in2\[25\] _03750_ VGND VGND VPWR VPWR _04035_ sky130_fd_sc_hd__nand2_1
X_15611_ _05892_ _05929_ _05930_ VGND VGND VPWR VPWR _05931_ sky130_fd_sc_hd__and3_1
X_12823_ _02895_ _02915_ VGND VGND VPWR VPWR _02916_ sky130_fd_sc_hd__xnor2_1
X_16591_ _06990_ _06991_ VGND VGND VPWR VPWR _06992_ sky130_fd_sc_hd__or2_1
XFILLER_0_97_863 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18330_ _07371_ _08141_ _08884_ _06721_ VGND VGND VPWR VPWR _08885_ sky130_fd_sc_hd__o211a_1
X_15542_ _05848_ _05854_ VGND VGND VPWR VPWR _05857_ sky130_fd_sc_hd__nand2_1
XTAP_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12754_ _02462_ _02464_ VGND VGND VPWR VPWR _02847_ sky130_fd_sc_hd__xor2_2
XTAP_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11705_ _01791_ _01797_ VGND VGND VPWR VPWR _01798_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_127_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18261_ _08736_ _08809_ VGND VGND VPWR VPWR _08810_ sky130_fd_sc_hd__xnor2_2
X_15473_ _05596_ _05699_ _05697_ VGND VGND VPWR VPWR _05782_ sky130_fd_sc_hd__a21oi_2
XTAP_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12685_ _02744_ _02752_ _02775_ VGND VGND VPWR VPWR _02778_ sky130_fd_sc_hd__a21oi_1
XTAP_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17212_ _07586_ _07587_ _07667_ VGND VGND VPWR VPWR _07669_ sky130_fd_sc_hd__nor3_1
X_14424_ _04496_ _04631_ _04637_ VGND VGND VPWR VPWR _04638_ sky130_fd_sc_hd__nor3_1
XFILLER_0_71_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11636_ _01221_ _01693_ VGND VGND VPWR VPWR _01729_ sky130_fd_sc_hd__nor2_1
X_18192_ _08660_ _08697_ _08734_ VGND VGND VPWR VPWR _08736_ sky130_fd_sc_hd__o21ba_2
XFILLER_0_21_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17143_ _04725_ _07592_ VGND VGND VPWR VPWR _07593_ sky130_fd_sc_hd__nand2_4
X_11567_ ApproximateM_inst.lob_16.lob2.genblk1\[5\].genblk1.mux.sel _03903_ VGND VGND
+ VPWR VPWR _01660_ sky130_fd_sc_hd__nand2_1
XFILLER_0_107_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14355_ _03164_ _03159_ _04561_ _03916_ VGND VGND VPWR VPWR _04562_ sky130_fd_sc_hd__o211a_1
XFILLER_0_123_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13306_ _05747_ _00513_ VGND VGND VPWR VPWR _03415_ sky130_fd_sc_hd__nand2_1
X_10518_ _00607_ _00608_ _00609_ VGND VGND VPWR VPWR _00611_ sky130_fd_sc_hd__a21o_1
X_14286_ _04470_ _04472_ _04486_ VGND VGND VPWR VPWR _04487_ sky130_fd_sc_hd__a21o_1
XFILLER_0_123_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17074_ _07514_ _07517_ VGND VGND VPWR VPWR _07518_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_24_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11498_ _00806_ _06591_ _00210_ _04220_ VGND VGND VPWR VPWR _01591_ sky130_fd_sc_hd__and4_1
X_13237_ _03337_ _03338_ _03297_ VGND VGND VPWR VPWR _03340_ sky130_fd_sc_hd__a21o_1
XFILLER_0_21_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16025_ _06372_ _06375_ _06376_ VGND VGND VPWR VPWR _06377_ sky130_fd_sc_hd__a21bo_1
X_10449_ _00385_ _00392_ _00541_ VGND VGND VPWR VPWR _00542_ sky130_fd_sc_hd__a21o_1
XFILLER_0_0_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13168_ _00676_ _00689_ VGND VGND VPWR VPWR _03267_ sky130_fd_sc_hd__or2_2
X_12119_ _05638_ _00774_ _00176_ _05562_ VGND VGND VPWR VPWR _02212_ sky130_fd_sc_hd__a22o_1
X_17976_ _08499_ _08500_ VGND VGND VPWR VPWR _08501_ sky130_fd_sc_hd__xor2_1
X_13099_ _03191_ VGND VGND VPWR VPWR _03192_ sky130_fd_sc_hd__inv_2
X_16927_ _07257_ VGND VGND VPWR VPWR _07358_ sky130_fd_sc_hd__inv_2
X_16858_ _02099_ _06723_ _07255_ _07282_ VGND VGND VPWR VPWR _09417_ sky130_fd_sc_hd__o22a_2
X_15809_ _06145_ _03906_ _03907_ _03909_ _02980_ _02978_ VGND VGND VPWR VPWR _06146_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_153_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_149_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16789_ _07026_ VGND VGND VPWR VPWR _07207_ sky130_fd_sc_hd__clkbuf_4
X_18528_ net68 _09096_ VGND VGND VPWR VPWR _09097_ sky130_fd_sc_hd__nor2_4
XFILLER_0_62_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_896 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_146_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18459_ _02938_ _09023_ _03930_ VGND VGND VPWR VPWR _09024_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_7_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_423 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09528_ _04362_ VGND VGND VPWR VPWR _04373_ sky130_fd_sc_hd__buf_6
XPHY_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09459_ _03607_ VGND VGND VPWR VPWR _03618_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_47_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12470_ _01113_ _02099_ VGND VGND VPWR VPWR _02563_ sky130_fd_sc_hd__nor2_2
XFILLER_0_136_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_152_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11421_ _01508_ _01513_ VGND VGND VPWR VPWR _01514_ sky130_fd_sc_hd__or2b_1
XFILLER_0_34_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14140_ _04325_ _04326_ VGND VGND VPWR VPWR _04327_ sky130_fd_sc_hd__and2_1
X_11352_ _01442_ _01443_ _01375_ _01376_ VGND VGND VPWR VPWR _01445_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_104_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_104_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10303_ _00380_ _00381_ _00395_ VGND VGND VPWR VPWR _00396_ sky130_fd_sc_hd__a21o_1
XFILLER_0_120_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14071_ _03199_ _04251_ VGND VGND VPWR VPWR _04252_ sky130_fd_sc_hd__nand2_1
X_11283_ _01267_ _01365_ VGND VGND VPWR VPWR _01376_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13022_ _03106_ _03114_ _03061_ VGND VGND VPWR VPWR _03115_ sky130_fd_sc_hd__mux2_1
X_10234_ _00306_ _00307_ _00325_ VGND VGND VPWR VPWR _00327_ sky130_fd_sc_hd__nand3_1
X_17830_ _03197_ _05625_ _08338_ _08341_ VGND VGND VPWR VPWR _08342_ sky130_fd_sc_hd__a211o_1
X_10165_ _00254_ _00257_ VGND VGND VPWR VPWR _00258_ sky130_fd_sc_hd__xnor2_1
X_17761_ _07751_ net145 VGND VGND VPWR VPWR _08266_ sky130_fd_sc_hd__nand2_1
X_14973_ _05229_ _05236_ VGND VGND VPWR VPWR _05237_ sky130_fd_sc_hd__or2_1
X_10096_ _00173_ VGND VGND VPWR VPWR _00189_ sky130_fd_sc_hd__buf_2
X_16712_ _06951_ VGND VGND VPWR VPWR _07124_ sky130_fd_sc_hd__buf_2
X_13924_ _03962_ VGND VGND VPWR VPWR _04091_ sky130_fd_sc_hd__inv_2
X_17692_ _08189_ _08190_ VGND VGND VPWR VPWR _08192_ sky130_fd_sc_hd__nand2_1
X_16643_ _07017_ _07048_ VGND VGND VPWR VPWR _07049_ sky130_fd_sc_hd__xor2_1
XFILLER_0_16_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13855_ _00204_ _01866_ _04015_ VGND VGND VPWR VPWR _04016_ sky130_fd_sc_hd__nand3_1
XFILLER_0_57_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12806_ _01465_ _01466_ _00854_ _02898_ VGND VGND VPWR VPWR _02899_ sky130_fd_sc_hd__a211o_1
X_16574_ _06749_ _06891_ _06970_ _06972_ VGND VGND VPWR VPWR _06974_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_29_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13786_ _03848_ _03782_ cla_inst.in1\[22\] VGND VGND VPWR VPWR _03940_ sky130_fd_sc_hd__and3_1
X_10998_ _01089_ _01090_ VGND VGND VPWR VPWR _01091_ sky130_fd_sc_hd__and2b_1
XFILLER_0_85_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18313_ _08864_ _08866_ VGND VGND VPWR VPWR _08867_ sky130_fd_sc_hd__xnor2_1
XTAP_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15525_ _05836_ _05837_ VGND VGND VPWR VPWR _05838_ sky130_fd_sc_hd__xor2_1
XFILLER_0_123_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12737_ _02820_ _02828_ _02829_ VGND VGND VPWR VPWR _02830_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_57_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18244_ _08786_ _08790_ VGND VGND VPWR VPWR _08792_ sky130_fd_sc_hd__nand2_1
X_15456_ _05761_ _01317_ _05449_ _05762_ VGND VGND VPWR VPWR _05763_ sky130_fd_sc_hd__and4b_1
XFILLER_0_72_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12668_ _02759_ _02760_ VGND VGND VPWR VPWR _02761_ sky130_fd_sc_hd__or2_1
XFILLER_0_154_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14407_ _04612_ _04616_ _04618_ VGND VGND VPWR VPWR _04619_ sky130_fd_sc_hd__or3_2
XFILLER_0_53_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11619_ _01187_ _01188_ _01191_ VGND VGND VPWR VPWR _01712_ sky130_fd_sc_hd__a21o_1
X_18175_ _07195_ _07861_ _07745_ _07604_ VGND VGND VPWR VPWR _08717_ sky130_fd_sc_hd__o211a_1
X_15387_ _05530_ _05676_ _05687_ VGND VGND VPWR VPWR _05688_ sky130_fd_sc_hd__o21a_1
XFILLER_0_4_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12599_ _02683_ _02691_ VGND VGND VPWR VPWR _02692_ sky130_fd_sc_hd__or2b_1
XFILLER_0_52_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17126_ _02347_ _06920_ _06921_ VGND VGND VPWR VPWR _07575_ sky130_fd_sc_hd__a21o_1
XFILLER_0_13_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14338_ _04423_ _04424_ _04542_ _04543_ VGND VGND VPWR VPWR _04544_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_123_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17057_ _07497_ _07498_ VGND VGND VPWR VPWR _07499_ sky130_fd_sc_hd__xnor2_2
X_14269_ _04461_ _04462_ _04467_ VGND VGND VPWR VPWR _04468_ sky130_fd_sc_hd__nand3_4
XFILLER_0_150_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16008_ _02476_ _00167_ VGND VGND VPWR VPWR _06358_ sky130_fd_sc_hd__and2_1
XTAP_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17959_ _08363_ _08450_ _08481_ VGND VGND VPWR VPWR _08482_ sky130_fd_sc_hd__a21o_1
XFILLER_0_73_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_800 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_137_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11970_ _02022_ _02016_ _02021_ VGND VGND VPWR VPWR _02063_ sky130_fd_sc_hd__nor3_1
X_10921_ _00998_ _00999_ _01013_ VGND VGND VPWR VPWR _01014_ sky130_fd_sc_hd__a21o_2
X_13640_ _03778_ _03779_ VGND VGND VPWR VPWR _03780_ sky130_fd_sc_hd__nor2_1
X_10852_ ApproximateM_inst.lob_16.lob2.genblk1\[12\].genblk1.mux.sel net209 _03388_
+ _04493_ VGND VGND VPWR VPWR _00945_ sky130_fd_sc_hd__a22o_1
XFILLER_0_94_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13571_ _03703_ _03704_ VGND VGND VPWR VPWR _03705_ sky130_fd_sc_hd__nor2_1
X_10783_ _00870_ _00875_ VGND VGND VPWR VPWR _00876_ sky130_fd_sc_hd__and2b_1
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15310_ _05503_ _05506_ _05603_ VGND VGND VPWR VPWR _05604_ sky130_fd_sc_hd__a21oi_1
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12522_ _02604_ _02613_ net137 _02614_ VGND VGND VPWR VPWR _02615_ sky130_fd_sc_hd__a211o_1
XFILLER_0_82_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16290_ _06664_ VGND VGND VPWR VPWR _06665_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_137_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_151_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15241_ _05320_ _05439_ VGND VGND VPWR VPWR _05528_ sky130_fd_sc_hd__and2_1
X_12453_ _05638_ ApproximateM_inst.lob_16.lob1.genblk1\[1\].genblk1.mux.sel _07581_
+ _05562_ VGND VGND VPWR VPWR _02546_ sky130_fd_sc_hd__a22o_1
XFILLER_0_152_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11404_ _01494_ _01495_ _01451_ _01444_ VGND VGND VPWR VPWR _01497_ sky130_fd_sc_hd__o211a_1
XFILLER_0_105_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15172_ _05444_ _05451_ VGND VGND VPWR VPWR _05454_ sky130_fd_sc_hd__nand2_1
XFILLER_0_50_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12384_ _05834_ _00357_ _07657_ _02476_ VGND VGND VPWR VPWR _02477_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_105_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14123_ _04302_ _04117_ _04308_ VGND VGND VPWR VPWR _04309_ sky130_fd_sc_hd__o21a_1
X_11335_ _01426_ _01427_ VGND VGND VPWR VPWR _01428_ sky130_fd_sc_hd__xnor2_2
X_18931_ clknet_4_12_0_clk _00085_ VGND VGND VPWR VPWR cla_inst.in2\[17\] sky130_fd_sc_hd__dfxtp_2
X_11266_ _01356_ VGND VGND VPWR VPWR _01359_ sky130_fd_sc_hd__clkbuf_8
X_14054_ _04061_ _04060_ VGND VGND VPWR VPWR _04234_ sky130_fd_sc_hd__or2b_1
X_10217_ _08724_ _00309_ VGND VGND VPWR VPWR _00310_ sky130_fd_sc_hd__nand2_1
XFILLER_0_120_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13005_ _02489_ VGND VGND VPWR VPWR _03098_ sky130_fd_sc_hd__buf_4
X_18862_ clknet_4_5_0_clk net288 VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__dfxtp_1
X_11197_ _00967_ _01274_ _01288_ _01289_ VGND VGND VPWR VPWR _01290_ sky130_fd_sc_hd__o211a_2
XFILLER_0_94_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17813_ _08253_ _08254_ _08323_ VGND VGND VPWR VPWR _08324_ sky130_fd_sc_hd__nand3_1
X_10148_ _07624_ _00240_ VGND VGND VPWR VPWR _00241_ sky130_fd_sc_hd__xnor2_1
X_18793_ _09304_ VGND VGND VPWR VPWR _00088_ sky130_fd_sc_hd__buf_1
XFILLER_0_89_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17744_ _08225_ _08229_ _08248_ _06723_ _01671_ VGND VGND VPWR VPWR _09395_ sky130_fd_sc_hd__o32a_1
X_14956_ _05216_ _05217_ VGND VGND VPWR VPWR _05218_ sky130_fd_sc_hd__xor2_1
X_10079_ _00171_ VGND VGND VPWR VPWR _00172_ sky130_fd_sc_hd__buf_4
X_13907_ _04068_ _04071_ VGND VGND VPWR VPWR _04073_ sky130_fd_sc_hd__nand2_1
X_17675_ _08057_ _08058_ VGND VGND VPWR VPWR _08173_ sky130_fd_sc_hd__or2_1
X_14887_ _05021_ _05023_ VGND VGND VPWR VPWR _05143_ sky130_fd_sc_hd__nand2_1
X_16626_ _07028_ _07029_ VGND VGND VPWR VPWR _07030_ sky130_fd_sc_hd__xnor2_1
X_13838_ _03805_ _03807_ _03996_ VGND VGND VPWR VPWR _03997_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_134_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16557_ _04449_ _04471_ _03184_ VGND VGND VPWR VPWR _06955_ sky130_fd_sc_hd__o21a_1
X_13769_ _03916_ _03917_ _03919_ _03921_ VGND VGND VPWR VPWR _03922_ sky130_fd_sc_hd__a211o_1
XFILLER_0_45_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15508_ _05813_ _05817_ _05818_ VGND VGND VPWR VPWR _05819_ sky130_fd_sc_hd__and3_1
XFILLER_0_57_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16488_ _06878_ _06879_ _00194_ VGND VGND VPWR VPWR _06880_ sky130_fd_sc_hd__a21bo_2
XFILLER_0_45_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18227_ _08739_ _08749_ VGND VGND VPWR VPWR _08773_ sky130_fd_sc_hd__and2b_1
X_15439_ _02998_ _03153_ VGND VGND VPWR VPWR _05744_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_251 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18158_ _07751_ _08150_ _08625_ _08540_ VGND VGND VPWR VPWR _08698_ sky130_fd_sc_hd__a31o_1
X_17109_ _07554_ _07555_ VGND VGND VPWR VPWR _07556_ sky130_fd_sc_hd__xnor2_1
X_18089_ _00558_ _07390_ _08621_ VGND VGND VPWR VPWR _08623_ sky130_fd_sc_hd__a21o_1
XFILLER_0_13_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09931_ _08746_ VGND VGND VPWR VPWR _08757_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_7_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09862_ _06982_ _07962_ _07951_ _07995_ VGND VGND VPWR VPWR _08006_ sky130_fd_sc_hd__nand4_1
XTAP_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09793_ _07243_ VGND VGND VPWR VPWR _07254_ sky130_fd_sc_hd__buf_4
XTAP_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_134_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_134_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11120_ _05682_ _04700_ _01211_ _01212_ VGND VGND VPWR VPWR _01213_ sky130_fd_sc_hd__a31o_1
X_11051_ _01134_ _01143_ VGND VGND VPWR VPWR _01144_ sky130_fd_sc_hd__nand2_1
XFILLER_0_102_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10002_ _07482_ _07908_ _09339_ _09340_ VGND VGND VPWR VPWR _09345_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_99_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14810_ _05056_ _05057_ _05058_ VGND VGND VPWR VPWR _05059_ sky130_fd_sc_hd__and3_1
X_15790_ _06097_ _06123_ VGND VGND VPWR VPWR _06125_ sky130_fd_sc_hd__or2_1
X_14741_ _04975_ _04976_ _04981_ VGND VGND VPWR VPWR _04983_ sky130_fd_sc_hd__a21o_1
Xwb_buttons_leds_151 VGND VGND VPWR VPWR wb_buttons_leds_151/HI led_enb[0] sky130_fd_sc_hd__conb_1
X_11953_ _01106_ _00515_ _02044_ _02045_ VGND VGND VPWR VPWR _02046_ sky130_fd_sc_hd__or4_4
Xwb_buttons_leds_162 VGND VGND VPWR VPWR wb_buttons_leds_162/HI led_enb[11] sky130_fd_sc_hd__conb_1
XFILLER_0_98_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10904_ _00990_ _00996_ VGND VGND VPWR VPWR _00997_ sky130_fd_sc_hd__and2_1
X_17460_ _07936_ _07937_ VGND VGND VPWR VPWR _07938_ sky130_fd_sc_hd__xnor2_2
X_14672_ _00125_ _00443_ _05050_ _00151_ VGND VGND VPWR VPWR _04909_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_58_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11884_ _01871_ _01888_ _01889_ _01887_ VGND VGND VPWR VPWR _01977_ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16411_ _06508_ _06783_ _06784_ _06796_ VGND VGND VPWR VPWR _06797_ sky130_fd_sc_hd__a31o_1
X_13623_ _03758_ _03759_ net226 _03754_ VGND VGND VPWR VPWR _03762_ sky130_fd_sc_hd__a211o_1
X_10835_ _03771_ ApproximateM_inst.lob_16.lob1.genblk1\[7\].genblk1.mux.sel ApproximateM_inst.lob_16.lob1.genblk1\[6\].genblk1.mux.sel
+ cla_inst.in2\[16\] VGND VGND VPWR VPWR _00928_ sky130_fd_sc_hd__a22o_1
XFILLER_0_104_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17391_ _07860_ _07862_ VGND VGND VPWR VPWR _07863_ sky130_fd_sc_hd__and2_1
XFILLER_0_27_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16342_ _06721_ VGND VGND VPWR VPWR _06723_ sky130_fd_sc_hd__clkbuf_4
X_13554_ _03685_ _03686_ VGND VGND VPWR VPWR _03687_ sky130_fd_sc_hd__or2_1
X_10766_ _00857_ _00858_ VGND VGND VPWR VPWR _00859_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_54_335 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12505_ _02595_ _02597_ VGND VGND VPWR VPWR _02598_ sky130_fd_sc_hd__nand2_1
XFILLER_0_152_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16273_ _06559_ _06583_ _06584_ _06608_ _06647_ VGND VGND VPWR VPWR _06648_ sky130_fd_sc_hd__o311a_1
X_13485_ _00294_ cla_inst.in1\[24\] _05693_ _04504_ VGND VGND VPWR VPWR _03611_ sky130_fd_sc_hd__a22o_1
X_10697_ _04548_ _04482_ VGND VGND VPWR VPWR _00790_ sky130_fd_sc_hd__nand2_2
XFILLER_0_82_688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18012_ _07035_ _07933_ _08538_ VGND VGND VPWR VPWR _08540_ sky130_fd_sc_hd__or3b_2
X_15224_ _05428_ _05396_ _05509_ VGND VGND VPWR VPWR _05511_ sky130_fd_sc_hd__and3_1
XFILLER_0_63_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12436_ _02471_ _02528_ VGND VGND VPWR VPWR _02529_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_22_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15155_ _02987_ _03456_ _00513_ _02985_ VGND VGND VPWR VPWR _05435_ sky130_fd_sc_hd__a22o_1
XFILLER_0_140_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12367_ _02452_ _02458_ _02459_ VGND VGND VPWR VPWR _02460_ sky130_fd_sc_hd__or3_1
X_14106_ _04558_ _09248_ _04288_ _04289_ VGND VGND VPWR VPWR _04290_ sky130_fd_sc_hd__and4_1
X_11318_ _01410_ _01329_ VGND VGND VPWR VPWR _01411_ sky130_fd_sc_hd__or2_1
X_15086_ _05237_ _05359_ VGND VGND VPWR VPWR _05360_ sky130_fd_sc_hd__xnor2_1
X_12298_ _02295_ _02298_ _02297_ VGND VGND VPWR VPWR _02391_ sky130_fd_sc_hd__o21ai_1
X_14037_ _04212_ _04213_ _03997_ _04173_ VGND VGND VPWR VPWR _04215_ sky130_fd_sc_hd__a211oi_1
X_11249_ cla_inst.in2\[24\] _00174_ _00871_ _09179_ VGND VGND VPWR VPWR _01342_ sky130_fd_sc_hd__nand4_1
X_18914_ clknet_4_9_0_clk _00068_ VGND VGND VPWR VPWR ApproximateM_inst.lob_16.lob2.mux.sel
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_129_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18845_ clknet_4_1_0_clk net274 VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__dfxtp_1
X_18776_ _09290_ VGND VGND VPWR VPWR _00083_ sky130_fd_sc_hd__buf_1
X_15988_ _02977_ _00134_ VGND VGND VPWR VPWR _06336_ sky130_fd_sc_hd__or2_2
X_17727_ _02987_ _06511_ _01671_ VGND VGND VPWR VPWR _08230_ sky130_fd_sc_hd__a21o_1
XFILLER_0_54_54 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14939_ _05199_ _05077_ VGND VGND VPWR VPWR _05200_ sky130_fd_sc_hd__nor2_1
XFILLER_0_77_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_148_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17658_ _02200_ _06891_ VGND VGND VPWR VPWR _08154_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_298 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16609_ _02829_ _02820_ VGND VGND VPWR VPWR _07012_ sky130_fd_sc_hd__xor2_1
XFILLER_0_148_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17589_ _08065_ _08078_ VGND VGND VPWR VPWR _08079_ sky130_fd_sc_hd__xor2_1
XFILLER_0_147_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold100 net100 VGND VGND VPWR VPWR net263 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold111 _00011_ VGND VGND VPWR VPWR net274 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_574 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold122 net88 VGND VGND VPWR VPWR net285 sky130_fd_sc_hd__dlygate4sd3_1
Xhold133 _00004_ VGND VGND VPWR VPWR net296 sky130_fd_sc_hd__dlygate4sd3_1
Xhold144 _00014_ VGND VGND VPWR VPWR net307 sky130_fd_sc_hd__dlygate4sd3_1
Xhold155 op_code\[3\] VGND VGND VPWR VPWR net318 sky130_fd_sc_hd__clkbuf_2
X_09914_ _04438_ _05388_ _05497_ _04646_ VGND VGND VPWR VPWR _08572_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09845_ _07788_ _07384_ _07810_ VGND VGND VPWR VPWR _07820_ sky130_fd_sc_hd__and3_1
XTAP_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09776_ ApproximateM_inst.lob_16.lob2.genblk1\[3\].genblk1.mux.sel VGND VGND VPWR
+ VPWR _07069_ sky130_fd_sc_hd__buf_6
XTAP_2305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10620_ _00700_ _00701_ _00711_ VGND VGND VPWR VPWR _00713_ sky130_fd_sc_hd__and3_1
XFILLER_0_63_132 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10551_ _05453_ VGND VGND VPWR VPWR _00644_ sky130_fd_sc_hd__buf_4
XFILLER_0_119_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13270_ _03224_ _03225_ _03236_ VGND VGND VPWR VPWR _03375_ sky130_fd_sc_hd__nor3_1
X_10482_ _00559_ _00574_ VGND VGND VPWR VPWR _00575_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_134_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12221_ _02302_ _02304_ _02305_ VGND VGND VPWR VPWR _02314_ sky130_fd_sc_hd__nor3_1
XFILLER_0_122_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12152_ _05584_ net206 _00179_ _05562_ VGND VGND VPWR VPWR _02245_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11103_ _01193_ _01194_ _01195_ VGND VGND VPWR VPWR _01196_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_102_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12083_ _02175_ _01999_ VGND VGND VPWR VPWR _02176_ sky130_fd_sc_hd__nor2_1
X_16960_ _06571_ _06653_ _07194_ _07290_ VGND VGND VPWR VPWR _07393_ sky130_fd_sc_hd__or4_2
X_11034_ _07232_ _07254_ _05333_ _05039_ VGND VGND VPWR VPWR _01127_ sky130_fd_sc_hd__nand4_2
X_15911_ _06244_ _06253_ VGND VGND VPWR VPWR _06255_ sky130_fd_sc_hd__or2_1
X_16891_ _07218_ VGND VGND VPWR VPWR _07318_ sky130_fd_sc_hd__clkbuf_4
X_18630_ net310 _09097_ _09177_ _09176_ VGND VGND VPWR VPWR _00035_ sky130_fd_sc_hd__o211a_1
X_15842_ _06128_ _06131_ VGND VGND VPWR VPWR _06182_ sky130_fd_sc_hd__nand2_1
X_18561_ net311 _09098_ _09130_ _09126_ VGND VGND VPWR VPWR _00006_ sky130_fd_sc_hd__o211a_1
X_15773_ _06104_ _06106_ VGND VGND VPWR VPWR _06107_ sky130_fd_sc_hd__and2_1
X_12985_ _03066_ _03076_ _03077_ VGND VGND VPWR VPWR _03078_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17512_ _07970_ _07994_ VGND VGND VPWR VPWR _07996_ sky130_fd_sc_hd__xnor2_1
X_14724_ _04924_ VGND VGND VPWR VPWR _04965_ sky130_fd_sc_hd__inv_2
X_11936_ _01081_ _03826_ _03399_ _01082_ VGND VGND VPWR VPWR _02029_ sky130_fd_sc_hd__a22o_1
X_18492_ _02939_ net115 _02960_ VGND VGND VPWR VPWR _09060_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_59_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17443_ _03080_ _03062_ _06724_ _03536_ VGND VGND VPWR VPWR _07921_ sky130_fd_sc_hd__a31o_1
X_14655_ _04888_ _04889_ VGND VGND VPWR VPWR _04890_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11867_ _01946_ _01959_ VGND VGND VPWR VPWR _01960_ sky130_fd_sc_hd__or2_1
XFILLER_0_129_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_129_359 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13606_ _03527_ _03743_ VGND VGND VPWR VPWR _03744_ sky130_fd_sc_hd__nand2_1
X_10818_ cla_inst.in2\[17\] ApproximateM_inst.lob_16.lob1.genblk1\[6\].genblk1.mux.sel
+ _00179_ _03520_ VGND VGND VPWR VPWR _00911_ sky130_fd_sc_hd__a22o_1
X_17374_ _07042_ _07721_ _07844_ VGND VGND VPWR VPWR _07845_ sky130_fd_sc_hd__o21ba_1
X_14586_ _04812_ _04814_ VGND VGND VPWR VPWR _04815_ sky130_fd_sc_hd__xnor2_1
X_11798_ _01704_ _01705_ _01706_ _01642_ VGND VGND VPWR VPWR _01891_ sky130_fd_sc_hd__o22a_1
XFILLER_0_28_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16325_ _06701_ _06703_ _03060_ VGND VGND VPWR VPWR _06704_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13537_ _03426_ _03428_ _03666_ VGND VGND VPWR VPWR _03668_ sky130_fd_sc_hd__or3b_1
XFILLER_0_153_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10749_ _06971_ _06722_ _07951_ _07995_ VGND VGND VPWR VPWR _00842_ sky130_fd_sc_hd__and4_1
XFILLER_0_54_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16256_ _06621_ _06628_ _03099_ VGND VGND VPWR VPWR _06629_ sky130_fd_sc_hd__mux2_1
X_13468_ _03589_ net225 _03588_ VGND VGND VPWR VPWR _03592_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_140_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_738 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15207_ _05374_ _05373_ VGND VGND VPWR VPWR _05492_ sky130_fd_sc_hd__or2b_1
XFILLER_0_23_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12419_ _02414_ _02511_ VGND VGND VPWR VPWR _02512_ sky130_fd_sc_hd__and2_1
XFILLER_0_112_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16187_ _06477_ _03029_ _06543_ _06546_ _06553_ VGND VGND VPWR VPWR _06554_ sky130_fd_sc_hd__o32a_2
X_13399_ _03469_ _03470_ _03514_ _03515_ VGND VGND VPWR VPWR _03517_ sky130_fd_sc_hd__a22o_1
XFILLER_0_112_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15138_ _05407_ _05416_ VGND VGND VPWR VPWR _05417_ sky130_fd_sc_hd__or2_1
X_15069_ _05339_ _05340_ VGND VGND VPWR VPWR _05341_ sky130_fd_sc_hd__and2_1
XFILLER_0_65_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09630_ _05322_ VGND VGND VPWR VPWR _05486_ sky130_fd_sc_hd__buf_4
X_18828_ net27 net28 _09109_ _09330_ VGND VGND VPWR VPWR _00100_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_65_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09561_ _04668_ _04722_ VGND VGND VPWR VPWR _04733_ sky130_fd_sc_hd__and2b_1
X_18759_ _00644_ net36 _09276_ VGND VGND VPWR VPWR _09277_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09492_ _03706_ _03957_ _03946_ VGND VGND VPWR VPWR _03979_ sky130_fd_sc_hd__a21o_1
XFILLER_0_66_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_362 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09828_ _07537_ VGND VGND VPWR VPWR _07635_ sky130_fd_sc_hd__clkbuf_4
X_09759_ _06526_ _06537_ _04973_ _06191_ VGND VGND VPWR VPWR _06884_ sky130_fd_sc_hd__o211ai_1
XTAP_2102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12770_ _02860_ _02861_ _02862_ VGND VGND VPWR VPWR _02863_ sky130_fd_sc_hd__or3b_1
XFILLER_0_96_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11721_ _03782_ _09179_ _07581_ _03848_ VGND VGND VPWR VPWR _01814_ sky130_fd_sc_hd__a22o_1
XFILLER_0_68_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_599 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14440_ _03321_ _04591_ _01005_ _00112_ VGND VGND VPWR VPWR _04655_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_49_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11652_ _00204_ VGND VGND VPWR VPWR _01745_ sky130_fd_sc_hd__buf_4
XTAP_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10603_ _00491_ _00535_ net164 _00695_ VGND VGND VPWR VPWR _00696_ sky130_fd_sc_hd__a211oi_4
X_14371_ _04577_ _04578_ VGND VGND VPWR VPWR _04579_ sky130_fd_sc_hd__nor2_2
XFILLER_0_153_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11583_ _01673_ _01675_ VGND VGND VPWR VPWR _01676_ sky130_fd_sc_hd__nor2_1
XFILLER_0_135_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16110_ _02983_ _02257_ _03181_ _06467_ _06468_ VGND VGND VPWR VPWR _06469_ sky130_fd_sc_hd__o311a_1
X_13322_ _03408_ _03409_ _03429_ _03430_ VGND VGND VPWR VPWR _03433_ sky130_fd_sc_hd__nand4_4
XFILLER_0_24_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10534_ _05017_ _05964_ _00624_ _00625_ VGND VGND VPWR VPWR _00627_ sky130_fd_sc_hd__a22o_1
X_17090_ _07533_ _07534_ VGND VGND VPWR VPWR _07535_ sky130_fd_sc_hd__nor2_1
XFILLER_0_150_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16041_ _02998_ _04647_ VGND VGND VPWR VPWR _06394_ sky130_fd_sc_hd__or2_1
XFILLER_0_134_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13253_ _03355_ _03357_ VGND VGND VPWR VPWR _03358_ sky130_fd_sc_hd__and2_1
X_10465_ _00557_ VGND VGND VPWR VPWR _00558_ sky130_fd_sc_hd__buf_4
XFILLER_0_122_568 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12204_ _02274_ _02296_ VGND VGND VPWR VPWR _02297_ sky130_fd_sc_hd__xor2_1
X_10396_ _00467_ _00486_ _00487_ _00488_ VGND VGND VPWR VPWR _00489_ sky130_fd_sc_hd__nand4_2
X_13184_ _03282_ _03283_ VGND VGND VPWR VPWR _03284_ sky130_fd_sc_hd__xor2_2
XFILLER_0_20_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12135_ _02224_ _02225_ _02227_ VGND VGND VPWR VPWR _02228_ sky130_fd_sc_hd__or3_2
X_17992_ _04630_ _06392_ _06391_ VGND VGND VPWR VPWR _08519_ sky130_fd_sc_hd__a21oi_1
X_16943_ _03198_ _04559_ _07365_ _07375_ VGND VGND VPWR VPWR _07376_ sky130_fd_sc_hd__a211o_1
X_12066_ _02136_ _02137_ _02154_ _02158_ VGND VGND VPWR VPWR _02159_ sky130_fd_sc_hd__a211oi_1
X_11017_ _01107_ _01109_ VGND VGND VPWR VPWR _01110_ sky130_fd_sc_hd__and2_1
X_16874_ _07298_ _07299_ VGND VGND VPWR VPWR _07300_ sky130_fd_sc_hd__nand2_1
X_15825_ _03016_ _03072_ _06091_ _06090_ VGND VGND VPWR VPWR _06163_ sky130_fd_sc_hd__a31o_1
X_18613_ net281 _09157_ _09167_ _09162_ VGND VGND VPWR VPWR _00027_ sky130_fd_sc_hd__o211a_1
X_18544_ net13 net2 net24 VGND VGND VPWR VPWR _09115_ sky130_fd_sc_hd__or3b_4
X_15756_ _03007_ _03142_ VGND VGND VPWR VPWR _06088_ sky130_fd_sc_hd__nand2_1
XFILLER_0_87_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12968_ _03060_ VGND VGND VPWR VPWR _03061_ sky130_fd_sc_hd__buf_4
XFILLER_0_48_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14707_ _04691_ _04692_ _04816_ _04817_ VGND VGND VPWR VPWR _04947_ sky130_fd_sc_hd__and4b_1
XFILLER_0_75_706 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11919_ ApproximateM_inst.lob_16.lob2.genblk1\[10\].genblk1.mux.sel _05290_ net207
+ _00179_ VGND VGND VPWR VPWR _02012_ sky130_fd_sc_hd__and4_1
X_18475_ _09038_ _09040_ VGND VGND VPWR VPWR _09041_ sky130_fd_sc_hd__xnor2_1
X_15687_ _05938_ _05941_ _06012_ VGND VGND VPWR VPWR _06014_ sky130_fd_sc_hd__a21oi_1
XTAP_2680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12899_ _02991_ VGND VGND VPWR VPWR _02992_ sky130_fd_sc_hd__buf_2
XFILLER_0_129_134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17426_ _07900_ _07901_ VGND VGND VPWR VPWR _07902_ sky130_fd_sc_hd__and2b_1
X_14638_ _07515_ _01962_ _01575_ _03008_ VGND VGND VPWR VPWR _04871_ sky130_fd_sc_hd__a22o_1
XTAP_1990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17357_ _07657_ net168 _07825_ VGND VGND VPWR VPWR _07826_ sky130_fd_sc_hd__and3_1
X_14569_ _04775_ _04794_ _04795_ VGND VGND VPWR VPWR _04796_ sky130_fd_sc_hd__nor3_2
XFILLER_0_83_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16308_ _02980_ _01503_ VGND VGND VPWR VPWR _06685_ sky130_fd_sc_hd__nand2_1
XFILLER_0_125_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17288_ _06871_ _07032_ _00213_ VGND VGND VPWR VPWR _07751_ sky130_fd_sc_hd__a21boi_4
XFILLER_0_70_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16239_ _03064_ _06609_ _03089_ VGND VGND VPWR VPWR _06610_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09613_ _05290_ VGND VGND VPWR VPWR _05301_ sky130_fd_sc_hd__buf_4
X_09544_ ApproximateM_inst.lob_16.lob2.genblk1\[11\].genblk1.mux.sel VGND VGND VPWR
+ VPWR _04548_ sky130_fd_sc_hd__buf_4
XFILLER_0_39_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09475_ _03782_ VGND VGND VPWR VPWR _03793_ sky130_fd_sc_hd__buf_6
XFILLER_0_93_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_783 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_117_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_658 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10250_ _07232_ _07254_ cla_inst.in1\[28\] _07374_ VGND VGND VPWR VPWR _00343_ sky130_fd_sc_hd__and4_1
X_10181_ _09027_ _09341_ _09345_ _09343_ VGND VGND VPWR VPWR _00274_ sky130_fd_sc_hd__or4b_4
XFILLER_0_100_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13940_ _04092_ _03945_ _04106_ VGND VGND VPWR VPWR _04108_ sky130_fd_sc_hd__nor3_1
X_13871_ _04031_ _04032_ VGND VGND VPWR VPWR _04033_ sky130_fd_sc_hd__nor2_2
XFILLER_0_69_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15610_ _05927_ _05928_ _05828_ _05893_ VGND VGND VPWR VPWR _05930_ sky130_fd_sc_hd__a211o_1
X_12822_ _02913_ _02914_ VGND VGND VPWR VPWR _02915_ sky130_fd_sc_hd__and2_1
X_16590_ _06908_ _06910_ _06909_ VGND VGND VPWR VPWR _06991_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_96_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15541_ _05848_ _05854_ VGND VGND VPWR VPWR _05855_ sky130_fd_sc_hd__or2_1
XTAP_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_875 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_96_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12753_ _02529_ _02589_ _02844_ _02845_ VGND VGND VPWR VPWR _02846_ sky130_fd_sc_hd__o31ai_4
XTAP_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11704_ _01795_ _01796_ VGND VGND VPWR VPWR _01797_ sky130_fd_sc_hd__and2_1
X_18260_ _08807_ _08808_ VGND VGND VPWR VPWR _08809_ sky130_fd_sc_hd__and2_1
X_15472_ _05778_ _05779_ VGND VGND VPWR VPWR _05781_ sky130_fd_sc_hd__or2_1
XTAP_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12684_ _02710_ _02745_ VGND VGND VPWR VPWR _02777_ sky130_fd_sc_hd__xor2_1
XTAP_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_424 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17211_ _07663_ _07666_ VGND VGND VPWR VPWR _07667_ sky130_fd_sc_hd__xnor2_1
X_14423_ _04634_ _04636_ VGND VGND VPWR VPWR _04637_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_127_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11635_ _07853_ _00461_ _01220_ VGND VGND VPWR VPWR _01728_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_112_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18191_ _08655_ _08733_ VGND VGND VPWR VPWR _08734_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_37_474 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_112_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17142_ _06889_ VGND VGND VPWR VPWR _07592_ sky130_fd_sc_hd__buf_4
X_14354_ _03164_ _03163_ VGND VGND VPWR VPWR _04561_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11566_ _06008_ ApproximateM_inst.lob_16.lob2.genblk1\[6\].genblk1.mux.sel ApproximateM_inst.lob_16.lob1.genblk1\[11\].genblk1.mux.sel
+ VGND VGND VPWR VPWR _01659_ sky130_fd_sc_hd__and3_1
XFILLER_0_13_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_123_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13305_ _09311_ _03412_ _03413_ VGND VGND VPWR VPWR _03414_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_150_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10517_ _00607_ _00608_ _00609_ VGND VGND VPWR VPWR _00610_ sky130_fd_sc_hd__nand3_1
X_17073_ _06581_ _07516_ VGND VGND VPWR VPWR _07517_ sky130_fd_sc_hd__nor2_1
XFILLER_0_12_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14285_ _04484_ _04485_ VGND VGND VPWR VPWR _04486_ sky130_fd_sc_hd__and2_1
XFILLER_0_150_652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11497_ _06591_ _00210_ _03607_ _05399_ VGND VGND VPWR VPWR _01590_ sky130_fd_sc_hd__a22o_1
XFILLER_0_123_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16024_ _06374_ _03107_ VGND VGND VPWR VPWR _06376_ sky130_fd_sc_hd__nand2_1
X_13236_ _03297_ _03337_ _03338_ VGND VGND VPWR VPWR _03339_ sky130_fd_sc_hd__nand3_4
X_10448_ _00386_ _00391_ VGND VGND VPWR VPWR _00541_ sky130_fd_sc_hd__and2b_1
XFILLER_0_21_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13167_ _03263_ _03264_ _00634_ _00660_ VGND VGND VPWR VPWR _03266_ sky130_fd_sc_hd__o211a_2
X_10379_ _08713_ _06732_ _00470_ _00471_ VGND VGND VPWR VPWR _00472_ sky130_fd_sc_hd__and4_2
XFILLER_0_21_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12118_ _05562_ _05584_ _04242_ net206 VGND VGND VPWR VPWR _02211_ sky130_fd_sc_hd__and4_1
X_17975_ _08381_ _08396_ _08394_ VGND VGND VPWR VPWR _08500_ sky130_fd_sc_hd__a21o_1
X_13098_ _03185_ _03190_ _02489_ VGND VGND VPWR VPWR _03191_ sky130_fd_sc_hd__mux2_1
X_12049_ _02058_ _02141_ VGND VGND VPWR VPWR _02142_ sky130_fd_sc_hd__xnor2_1
X_16926_ _07289_ _00248_ _06673_ VGND VGND VPWR VPWR _07357_ sky130_fd_sc_hd__or3_2
XFILLER_0_137_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16857_ _07256_ _07261_ _07262_ _07279_ _07281_ VGND VGND VPWR VPWR _07282_ sky130_fd_sc_hd__a311o_1
X_15808_ _03054_ _03058_ _03050_ VGND VGND VPWR VPWR _06145_ sky130_fd_sc_hd__mux2_1
X_16788_ _06652_ _06764_ _06944_ _07115_ VGND VGND VPWR VPWR _07206_ sky130_fd_sc_hd__or4_1
XFILLER_0_153_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15739_ _06068_ _06069_ VGND VGND VPWR VPWR _06070_ sky130_fd_sc_hd__nor2_1
XFILLER_0_75_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18527_ net34 net67 VGND VGND VPWR VPWR _09096_ sky130_fd_sc_hd__nand2_1
X_18458_ _02920_ _08985_ _02918_ VGND VGND VPWR VPWR _09023_ sky130_fd_sc_hd__o21a_1
XFILLER_0_8_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17409_ _07881_ _07882_ VGND VGND VPWR VPWR _07883_ sky130_fd_sc_hd__and2_1
XFILLER_0_16_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18389_ _07743_ _08947_ VGND VGND VPWR VPWR _08948_ sky130_fd_sc_hd__or2_1
XFILLER_0_28_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_606 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09527_ ApproximateM_inst.lob_16.lob2.genblk1\[12\].genblk1.mux.sel VGND VGND VPWR
+ VPWR _04362_ sky130_fd_sc_hd__buf_4
XFILLER_0_149_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09458_ ApproximateM_inst.lob_16.lob1.genblk1\[7\].genblk1.mux.sel VGND VGND VPWR
+ VPWR _03607_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_93_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11420_ _01511_ _01512_ VGND VGND VPWR VPWR _01513_ sky130_fd_sc_hd__xor2_1
XFILLER_0_62_742 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_117_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11351_ _01375_ _01376_ _01442_ _01443_ VGND VGND VPWR VPWR _01444_ sky130_fd_sc_hd__a211o_1
XFILLER_0_61_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10302_ _00383_ _00394_ VGND VGND VPWR VPWR _00395_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_104_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14070_ _03539_ _04248_ _04250_ VGND VGND VPWR VPWR _04251_ sky130_fd_sc_hd__o21ai_1
X_11282_ _01362_ _01338_ _01363_ VGND VGND VPWR VPWR _01375_ sky130_fd_sc_hd__or3_1
XFILLER_0_120_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13021_ _03110_ _03113_ _03090_ VGND VGND VPWR VPWR _03114_ sky130_fd_sc_hd__mux2_1
X_10233_ _00306_ _00307_ _00325_ VGND VGND VPWR VPWR _00326_ sky130_fd_sc_hd__a21o_2
XFILLER_0_120_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10164_ _00255_ _00256_ VGND VGND VPWR VPWR _00257_ sky130_fd_sc_hd__and2b_1
X_14972_ _05233_ _05234_ VGND VGND VPWR VPWR _05236_ sky130_fd_sc_hd__xor2_1
X_10095_ _00186_ _00187_ VGND VGND VPWR VPWR _00188_ sky130_fd_sc_hd__or2_1
X_17760_ _08263_ _08264_ VGND VGND VPWR VPWR _08265_ sky130_fd_sc_hd__xnor2_1
X_13923_ _03368_ _01678_ _04021_ VGND VGND VPWR VPWR _04090_ sky130_fd_sc_hd__nand3_1
XFILLER_0_89_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16711_ _07119_ _07121_ VGND VGND VPWR VPWR _07122_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_107_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17691_ _07207_ _07649_ _07780_ _06947_ VGND VGND VPWR VPWR _08190_ sky130_fd_sc_hd__a22o_1
X_16642_ _07019_ _07046_ VGND VGND VPWR VPWR _07048_ sky130_fd_sc_hd__xnor2_1
X_13854_ _04013_ _04014_ VGND VGND VPWR VPWR _04015_ sky130_fd_sc_hd__xnor2_1
X_12805_ _00824_ _00853_ _00852_ VGND VGND VPWR VPWR _02898_ sky130_fd_sc_hd__a21oi_1
X_16573_ _06970_ _06972_ _06749_ _06891_ VGND VGND VPWR VPWR _06973_ sky130_fd_sc_hd__o211a_1
X_13785_ _03934_ _03936_ _03937_ VGND VGND VPWR VPWR _03939_ sky130_fd_sc_hd__a21o_1
X_10997_ _06971_ _06689_ _01087_ _01088_ VGND VGND VPWR VPWR _01090_ sky130_fd_sc_hd__a22o_1
XFILLER_0_96_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15524_ _02998_ _05652_ VGND VGND VPWR VPWR _05837_ sky130_fd_sc_hd__nand2_1
X_18312_ _08638_ _08787_ _07604_ _07859_ VGND VGND VPWR VPWR _08866_ sky130_fd_sc_hd__o211a_1
XFILLER_0_32_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12736_ _02797_ _02795_ VGND VGND VPWR VPWR _02829_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_32_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18243_ _08786_ _08790_ VGND VGND VPWR VPWR _08791_ sky130_fd_sc_hd__or2_1
XFILLER_0_154_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15455_ _07515_ _05758_ _05986_ _03008_ VGND VGND VPWR VPWR _05762_ sky130_fd_sc_hd__a22o_1
X_12667_ _02719_ _02725_ VGND VGND VPWR VPWR _02760_ sky130_fd_sc_hd__xnor2_1
X_14406_ _03014_ _02124_ _04615_ _04617_ VGND VGND VPWR VPWR _04618_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_65_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11618_ _01614_ _01616_ _01613_ VGND VGND VPWR VPWR _01711_ sky130_fd_sc_hd__a21o_1
X_18174_ _07109_ _07859_ _08640_ _08639_ VGND VGND VPWR VPWR _08716_ sky130_fd_sc_hd__a31o_1
X_15386_ _05685_ _05686_ VGND VGND VPWR VPWR _05687_ sky130_fd_sc_hd__and2_1
XFILLER_0_5_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12598_ _02683_ _02684_ _02690_ VGND VGND VPWR VPWR _02691_ sky130_fd_sc_hd__or3_1
XFILLER_0_41_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17125_ _00558_ _06437_ _07573_ VGND VGND VPWR VPWR _07574_ sky130_fd_sc_hd__o21a_1
X_14337_ _04540_ _04541_ _04425_ _04382_ VGND VGND VPWR VPWR _04543_ sky130_fd_sc_hd__o211a_1
X_11549_ _01564_ _01604_ _01640_ _01641_ VGND VGND VPWR VPWR _01642_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_52_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17056_ _06764_ _07194_ VGND VGND VPWR VPWR _07498_ sky130_fd_sc_hd__nor2_1
X_14268_ _04463_ _04466_ VGND VGND VPWR VPWR _04467_ sky130_fd_sc_hd__xor2_2
XFILLER_0_122_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16007_ _02476_ _00167_ VGND VGND VPWR VPWR _06357_ sky130_fd_sc_hd__nor2_1
X_13219_ _00125_ VGND VGND VPWR VPWR _03321_ sky130_fd_sc_hd__clkbuf_4
XTAP_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14199_ _04222_ _04225_ VGND VGND VPWR VPWR _04392_ sky130_fd_sc_hd__and2b_1
XTAP_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17958_ _08469_ _08480_ VGND VGND VPWR VPWR _08481_ sky130_fd_sc_hd__xnor2_1
X_16909_ _07336_ _07337_ VGND VGND VPWR VPWR _07338_ sky130_fd_sc_hd__and2_1
X_17889_ _08298_ _08309_ VGND VGND VPWR VPWR _08406_ sky130_fd_sc_hd__or2b_1
XFILLER_0_73_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10920_ _01007_ _01012_ VGND VGND VPWR VPWR _01013_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_79_650 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10851_ ApproximateM_inst.lob_16.lob2.genblk1\[13\].genblk1.mux.sel ApproximateM_inst.lob_16.lob2.genblk1\[12\].genblk1.mux.sel
+ net209 _03388_ VGND VGND VPWR VPWR _00944_ sky130_fd_sc_hd__and4_1
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13570_ _00148_ _00149_ _04154_ _00563_ VGND VGND VPWR VPWR _03704_ sky130_fd_sc_hd__and4_1
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10782_ _00190_ _00192_ _00134_ _00108_ _00874_ VGND VGND VPWR VPWR _00875_ sky130_fd_sc_hd__a41o_1
XFILLER_0_94_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12521_ _02560_ _02562_ _02564_ _02558_ VGND VGND VPWR VPWR _02614_ sky130_fd_sc_hd__o31a_1
XFILLER_0_66_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15240_ _05443_ _05455_ VGND VGND VPWR VPWR _05527_ sky130_fd_sc_hd__and2_1
XPHY_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12452_ _02494_ _02492_ _02493_ VGND VGND VPWR VPWR _02545_ sky130_fd_sc_hd__nand3_1
XFILLER_0_124_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11403_ _01451_ _01444_ _01494_ _01495_ VGND VGND VPWR VPWR _01496_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_152_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15171_ _05444_ _05451_ VGND VGND VPWR VPWR _05452_ sky130_fd_sc_hd__or2_1
XFILLER_0_22_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12383_ _00645_ VGND VGND VPWR VPWR _02476_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_151_257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14122_ _04305_ _04306_ VGND VGND VPWR VPWR _04308_ sky130_fd_sc_hd__xnor2_1
X_11334_ _00195_ _00702_ _00127_ _07559_ _01344_ VGND VGND VPWR VPWR _01427_ sky130_fd_sc_hd__a41o_1
XFILLER_0_22_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14053_ _04230_ _04232_ VGND VGND VPWR VPWR _04233_ sky130_fd_sc_hd__nor2_2
X_18930_ clknet_4_10_0_clk _00084_ VGND VGND VPWR VPWR cla_inst.in2\[16\] sky130_fd_sc_hd__dfxtp_2
X_11265_ _01356_ _01357_ _01110_ VGND VGND VPWR VPWR _01358_ sky130_fd_sc_hd__and3_1
XFILLER_0_120_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13004_ _03093_ _03096_ _03090_ VGND VGND VPWR VPWR _03097_ sky130_fd_sc_hd__mux2_1
X_10216_ _00308_ VGND VGND VPWR VPWR _00309_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_101_880 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18861_ clknet_4_7_0_clk net282 VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__dfxtp_1
X_11196_ _01279_ _01287_ _01286_ VGND VGND VPWR VPWR _01289_ sky130_fd_sc_hd__o21ai_1
X_17812_ _08320_ _08321_ VGND VGND VPWR VPWR _08323_ sky130_fd_sc_hd__nand2_1
X_10147_ _00236_ _00239_ VGND VGND VPWR VPWR _00240_ sky130_fd_sc_hd__xnor2_1
X_18792_ _09298_ _09302_ VGND VGND VPWR VPWR _09304_ sky130_fd_sc_hd__and2_1
XFILLER_0_27_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14955_ _02985_ _02988_ _09311_ _08224_ _05105_ VGND VGND VPWR VPWR _05217_ sky130_fd_sc_hd__a41o_1
X_17743_ _07256_ _08234_ _08236_ _08247_ VGND VGND VPWR VPWR _08248_ sky130_fd_sc_hd__a31o_1
XFILLER_0_89_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10078_ _04242_ VGND VGND VPWR VPWR _00171_ sky130_fd_sc_hd__buf_4
X_13906_ _04068_ _04071_ VGND VGND VPWR VPWR _04072_ sky130_fd_sc_hd__or2_1
X_14886_ _05032_ _05030_ VGND VGND VPWR VPWR _05142_ sky130_fd_sc_hd__and2b_1
X_17674_ _08070_ _08072_ _08069_ VGND VGND VPWR VPWR _08172_ sky130_fd_sc_hd__o21ai_1
X_13837_ _03792_ _03995_ VGND VGND VPWR VPWR _03996_ sky130_fd_sc_hd__xnor2_1
X_16625_ _06653_ _06874_ VGND VGND VPWR VPWR _07029_ sky130_fd_sc_hd__nor2_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16556_ _06812_ _06529_ _06953_ VGND VGND VPWR VPWR _06954_ sky130_fd_sc_hd__or3_1
X_13768_ _03920_ VGND VGND VPWR VPWR _03921_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_84_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_127_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15507_ _00115_ _00339_ _05814_ _05815_ VGND VGND VPWR VPWR _05818_ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12719_ _02789_ _02811_ VGND VGND VPWR VPWR _02812_ sky130_fd_sc_hd__or2b_1
XFILLER_0_72_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16487_ _06812_ _06529_ _06530_ VGND VGND VPWR VPWR _06879_ sky130_fd_sc_hd__or3_1
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_128_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13699_ _03843_ _03844_ VGND VGND VPWR VPWR _03845_ sky130_fd_sc_hd__xor2_1
X_15438_ _05741_ _05742_ VGND VGND VPWR VPWR _05743_ sky130_fd_sc_hd__nor2_1
X_18226_ _08750_ _08756_ _08772_ _06721_ _06776_ VGND VGND VPWR VPWR _09402_ sky130_fd_sc_hd__o32a_2
XFILLER_0_5_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_131_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15369_ _00591_ _05652_ _05667_ VGND VGND VPWR VPWR _05668_ sky130_fd_sc_hd__and3_1
X_18157_ _08662_ _08664_ VGND VGND VPWR VPWR _08697_ sky130_fd_sc_hd__and2b_1
XFILLER_0_142_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17108_ _07443_ _07445_ VGND VGND VPWR VPWR _07555_ sky130_fd_sc_hd__or2_1
X_18088_ _02259_ _07387_ _08621_ VGND VGND VPWR VPWR _08622_ sky130_fd_sc_hd__or3b_1
XFILLER_0_40_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09930_ cla_inst.in1\[21\] VGND VGND VPWR VPWR _08746_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_110_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17039_ _07458_ _07465_ _07479_ VGND VGND VPWR VPWR _07480_ sky130_fd_sc_hd__and3_1
XFILLER_0_1_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09861_ _07973_ cla_inst.in1\[23\] cla_inst.in1\[22\] _07984_ VGND VGND VPWR VPWR
+ _07995_ sky130_fd_sc_hd__a22o_1
XFILLER_0_68_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09792_ ApproximateM_inst.lob_16.lob2.genblk1\[3\].genblk1.mux.sel VGND VGND VPWR
+ VPWR _07243_ sky130_fd_sc_hd__buf_4
XTAP_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_114_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11050_ _01134_ _01135_ _01142_ VGND VGND VPWR VPWR _01143_ sky130_fd_sc_hd__nand3_2
XFILLER_0_101_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10001_ _09027_ _09341_ _09342_ _09343_ VGND VGND VPWR VPWR _09344_ sky130_fd_sc_hd__and4bb_2
X_14740_ _04975_ _04976_ _04981_ VGND VGND VPWR VPWR _04982_ sky130_fd_sc_hd__nand3_2
XFILLER_0_99_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11952_ _01575_ VGND VGND VPWR VPWR _02045_ sky130_fd_sc_hd__clkinv_4
Xwb_buttons_leds_152 VGND VGND VPWR VPWR wb_buttons_leds_152/HI led_enb[1] sky130_fd_sc_hd__conb_1
Xwb_buttons_leds_163 VGND VGND VPWR VPWR wb_buttons_leds_163/HI o_wb_stall sky130_fd_sc_hd__conb_1
X_10903_ _00991_ _00995_ VGND VGND VPWR VPWR _00996_ sky130_fd_sc_hd__xor2_2
X_14671_ _04747_ _04748_ _04746_ VGND VGND VPWR VPWR _04907_ sky130_fd_sc_hd__o21ai_1
X_11883_ _01944_ _01973_ _01974_ _01975_ VGND VGND VPWR VPWR _01976_ sky130_fd_sc_hd__or4_4
X_16410_ _02823_ _06785_ _06795_ VGND VGND VPWR VPWR _06796_ sky130_fd_sc_hd__o21ai_1
X_13622_ _03590_ _03754_ _03758_ net336 VGND VGND VPWR VPWR _03761_ sky130_fd_sc_hd__o211ai_4
X_10834_ cla_inst.in2\[16\] ApproximateM_inst.lob_16.lob2.genblk2.mux_final.sel ApproximateM_inst.lob_16.lob1.genblk1\[7\].genblk1.mux.sel
+ ApproximateM_inst.lob_16.lob1.genblk1\[6\].genblk1.mux.sel VGND VGND VPWR VPWR _00927_
+ sky130_fd_sc_hd__and4_1
X_17390_ _06561_ _07124_ _07516_ _07861_ VGND VGND VPWR VPWR _07862_ sky130_fd_sc_hd__or4_1
XFILLER_0_66_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16341_ _06720_ VGND VGND VPWR VPWR _06721_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_149_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13553_ _00203_ _01962_ VGND VGND VPWR VPWR _03686_ sky130_fd_sc_hd__nand2_1
XFILLER_0_94_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10765_ _00162_ _00230_ VGND VGND VPWR VPWR _00858_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_67_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_137_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12504_ _07352_ _00146_ _02595_ _02596_ VGND VGND VPWR VPWR _02597_ sky130_fd_sc_hd__nand4_2
XFILLER_0_137_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16272_ _03117_ _06630_ _06644_ _06645_ VGND VGND VPWR VPWR _06647_ sky130_fd_sc_hd__a211o_1
XFILLER_0_125_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13484_ _03990_ _06062_ _03385_ _03384_ _00459_ VGND VGND VPWR VPWR _03610_ sky130_fd_sc_hd__a32o_1
X_10696_ _00786_ _00787_ _00788_ VGND VGND VPWR VPWR _00789_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_152_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15223_ _05428_ _05396_ _05509_ VGND VGND VPWR VPWR _05510_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_81_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18011_ _07125_ _07706_ VGND VGND VPWR VPWR _08538_ sky130_fd_sc_hd__nor2_1
XFILLER_0_113_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12435_ _02460_ _02472_ _02527_ VGND VGND VPWR VPWR _02528_ sky130_fd_sc_hd__and3_1
XFILLER_0_22_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15154_ _02985_ _03456_ VGND VGND VPWR VPWR _05434_ sky130_fd_sc_hd__nand2_1
X_12366_ _02389_ _02457_ _02451_ _02456_ VGND VGND VPWR VPWR _02459_ sky130_fd_sc_hd__o211a_1
X_14105_ _04515_ _02188_ _00498_ _08169_ VGND VGND VPWR VPWR _04289_ sky130_fd_sc_hd__nand4_1
XFILLER_0_22_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11317_ _01324_ _01326_ VGND VGND VPWR VPWR _01410_ sky130_fd_sc_hd__and2b_1
X_15085_ _05350_ _05358_ VGND VGND VPWR VPWR _05359_ sky130_fd_sc_hd__xor2_1
XFILLER_0_22_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12297_ _02295_ _02297_ _02298_ VGND VGND VPWR VPWR _02390_ sky130_fd_sc_hd__or3_1
X_14036_ _03997_ _04173_ _04212_ _04213_ VGND VGND VPWR VPWR _04214_ sky130_fd_sc_hd__o211a_1
X_18913_ clknet_4_8_0_clk _00067_ VGND VGND VPWR VPWR cla_inst.in1\[31\] sky130_fd_sc_hd__dfxtp_1
X_11248_ _00203_ _01264_ VGND VGND VPWR VPWR _01341_ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_56 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18844_ clknet_4_0_0_clk net262 VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__dfxtp_1
X_11179_ _01147_ _01148_ _01237_ VGND VGND VPWR VPWR _01272_ sky130_fd_sc_hd__a21oi_1
X_18775_ _09273_ _09289_ VGND VGND VPWR VPWR _09290_ sky130_fd_sc_hd__and2_1
X_15987_ _06332_ _06333_ _06334_ _02677_ VGND VGND VPWR VPWR _06335_ sky130_fd_sc_hd__a31o_1
X_17726_ _02326_ _02467_ _08226_ _08228_ VGND VGND VPWR VPWR _08229_ sky130_fd_sc_hd__a31oi_4
X_14938_ _04946_ VGND VGND VPWR VPWR _05199_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17657_ _08151_ _08152_ VGND VGND VPWR VPWR _08153_ sky130_fd_sc_hd__nand2_1
X_14869_ _05121_ _05122_ VGND VGND VPWR VPWR _05123_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_147_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16608_ _06421_ _06996_ _06997_ _07005_ _07010_ VGND VGND VPWR VPWR _07011_ sky130_fd_sc_hd__a311o_1
X_17588_ _08076_ _08077_ VGND VGND VPWR VPWR _08078_ sky130_fd_sc_hd__or2_1
XFILLER_0_147_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16539_ _06826_ _06899_ VGND VGND VPWR VPWR _06935_ sky130_fd_sc_hd__nor2_1
XFILLER_0_46_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18209_ _08676_ _08677_ _08675_ VGND VGND VPWR VPWR _08754_ sky130_fd_sc_hd__a21o_1
XFILLER_0_5_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_531 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold101 _00029_ VGND VGND VPWR VPWR net264 sky130_fd_sc_hd__dlygate4sd3_1
Xhold112 net91 VGND VGND VPWR VPWR net275 sky130_fd_sc_hd__dlygate4sd3_1
Xhold123 _00018_ VGND VGND VPWR VPWR net286 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold134 net86 VGND VGND VPWR VPWR net297 sky130_fd_sc_hd__dlygate4sd3_1
Xhold145 net103 VGND VGND VPWR VPWR net308 sky130_fd_sc_hd__dlygate4sd3_1
X_09913_ _04646_ _04373_ _05333_ _05039_ VGND VGND VPWR VPWR _08561_ sky130_fd_sc_hd__and4_1
XFILLER_0_0_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09844_ _07799_ _07722_ VGND VGND VPWR VPWR _07810_ sky130_fd_sc_hd__and2_4
XTAP_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09775_ _07047_ VGND VGND VPWR VPWR _07058_ sky130_fd_sc_hd__buf_4
XTAP_2306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_247 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_139_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10550_ _00641_ _00642_ VGND VGND VPWR VPWR _00643_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_9_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_144 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10481_ _00572_ _00573_ VGND VGND VPWR VPWR _00574_ sky130_fd_sc_hd__and2_1
X_12220_ _02126_ _02128_ _02303_ VGND VGND VPWR VPWR _02313_ sky130_fd_sc_hd__or3_1
XFILLER_0_60_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12151_ _05562_ _05584_ net206 _00179_ VGND VGND VPWR VPWR _02244_ sky130_fd_sc_hd__and4_1
X_11102_ _01062_ _01067_ VGND VGND VPWR VPWR _01195_ sky130_fd_sc_hd__xnor2_2
X_12082_ _02173_ _02174_ VGND VGND VPWR VPWR _02175_ sky130_fd_sc_hd__or2b_1
X_11033_ _01096_ _01124_ _01125_ VGND VGND VPWR VPWR _01126_ sky130_fd_sc_hd__nand3_2
X_15910_ _06244_ _06253_ VGND VGND VPWR VPWR _06254_ sky130_fd_sc_hd__nand2_1
X_16890_ _07315_ _07316_ VGND VGND VPWR VPWR _07317_ sky130_fd_sc_hd__nor2_1
X_15841_ _06178_ _06179_ VGND VGND VPWR VPWR _06180_ sky130_fd_sc_hd__or2_2
XFILLER_0_99_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18560_ salida\[2\] _09114_ _09118_ salida\[34\] _09128_ VGND VGND VPWR VPWR _09130_
+ sky130_fd_sc_hd__a221o_1
X_15772_ _06026_ _06028_ _06103_ VGND VGND VPWR VPWR _06106_ sky130_fd_sc_hd__or3_1
X_12984_ _02981_ VGND VGND VPWR VPWR _03077_ sky130_fd_sc_hd__buf_4
X_17511_ _07974_ _07993_ VGND VGND VPWR VPWR _07994_ sky130_fd_sc_hd__xor2_1
X_14723_ _04934_ _04935_ VGND VGND VPWR VPWR _04964_ sky130_fd_sc_hd__and2_1
X_11935_ _01949_ _01957_ VGND VGND VPWR VPWR _02028_ sky130_fd_sc_hd__xnor2_2
X_18491_ _06248_ _06413_ _06412_ _06328_ VGND VGND VPWR VPWR _09058_ sky130_fd_sc_hd__o211a_1
XFILLER_0_59_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14654_ _00195_ _00702_ _06062_ _05257_ VGND VGND VPWR VPWR _04889_ sky130_fd_sc_hd__and4_1
X_17442_ _06736_ _06729_ _06731_ _06726_ _02977_ _02981_ VGND VGND VPWR VPWR _07920_
+ sky130_fd_sc_hd__mux4_1
X_11866_ _01949_ net176 _01958_ VGND VGND VPWR VPWR _01959_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_67_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13605_ _03355_ _03528_ VGND VGND VPWR VPWR _03743_ sky130_fd_sc_hd__or2b_1
XFILLER_0_95_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10817_ net227 net169 _04242_ _00179_ VGND VGND VPWR VPWR _00910_ sky130_fd_sc_hd__nand4_2
XFILLER_0_95_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14585_ _03368_ _04647_ _04645_ _04813_ VGND VGND VPWR VPWR _04814_ sky130_fd_sc_hd__a31oi_2
X_17373_ _06957_ _07194_ _07290_ _06961_ VGND VGND VPWR VPWR _07844_ sky130_fd_sc_hd__o22a_1
X_11797_ _01871_ _01887_ _01888_ _01889_ VGND VGND VPWR VPWR _01890_ sky130_fd_sc_hd__nand4_2
XFILLER_0_138_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13536_ _03426_ _03428_ _03666_ VGND VGND VPWR VPWR _03667_ sky130_fd_sc_hd__o21ba_1
X_16324_ _03152_ _06496_ _06702_ _06626_ VGND VGND VPWR VPWR _06703_ sky130_fd_sc_hd__o211a_1
X_10748_ _08006_ _00837_ _00840_ VGND VGND VPWR VPWR _00841_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_125_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16255_ _06627_ VGND VGND VPWR VPWR _06628_ sky130_fd_sc_hd__inv_2
XFILLER_0_36_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13467_ _03588_ _03589_ _03590_ VGND VGND VPWR VPWR _03591_ sky130_fd_sc_hd__or3_4
XFILLER_0_82_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10679_ ApproximateM_inst.lob_16.lob1.genblk1\[5\].genblk1.mux.sel VGND VGND VPWR
+ VPWR _00772_ sky130_fd_sc_hd__buf_6
XFILLER_0_153_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15206_ _05489_ _05490_ VGND VGND VPWR VPWR _05491_ sky130_fd_sc_hd__xor2_2
XFILLER_0_125_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12418_ _02401_ _02413_ VGND VGND VPWR VPWR _02511_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16186_ _03029_ _06420_ _06543_ _06552_ VGND VGND VPWR VPWR _06553_ sky130_fd_sc_hd__o31a_1
X_13398_ _03469_ _03470_ _03514_ _03515_ VGND VGND VPWR VPWR _03516_ sky130_fd_sc_hd__nand4_4
XFILLER_0_50_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15137_ _05411_ _05415_ VGND VGND VPWR VPWR _05416_ sky130_fd_sc_hd__nand2_2
X_12349_ _02372_ _02374_ _02375_ _02369_ VGND VGND VPWR VPWR _02442_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_49_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15068_ _05331_ _05338_ VGND VGND VPWR VPWR _05340_ sky130_fd_sc_hd__nand2_1
X_14019_ _04029_ _04037_ _04194_ VGND VGND VPWR VPWR _04195_ sky130_fd_sc_hd__a21o_1
X_18827_ net69 _09111_ net67 VGND VGND VPWR VPWR _09330_ sky130_fd_sc_hd__or3b_1
XFILLER_0_65_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09560_ _04668_ _04679_ _04711_ VGND VGND VPWR VPWR _04722_ sky130_fd_sc_hd__or3_1
X_18758_ _09250_ VGND VGND VPWR VPWR _09276_ sky130_fd_sc_hd__buf_4
X_17709_ _08086_ _08096_ _08209_ VGND VGND VPWR VPWR _08210_ sky130_fd_sc_hd__a21bo_1
X_09491_ _03706_ _03946_ _03957_ VGND VGND VPWR VPWR _03968_ sky130_fd_sc_hd__nand3_2
X_18689_ net44 _09189_ _09223_ VGND VGND VPWR VPWR _00054_ sky130_fd_sc_hd__o21a_1
XFILLER_0_77_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_144 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_112_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09827_ _07515_ _07537_ _07570_ _07613_ VGND VGND VPWR VPWR _07624_ sky130_fd_sc_hd__and4_1
X_09758_ _06819_ _06830_ _06852_ VGND VGND VPWR VPWR _06873_ sky130_fd_sc_hd__nand3_2
XTAP_2103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09689_ _05997_ _06116_ VGND VGND VPWR VPWR _06127_ sky130_fd_sc_hd__xnor2_4
XTAP_2136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11720_ _03848_ _01151_ _09179_ _07581_ VGND VGND VPWR VPWR _01813_ sky130_fd_sc_hd__and4_1
XTAP_2169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11651_ _01743_ VGND VGND VPWR VPWR _01744_ sky130_fd_sc_hd__inv_2
XTAP_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10602_ _00661_ net165 _00692_ _00693_ VGND VGND VPWR VPWR _00695_ sky130_fd_sc_hd__a2bb2oi_2
XFILLER_0_76_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14370_ _04001_ _07733_ _04575_ _04576_ VGND VGND VPWR VPWR _04578_ sky130_fd_sc_hd__o2bb2a_1
X_11582_ _07853_ _06482_ _01674_ VGND VGND VPWR VPWR _01675_ sky130_fd_sc_hd__and3_2
XFILLER_0_153_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13321_ _03408_ _03409_ _03429_ _03430_ VGND VGND VPWR VPWR _03431_ sky130_fd_sc_hd__a22o_1
XFILLER_0_52_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10533_ _04558_ _05964_ _00624_ _00625_ VGND VGND VPWR VPWR _00626_ sky130_fd_sc_hd__nand4_2
XFILLER_0_51_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16040_ _06391_ _06392_ _04630_ VGND VGND VPWR VPWR _06393_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_135_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13252_ _03353_ _03354_ VGND VGND VPWR VPWR _03357_ sky130_fd_sc_hd__nand2_1
X_10464_ _04012_ VGND VGND VPWR VPWR _00557_ sky130_fd_sc_hd__buf_6
XFILLER_0_122_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12203_ _02277_ _02279_ VGND VGND VPWR VPWR _02296_ sky130_fd_sc_hd__nor2_1
XFILLER_0_33_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13183_ _07091_ _00509_ VGND VGND VPWR VPWR _03283_ sky130_fd_sc_hd__nand2_1
XFILLER_0_60_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10395_ _00465_ _00466_ _00291_ _00431_ VGND VGND VPWR VPWR _00488_ sky130_fd_sc_hd__a211o_4
X_12134_ _02193_ _02226_ VGND VGND VPWR VPWR _02227_ sky130_fd_sc_hd__nand2_1
X_17991_ _04630_ _06391_ _06392_ VGND VGND VPWR VPWR _08517_ sky130_fd_sc_hd__and3_1
XFILLER_0_20_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16942_ _06680_ _07367_ _07369_ _07373_ VGND VGND VPWR VPWR _07375_ sky130_fd_sc_hd__or4_1
X_12065_ _02154_ _02156_ _02157_ VGND VGND VPWR VPWR _02158_ sky130_fd_sc_hd__nor3_1
X_11016_ _07788_ _05975_ _01108_ VGND VGND VPWR VPWR _01109_ sky130_fd_sc_hd__and3_2
X_16873_ _07200_ _07296_ VGND VGND VPWR VPWR _07299_ sky130_fd_sc_hd__nand2_1
X_18612_ salida\[23\] _09159_ _09160_ salida\[55\] _09163_ VGND VGND VPWR VPWR _09167_
+ sky130_fd_sc_hd__a221o_1
X_15824_ _06115_ _06113_ VGND VGND VPWR VPWR _06162_ sky130_fd_sc_hd__and2b_1
XFILLER_0_35_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18543_ _09113_ VGND VGND VPWR VPWR _09114_ sky130_fd_sc_hd__buf_2
X_15755_ _06034_ _06058_ _06059_ VGND VGND VPWR VPWR _06087_ sky130_fd_sc_hd__nand3_1
X_12967_ _02489_ VGND VGND VPWR VPWR _03060_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_59_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14706_ _04942_ _04945_ VGND VGND VPWR VPWR _04946_ sky130_fd_sc_hd__xor2_2
X_11918_ _01922_ _02010_ VGND VGND VPWR VPWR _02011_ sky130_fd_sc_hd__xnor2_1
X_18474_ _03108_ _03760_ _08047_ _09039_ VGND VGND VPWR VPWR _09040_ sky130_fd_sc_hd__o31a_1
X_12898_ _00148_ VGND VGND VPWR VPWR _02991_ sky130_fd_sc_hd__clkbuf_4
X_15686_ _05938_ _05941_ _06012_ VGND VGND VPWR VPWR _06013_ sky130_fd_sc_hd__and3_1
XFILLER_0_75_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17425_ _07821_ _07786_ _07899_ VGND VGND VPWR VPWR _07901_ sky130_fd_sc_hd__or3b_2
XFILLER_0_27_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14637_ _03008_ _07515_ _01962_ _02124_ VGND VGND VPWR VPWR _04870_ sky130_fd_sc_hd__and4_1
XFILLER_0_74_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11849_ _01841_ _01882_ _01883_ _01881_ VGND VGND VPWR VPWR _01942_ sky130_fd_sc_hd__a22o_1
XTAP_1980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14568_ _04776_ _04664_ _04793_ VGND VGND VPWR VPWR _04795_ sky130_fd_sc_hd__and3_1
XFILLER_0_71_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17356_ _04034_ _06889_ VGND VGND VPWR VPWR _07825_ sky130_fd_sc_hd__and2_1
XFILLER_0_144_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16307_ _06332_ _06545_ _06681_ _01503_ _06683_ VGND VGND VPWR VPWR _06684_ sky130_fd_sc_hd__a221o_1
XFILLER_0_27_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13519_ _03622_ _03623_ _03646_ VGND VGND VPWR VPWR _03648_ sky130_fd_sc_hd__and3_1
X_14499_ _04712_ _04713_ _04718_ VGND VGND VPWR VPWR _04719_ sky130_fd_sc_hd__nand3_1
X_17287_ _07302_ _07303_ _07130_ _07126_ VGND VGND VPWR VPWR _07750_ sky130_fd_sc_hd__or4_1
XFILLER_0_153_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16238_ _09263_ _03074_ VGND VGND VPWR VPWR _06609_ sky130_fd_sc_hd__or2_1
XFILLER_0_23_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16169_ _03184_ VGND VGND VPWR VPWR _06534_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09612_ ApproximateM_inst.lob_16.lob2.genblk1\[9\].genblk1.mux.sel VGND VGND VPWR
+ VPWR _05290_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_78_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09543_ _04406_ _04526_ VGND VGND VPWR VPWR _04537_ sky130_fd_sc_hd__or2_4
XFILLER_0_92_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09474_ _03771_ VGND VGND VPWR VPWR _03782_ sky130_fd_sc_hd__buf_4
XFILLER_0_116_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire119 _03888_ VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__buf_1
XFILLER_0_46_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_116_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10180_ _09348_ _00270_ _00271_ _00272_ VGND VGND VPWR VPWR _00273_ sky130_fd_sc_hd__nand4_4
X_13870_ cla_inst.in2\[27\] cla_inst.in2\[26\] _03903_ _03914_ VGND VGND VPWR VPWR
+ _04032_ sky130_fd_sc_hd__and4_2
XFILLER_0_88_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12821_ _02911_ _02912_ _01492_ _01494_ VGND VGND VPWR VPWR _02914_ sky130_fd_sc_hd__a211o_2
X_15540_ _05851_ _05853_ VGND VGND VPWR VPWR _05854_ sky130_fd_sc_hd__or2_1
XTAP_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12752_ _02528_ _02587_ _02471_ VGND VGND VPWR VPWR _02845_ sky130_fd_sc_hd__o21ai_1
XTAP_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11703_ _01764_ _01792_ _01794_ VGND VGND VPWR VPWR _01796_ sky130_fd_sc_hd__or3_1
X_15471_ _05776_ _05777_ _05674_ VGND VGND VPWR VPWR _05779_ sky130_fd_sc_hd__o21a_1
XTAP_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12683_ _02744_ _02752_ _02775_ VGND VGND VPWR VPWR _02776_ sky130_fd_sc_hd__and3_1
XTAP_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14422_ _00253_ _00460_ VGND VGND VPWR VPWR _04636_ sky130_fd_sc_hd__nand2_1
XTAP_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17210_ _06750_ _07665_ _07543_ _07541_ VGND VGND VPWR VPWR _07666_ sky130_fd_sc_hd__a31oi_2
X_11634_ _01221_ _01693_ VGND VGND VPWR VPWR _01727_ sky130_fd_sc_hd__and2_1
XFILLER_0_154_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18190_ _08731_ _08732_ VGND VGND VPWR VPWR _08733_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_126_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14353_ _03138_ _03147_ _03185_ _03190_ _03062_ _02979_ VGND VGND VPWR VPWR _04560_
+ sky130_fd_sc_hd__mux4_1
X_17141_ _06937_ _07314_ VGND VGND VPWR VPWR _07590_ sky130_fd_sc_hd__nor2_1
X_11565_ _06982_ _01005_ _01656_ _01657_ VGND VGND VPWR VPWR _01658_ sky130_fd_sc_hd__a31o_1
XFILLER_0_25_648 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13304_ _06051_ _09303_ _07733_ _06040_ VGND VGND VPWR VPWR _03413_ sky130_fd_sc_hd__a22o_1
XFILLER_0_80_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10516_ _00433_ _00434_ _00432_ VGND VGND VPWR VPWR _00609_ sky130_fd_sc_hd__a21bo_1
X_17072_ _07410_ VGND VGND VPWR VPWR _07516_ sky130_fd_sc_hd__clkbuf_4
X_14284_ _04309_ _04473_ _04483_ VGND VGND VPWR VPWR _04485_ sky130_fd_sc_hd__or3_1
XFILLER_0_24_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11496_ _01587_ _01588_ VGND VGND VPWR VPWR _01589_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_122_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_134_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_664 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13235_ _03335_ _03336_ _00690_ _00692_ VGND VGND VPWR VPWR _03338_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_21_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16023_ _06374_ _03107_ VGND VGND VPWR VPWR _06375_ sky130_fd_sc_hd__or2_1
X_10447_ _00383_ _00394_ VGND VGND VPWR VPWR _00540_ sky130_fd_sc_hd__and2_1
XFILLER_0_110_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_122_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13166_ _00634_ _00660_ _03263_ _03264_ VGND VGND VPWR VPWR _03265_ sky130_fd_sc_hd__a211oi_2
X_10378_ _05508_ _05464_ _00308_ _05964_ VGND VGND VPWR VPWR _00471_ sky130_fd_sc_hd__nand4_1
X_12117_ _02181_ _02204_ _02209_ VGND VGND VPWR VPWR _02210_ sky130_fd_sc_hd__or3_1
X_17974_ _08497_ _08498_ VGND VGND VPWR VPWR _08499_ sky130_fd_sc_hd__and2_1
X_13097_ _03187_ _03189_ _03047_ VGND VGND VPWR VPWR _03190_ sky130_fd_sc_hd__mux2_1
X_12048_ _01905_ _02060_ VGND VGND VPWR VPWR _02141_ sky130_fd_sc_hd__nand2_1
X_16925_ _07289_ _07355_ _00248_ VGND VGND VPWR VPWR _07356_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_46_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16856_ _02776_ _02834_ _07280_ VGND VGND VPWR VPWR _07281_ sky130_fd_sc_hd__o21a_1
XFILLER_0_88_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15807_ _03034_ _06143_ _04247_ VGND VGND VPWR VPWR _06144_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16787_ _07203_ _07204_ VGND VGND VPWR VPWR _07205_ sky130_fd_sc_hd__nor2_1
X_13999_ _03985_ _03999_ VGND VGND VPWR VPWR _04173_ sky130_fd_sc_hd__and2_1
XFILLER_0_62_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18526_ _09074_ _09081_ _09095_ _06721_ _00516_ VGND VGND VPWR VPWR _09410_ sky130_fd_sc_hd__o32a_1
XFILLER_0_153_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15738_ _05994_ _06067_ VGND VGND VPWR VPWR _06069_ sky130_fd_sc_hd__and2_1
XFILLER_0_47_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18457_ _09020_ _09021_ VGND VGND VPWR VPWR _09022_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_118_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15669_ _05920_ _05993_ VGND VGND VPWR VPWR _05994_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_145_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17408_ _07731_ _07767_ _07880_ VGND VGND VPWR VPWR _07882_ sky130_fd_sc_hd__or3_1
XFILLER_0_44_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18388_ _03760_ _08047_ VGND VGND VPWR VPWR _08947_ sky130_fd_sc_hd__nor2_1
XFILLER_0_90_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17339_ _04853_ _06371_ _06370_ VGND VGND VPWR VPWR _07807_ sky130_fd_sc_hd__a21o_1
XFILLER_0_70_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_114_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19009_ clknet_4_1_0_clk _09376_ VGND VGND VPWR VPWR salida\[62\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_141_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_140_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09526_ _04340_ VGND VGND VPWR VPWR _04351_ sky130_fd_sc_hd__buf_6
XFILLER_0_39_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_148_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09457_ _03366_ VGND VGND VPWR VPWR _03596_ sky130_fd_sc_hd__buf_4
XFILLER_0_137_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_559 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_149_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_710 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11350_ _01440_ _01441_ _01337_ _01377_ VGND VGND VPWR VPWR _01443_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_132_620 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10301_ _00384_ _00393_ VGND VGND VPWR VPWR _00394_ sky130_fd_sc_hd__xnor2_1
X_11281_ _01371_ _01372_ _01370_ _01373_ VGND VGND VPWR VPWR _01374_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_105_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_120_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13020_ _03023_ _03112_ VGND VGND VPWR VPWR _03113_ sky130_fd_sc_hd__nand2_1
X_10232_ _00316_ _00324_ VGND VGND VPWR VPWR _00325_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_30_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10163_ _00175_ _03618_ _00218_ _00173_ VGND VGND VPWR VPWR _00256_ sky130_fd_sc_hd__a22o_1
XFILLER_0_100_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14971_ _00362_ _05856_ VGND VGND VPWR VPWR _05234_ sky130_fd_sc_hd__nand2_1
X_10094_ _00170_ _00172_ _00182_ _00185_ VGND VGND VPWR VPWR _00187_ sky130_fd_sc_hd__a22oi_1
X_16710_ _07022_ _07027_ _07120_ VGND VGND VPWR VPWR _07121_ sky130_fd_sc_hd__a21oi_1
X_13922_ _04018_ _04020_ VGND VGND VPWR VPWR _04089_ sky130_fd_sc_hd__or2b_1
X_17690_ _07302_ _07303_ _07516_ _07511_ VGND VGND VPWR VPWR _08189_ sky130_fd_sc_hd__or4_1
XFILLER_0_88_117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16641_ _07021_ _07045_ VGND VGND VPWR VPWR _07046_ sky130_fd_sc_hd__xnor2_1
X_13853_ _03839_ _03842_ _03840_ VGND VGND VPWR VPWR _04014_ sky130_fd_sc_hd__o21ba_2
XFILLER_0_88_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12804_ _01486_ _01487_ VGND VGND VPWR VPWR _02897_ sky130_fd_sc_hd__nand2_1
XFILLER_0_85_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16572_ _06882_ _06883_ VGND VGND VPWR VPWR _06972_ sky130_fd_sc_hd__and2b_1
X_13784_ _03934_ _03936_ _03937_ VGND VGND VPWR VPWR _03938_ sky130_fd_sc_hd__nand3_1
X_10996_ _06971_ _06689_ _01087_ _01088_ VGND VGND VPWR VPWR _01089_ sky130_fd_sc_hd__and4_1
XFILLER_0_69_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18311_ _08862_ _08863_ VGND VGND VPWR VPWR _08864_ sky130_fd_sc_hd__nor2_1
XTAP_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15523_ _05832_ _05835_ VGND VGND VPWR VPWR _05836_ sky130_fd_sc_hd__nand2_1
XTAP_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_96_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12735_ _02826_ _02827_ VGND VGND VPWR VPWR _02828_ sky130_fd_sc_hd__and2_1
XFILLER_0_139_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18242_ _08787_ _08788_ VGND VGND VPWR VPWR _08790_ sky130_fd_sc_hd__xor2_1
X_15454_ _03008_ _07515_ _05758_ _05986_ VGND VGND VPWR VPWR _05761_ sky130_fd_sc_hd__and4_1
XFILLER_0_44_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12666_ _02754_ _02756_ _02757_ _02758_ VGND VGND VPWR VPWR _02759_ sky130_fd_sc_hd__or4_2
XFILLER_0_127_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_795 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14405_ _04614_ VGND VGND VPWR VPWR _04617_ sky130_fd_sc_hd__inv_2
X_11617_ _01610_ _01619_ _01708_ _01709_ VGND VGND VPWR VPWR _01710_ sky130_fd_sc_hd__o211ai_2
X_18173_ _08712_ _08714_ VGND VGND VPWR VPWR _08715_ sky130_fd_sc_hd__or2_1
X_15385_ _05677_ _05684_ VGND VGND VPWR VPWR _05686_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12597_ _02687_ _02688_ _02689_ VGND VGND VPWR VPWR _02690_ sky130_fd_sc_hd__or3_1
XFILLER_0_154_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17124_ _06424_ _06438_ VGND VGND VPWR VPWR _07573_ sky130_fd_sc_hd__nor2_1
X_14336_ _04425_ _04382_ _04540_ _04541_ VGND VGND VPWR VPWR _04542_ sky130_fd_sc_hd__a211oi_2
X_11548_ _01621_ _01639_ _01638_ VGND VGND VPWR VPWR _01641_ sky130_fd_sc_hd__o21a_1
XFILLER_0_107_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14267_ _04464_ _04465_ VGND VGND VPWR VPWR _04466_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_122_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17055_ _06657_ _07396_ VGND VGND VPWR VPWR _07497_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11479_ _08724_ _04067_ _01570_ _01571_ VGND VGND VPWR VPWR _01572_ sky130_fd_sc_hd__a31o_1
XFILLER_0_122_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13218_ _00681_ _00682_ VGND VGND VPWR VPWR _03320_ sky130_fd_sc_hd__nor2_1
X_16006_ _06354_ _06355_ _01829_ VGND VGND VPWR VPWR _06356_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_21_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14198_ _04387_ _04388_ _04389_ VGND VGND VPWR VPWR _04391_ sky130_fd_sc_hd__o21a_1
XTAP_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_567 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13149_ _03245_ _03246_ VGND VGND VPWR VPWR _03247_ sky130_fd_sc_hd__xor2_2
XTAP_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17957_ _08470_ _08479_ VGND VGND VPWR VPWR _08480_ sky130_fd_sc_hd__xnor2_1
X_16908_ _06665_ _07332_ _07335_ VGND VGND VPWR VPWR _07337_ sky130_fd_sc_hd__o21ai_1
X_17888_ _08403_ _08404_ VGND VGND VPWR VPWR _08405_ sky130_fd_sc_hd__or2_1
X_16839_ _07259_ _07260_ VGND VGND VPWR VPWR _07262_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18509_ _00516_ _09076_ _06512_ VGND VGND VPWR VPWR _09077_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_145_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10850_ ApproximateM_inst.lob_16.lob2.genblk1\[11\].genblk1.mux.sel _03903_ VGND
+ VGND VPWR VPWR _00943_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09509_ _04099_ _04132_ _04143_ _04154_ VGND VGND VPWR VPWR _04165_ sky130_fd_sc_hd__and4_1
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10781_ _00169_ _00180_ _00872_ _00873_ VGND VGND VPWR VPWR _00874_ sky130_fd_sc_hd__and4_1
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12520_ _02605_ _02606_ _02612_ VGND VGND VPWR VPWR _02613_ sky130_fd_sc_hd__or3_4
XFILLER_0_149_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12451_ _02498_ _02543_ VGND VGND VPWR VPWR _02544_ sky130_fd_sc_hd__nand2_1
XFILLER_0_136_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_220 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_152_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11402_ _01492_ _01493_ _01452_ _01453_ VGND VGND VPWR VPWR _01495_ sky130_fd_sc_hd__o211a_1
XFILLER_0_151_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15170_ _05448_ _05450_ VGND VGND VPWR VPWR _05451_ sky130_fd_sc_hd__or2_1
XFILLER_0_117_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12382_ _02425_ _02474_ VGND VGND VPWR VPWR _02475_ sky130_fd_sc_hd__nor2_1
XFILLER_0_151_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_90 _08880_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14121_ _02533_ _03456_ _04134_ _04133_ VGND VGND VPWR VPWR _04306_ sky130_fd_sc_hd__a31o_1
XFILLER_0_105_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_151_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11333_ _00874_ _01425_ VGND VGND VPWR VPWR _01426_ sky130_fd_sc_hd__or2_1
XFILLER_0_104_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_120_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_163 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14052_ _04228_ _04229_ _04089_ _04090_ VGND VGND VPWR VPWR _04232_ sky130_fd_sc_hd__o211a_1
X_11264_ _09354_ VGND VGND VPWR VPWR _01357_ sky130_fd_sc_hd__buf_4
X_13003_ _03040_ _03095_ VGND VGND VPWR VPWR _03096_ sky130_fd_sc_hd__nand2_1
X_10215_ _05693_ VGND VGND VPWR VPWR _00308_ sky130_fd_sc_hd__buf_4
XFILLER_0_120_678 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18860_ clknet_4_7_0_clk net284 VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__dfxtp_1
X_11195_ _01279_ _01286_ _01287_ VGND VGND VPWR VPWR _01288_ sky130_fd_sc_hd__or3_1
XFILLER_0_101_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17811_ _08318_ _08319_ VGND VGND VPWR VPWR _08321_ sky130_fd_sc_hd__or2_1
X_10146_ _00237_ _00238_ VGND VGND VPWR VPWR _00239_ sky130_fd_sc_hd__and2b_1
X_18791_ _03368_ net47 _09301_ VGND VGND VPWR VPWR _09302_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17742_ _06421_ _08237_ _08238_ _08240_ _08245_ VGND VGND VPWR VPWR _08247_ sky130_fd_sc_hd__a311o_1
X_14954_ _05214_ _05215_ VGND VGND VPWR VPWR _05216_ sky130_fd_sc_hd__xnor2_1
X_10077_ _00169_ VGND VGND VPWR VPWR _00170_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_27_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13905_ _03741_ _03746_ _03902_ _04070_ VGND VGND VPWR VPWR _04071_ sky130_fd_sc_hd__o31a_1
X_17673_ _08167_ _08170_ VGND VGND VPWR VPWR _08171_ sky130_fd_sc_hd__xor2_1
X_14885_ _04877_ _05029_ VGND VGND VPWR VPWR _05141_ sky130_fd_sc_hd__and2b_1
X_16624_ _07022_ _07027_ VGND VGND VPWR VPWR _07028_ sky130_fd_sc_hd__xnor2_1
X_13836_ _03993_ _03994_ VGND VGND VPWR VPWR _03995_ sky130_fd_sc_hd__and2_1
XFILLER_0_58_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16555_ _03804_ _03826_ _03399_ VGND VGND VPWR VPWR _06953_ sky130_fd_sc_hd__or3_1
XFILLER_0_128_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10979_ _01069_ _01070_ _01071_ VGND VGND VPWR VPWR _01072_ sky130_fd_sc_hd__a21o_1
X_13767_ _02972_ VGND VGND VPWR VPWR _03920_ sky130_fd_sc_hd__clkbuf_4
X_15506_ _05816_ VGND VGND VPWR VPWR _05817_ sky130_fd_sc_hd__inv_2
X_12718_ _02786_ _02787_ _02788_ _02782_ VGND VGND VPWR VPWR _02811_ sky130_fd_sc_hd__a31o_1
XFILLER_0_127_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16486_ _03184_ _06529_ net150 _03313_ VGND VGND VPWR VPWR _06878_ sky130_fd_sc_hd__a211o_1
XFILLER_0_45_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13698_ _00253_ _01575_ _03680_ _03679_ VGND VGND VPWR VPWR _03844_ sky130_fd_sc_hd__a31o_1
XFILLER_0_72_326 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18225_ _06426_ _06447_ _08758_ _08771_ VGND VGND VPWR VPWR _08772_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_143_704 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15437_ _02993_ _02996_ _00495_ _00339_ VGND VGND VPWR VPWR _05742_ sky130_fd_sc_hd__and4_1
XFILLER_0_84_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12649_ _02733_ _02739_ _02740_ _02741_ VGND VGND VPWR VPWR _02742_ sky130_fd_sc_hd__a211o_1
XFILLER_0_115_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_871 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18156_ _08695_ VGND VGND VPWR VPWR _08696_ sky130_fd_sc_hd__inv_2
X_15368_ _05665_ _05666_ VGND VGND VPWR VPWR _05667_ sky130_fd_sc_hd__nor2_1
XFILLER_0_25_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17107_ _07552_ _07553_ VGND VGND VPWR VPWR _07554_ sky130_fd_sc_hd__xnor2_1
X_14319_ _04514_ _04522_ VGND VGND VPWR VPWR _04523_ sky130_fd_sc_hd__xnor2_1
X_18087_ _08619_ _08620_ VGND VGND VPWR VPWR _08621_ sky130_fd_sc_hd__and2_1
X_15299_ _05590_ _05591_ VGND VGND VPWR VPWR _05592_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_1_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17038_ _03921_ _03120_ _04826_ _07468_ _07478_ VGND VGND VPWR VPWR _07479_ sky130_fd_sc_hd__o311a_1
XFILLER_0_1_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09860_ ApproximateM_inst.lob_16.lob2.genblk1\[4\].genblk1.mux.sel VGND VGND VPWR
+ VPWR _07984_ sky130_fd_sc_hd__buf_6
XTAP_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09791_ _07221_ VGND VGND VPWR VPWR _07232_ sky130_fd_sc_hd__buf_4
XTAP_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18989_ clknet_4_6_0_clk _09385_ VGND VGND VPWR VPWR salida\[42\] sky130_fd_sc_hd__dfxtp_1
XTAP_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10000_ _09005_ _09016_ net166 _06906_ VGND VGND VPWR VPWR _09343_ sky130_fd_sc_hd__a211o_1
X_09989_ cla_inst.in1\[29\] VGND VGND VPWR VPWR _09303_ sky130_fd_sc_hd__clkbuf_4
X_11951_ _04700_ VGND VGND VPWR VPWR _02044_ sky130_fd_sc_hd__clkinv_4
Xwb_buttons_leds_153 VGND VGND VPWR VPWR wb_buttons_leds_153/HI led_enb[2] sky130_fd_sc_hd__conb_1
X_10902_ _05497_ _00993_ _00994_ VGND VGND VPWR VPWR _00995_ sky130_fd_sc_hd__a21bo_1
X_14670_ _00115_ _05888_ _04784_ _04783_ VGND VGND VPWR VPWR _04906_ sky130_fd_sc_hd__a31o_1
X_11882_ _01943_ _01919_ _01941_ VGND VGND VPWR VPWR _01975_ sky130_fd_sc_hd__and3_1
X_13621_ _03755_ _03756_ _03757_ VGND VGND VPWR VPWR _03759_ sky130_fd_sc_hd__a21o_1
X_10833_ _00918_ _00919_ _00924_ VGND VGND VPWR VPWR _00926_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_66_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16340_ _02966_ _06459_ VGND VGND VPWR VPWR _06720_ sky130_fd_sc_hd__or2_2
X_10764_ _00828_ _00851_ _00827_ VGND VGND VPWR VPWR _00857_ sky130_fd_sc_hd__a21bo_2
X_13552_ _03682_ _03683_ VGND VGND VPWR VPWR _03685_ sky130_fd_sc_hd__xor2_1
XFILLER_0_66_164 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_109_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12503_ _07973_ _00196_ _01031_ _07221_ VGND VGND VPWR VPWR _02596_ sky130_fd_sc_hd__a22o_1
X_13483_ _03398_ _03400_ VGND VGND VPWR VPWR _03609_ sky130_fd_sc_hd__nand2_1
X_16271_ _03036_ _02965_ _06422_ VGND VGND VPWR VPWR _06645_ sky130_fd_sc_hd__or3_4
X_10695_ _04427_ _03739_ _03804_ _04635_ VGND VGND VPWR VPWR _00788_ sky130_fd_sc_hd__a22o_1
XFILLER_0_109_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18010_ _08535_ _08536_ VGND VGND VPWR VPWR _08537_ sky130_fd_sc_hd__xnor2_1
X_15222_ _05506_ _05507_ VGND VGND VPWR VPWR _05509_ sky130_fd_sc_hd__nand2_1
X_12434_ _02523_ _02526_ VGND VGND VPWR VPWR _02527_ sky130_fd_sc_hd__or2_1
XFILLER_0_35_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15153_ _02987_ _00665_ _05317_ VGND VGND VPWR VPWR _05433_ sky130_fd_sc_hd__and3_1
X_12365_ _02451_ _02456_ _02389_ _02457_ VGND VGND VPWR VPWR _02458_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_50_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_105_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14104_ _04438_ _07722_ _08169_ _04515_ VGND VGND VPWR VPWR _04288_ sky130_fd_sc_hd__a22o_1
X_11316_ _01407_ _01408_ VGND VGND VPWR VPWR _01409_ sky130_fd_sc_hd__nor2_1
XFILLER_0_132_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15084_ _05351_ _05357_ VGND VGND VPWR VPWR _05358_ sky130_fd_sc_hd__xor2_1
XFILLER_0_50_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12296_ _02385_ _02387_ _02388_ VGND VGND VPWR VPWR _02389_ sky130_fd_sc_hd__nor3_1
X_14035_ _04210_ _04211_ _04191_ VGND VGND VPWR VPWR _04213_ sky130_fd_sc_hd__o21ai_1
X_18912_ clknet_4_8_0_clk _00066_ VGND VGND VPWR VPWR cla_inst.in1\[30\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_38_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11247_ _00204_ _01248_ _01259_ VGND VGND VPWR VPWR _01340_ sky130_fd_sc_hd__and3_1
XFILLER_0_120_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18843_ clknet_4_0_0_clk net253 VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11178_ _01251_ _01270_ VGND VGND VPWR VPWR _01271_ sky130_fd_sc_hd__xnor2_1
X_10129_ _00220_ _00221_ VGND VGND VPWR VPWR _00222_ sky130_fd_sc_hd__or2_1
X_18774_ _06374_ net41 _09276_ VGND VGND VPWR VPWR _09289_ sky130_fd_sc_hd__mux2_1
X_15986_ _07711_ _00357_ _07657_ _02505_ VGND VGND VPWR VPWR _06334_ sky130_fd_sc_hd__a22o_1
XFILLER_0_54_12 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17725_ _03930_ _08227_ VGND VGND VPWR VPWR _08228_ sky130_fd_sc_hd__nand2_1
X_14937_ _05196_ _05197_ VGND VGND VPWR VPWR _05198_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17656_ _02044_ _06755_ _06764_ _07933_ VGND VGND VPWR VPWR _08152_ sky130_fd_sc_hd__or4_1
X_14868_ _04992_ _04998_ VGND VGND VPWR VPWR _05122_ sky130_fd_sc_hd__and2_1
X_16607_ _06543_ _06434_ _07006_ _07009_ VGND VGND VPWR VPWR _07010_ sky130_fd_sc_hd__a31o_1
X_13819_ _03974_ _03975_ VGND VGND VPWR VPWR _03976_ sky130_fd_sc_hd__xor2_2
X_17587_ _08074_ _08075_ _08066_ VGND VGND VPWR VPWR _08077_ sky130_fd_sc_hd__o21a_1
X_14799_ _05045_ _05046_ VGND VGND VPWR VPWR _05047_ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16538_ _06898_ _06897_ VGND VGND VPWR VPWR _06934_ sky130_fd_sc_hd__and2b_1
XFILLER_0_128_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_624 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16469_ _03120_ _03565_ _06850_ _06859_ VGND VGND VPWR VPWR _06860_ sky130_fd_sc_hd__o211a_1
XFILLER_0_73_679 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18208_ _08751_ _08752_ VGND VGND VPWR VPWR _08753_ sky130_fd_sc_hd__and2b_1
XFILLER_0_26_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18139_ _08675_ _08676_ _08677_ VGND VGND VPWR VPWR _08678_ sky130_fd_sc_hd__and3b_1
XFILLER_0_130_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_124_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold102 net93 VGND VGND VPWR VPWR net265 sky130_fd_sc_hd__dlygate4sd3_1
Xhold113 _00021_ VGND VGND VPWR VPWR net276 sky130_fd_sc_hd__dlygate4sd3_1
Xhold124 net99 VGND VGND VPWR VPWR net287 sky130_fd_sc_hd__dlygate4sd3_1
Xhold135 _00016_ VGND VGND VPWR VPWR net298 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold146 _00032_ VGND VGND VPWR VPWR net309 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09912_ _04558_ _05486_ VGND VGND VPWR VPWR _08550_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09843_ ApproximateM_inst.lob_16.lob2.mux.sel VGND VGND VPWR VPWR _07799_ sky130_fd_sc_hd__clkbuf_4
XTAP_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09774_ _07036_ VGND VGND VPWR VPWR _07047_ sky130_fd_sc_hd__clkbuf_8
XTAP_2307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_80 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10480_ _00571_ _00560_ _00561_ VGND VGND VPWR VPWR _00573_ sky130_fd_sc_hd__or3_1
XFILLER_0_44_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12150_ _06993_ _00166_ _02241_ _02242_ VGND VGND VPWR VPWR _02243_ sky130_fd_sc_hd__a31o_1
X_11101_ _01175_ _01171_ VGND VGND VPWR VPWR _01194_ sky130_fd_sc_hd__or2b_1
X_12081_ _02169_ _02081_ VGND VGND VPWR VPWR _02174_ sky130_fd_sc_hd__xor2_1
XFILLER_0_5_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11032_ _06971_ _05246_ _01094_ _01095_ VGND VGND VPWR VPWR _01125_ sky130_fd_sc_hd__a22o_1
X_15840_ _06121_ _06124_ _06177_ VGND VGND VPWR VPWR _06179_ sky130_fd_sc_hd__and3_1
X_15771_ _06026_ _06028_ _06103_ VGND VGND VPWR VPWR _06104_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_99_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12983_ _03070_ _03075_ _03050_ VGND VGND VPWR VPWR _03076_ sky130_fd_sc_hd__mux2_1
X_17510_ _07991_ _07992_ VGND VGND VPWR VPWR _07993_ sky130_fd_sc_hd__and2b_1
X_14722_ _00592_ _04900_ _04899_ VGND VGND VPWR VPWR _04963_ sky130_fd_sc_hd__and3_1
X_18490_ _06836_ _09055_ _09056_ VGND VGND VPWR VPWR _09057_ sky130_fd_sc_hd__or3_1
X_11934_ _02009_ _02024_ _02026_ VGND VGND VPWR VPWR _02027_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_59_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17441_ _06375_ _06545_ _07917_ _03108_ VGND VGND VPWR VPWR _07918_ sky130_fd_sc_hd__a22o_1
X_14653_ _00191_ _06094_ _00460_ _00189_ VGND VGND VPWR VPWR _04888_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_39_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11865_ _01953_ _01956_ VGND VGND VPWR VPWR _01958_ sky130_fd_sc_hd__and2_1
XFILLER_0_39_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13604_ _03358_ _03359_ _03527_ _03528_ VGND VGND VPWR VPWR _03742_ sky130_fd_sc_hd__and4_1
XFILLER_0_67_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10816_ _00772_ VGND VGND VPWR VPWR _00909_ sky130_fd_sc_hd__buf_6
X_17372_ _07714_ _07715_ _07712_ VGND VGND VPWR VPWR _07843_ sky130_fd_sc_hd__a21oi_1
X_14584_ _04643_ _04644_ VGND VGND VPWR VPWR _04813_ sky130_fd_sc_hd__and2b_1
X_11796_ _01885_ _01886_ _01881_ _01884_ VGND VGND VPWR VPWR _01889_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_28_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_144_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16323_ _03047_ _06499_ VGND VGND VPWR VPWR _06702_ sky130_fd_sc_hd__or2_1
XFILLER_0_137_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13535_ _03660_ _03665_ VGND VGND VPWR VPWR _03666_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_153_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10747_ _05671_ _00459_ _00838_ _00839_ _05388_ VGND VGND VPWR VPWR _00840_ sky130_fd_sc_hd__a32oi_2
XFILLER_0_40_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16254_ _03152_ _06622_ _06625_ _06626_ VGND VGND VPWR VPWR _06627_ sky130_fd_sc_hd__o211a_1
X_13466_ _03520_ _03498_ _05311_ cla_inst.in1\[17\] VGND VGND VPWR VPWR _03590_ sky130_fd_sc_hd__and4_4
X_10678_ cla_inst.in2\[19\] cla_inst.in2\[17\] ApproximateM_inst.lob_16.lob1.genblk1\[7\].genblk1.mux.sel
+ ApproximateM_inst.lob_16.lob1.genblk1\[5\].genblk1.mux.sel VGND VGND VPWR VPWR _00771_
+ sky130_fd_sc_hd__and4_2
XFILLER_0_36_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_152_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15205_ _02999_ _00339_ VGND VGND VPWR VPWR _05490_ sky130_fd_sc_hd__nand2_1
XFILLER_0_51_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12417_ _02484_ _02509_ VGND VGND VPWR VPWR _02510_ sky130_fd_sc_hd__xnor2_1
X_16185_ _03027_ _06420_ _06549_ _06551_ _02779_ VGND VGND VPWR VPWR _06552_ sky130_fd_sc_hd__a2111o_1
X_13397_ _03512_ _03513_ _03333_ _03335_ VGND VGND VPWR VPWR _03515_ sky130_fd_sc_hd__a211o_1
XFILLER_0_23_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15136_ _04409_ _05409_ _05413_ _05414_ VGND VGND VPWR VPWR _05415_ sky130_fd_sc_hd__o211a_4
X_12348_ _02435_ _02440_ VGND VGND VPWR VPWR _02441_ sky130_fd_sc_hd__or2_1
XFILLER_0_23_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15067_ _05331_ _05338_ VGND VGND VPWR VPWR _05339_ sky130_fd_sc_hd__or2_1
X_12279_ _02260_ _02371_ VGND VGND VPWR VPWR _02372_ sky130_fd_sc_hd__nor2_1
X_14018_ _04030_ _04036_ VGND VGND VPWR VPWR _04194_ sky130_fd_sc_hd__and2b_1
XFILLER_0_65_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18826_ _09329_ VGND VGND VPWR VPWR _00099_ sky130_fd_sc_hd__clkbuf_1
X_18757_ _09275_ VGND VGND VPWR VPWR _00077_ sky130_fd_sc_hd__buf_1
X_15969_ _03920_ _05095_ _06316_ VGND VGND VPWR VPWR _06317_ sky130_fd_sc_hd__a21oi_2
X_17708_ _08097_ _08084_ VGND VGND VPWR VPWR _08209_ sky130_fd_sc_hd__or2b_1
X_09490_ _03553_ _03563_ _03695_ VGND VGND VPWR VPWR _03957_ sky130_fd_sc_hd__a21o_1
XFILLER_0_78_727 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18688_ _01671_ _09183_ _09191_ VGND VGND VPWR VPWR _09223_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_81_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17639_ _08132_ _08133_ _06589_ VGND VGND VPWR VPWR _08134_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_93_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_147_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_129_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_830 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_131_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09826_ _07602_ VGND VGND VPWR VPWR _07613_ sky130_fd_sc_hd__clkbuf_8
X_09757_ _06819_ _06830_ _06852_ VGND VGND VPWR VPWR _06863_ sky130_fd_sc_hd__a21o_1
XTAP_2104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09688_ _06073_ _06105_ VGND VGND VPWR VPWR _06116_ sky130_fd_sc_hd__and2b_1
XTAP_2137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_900 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11650_ cla_inst.in2\[20\] _07646_ _09354_ _00877_ VGND VGND VPWR VPWR _01743_ sky130_fd_sc_hd__a22o_1
XTAP_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_154_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10601_ _00661_ _00662_ _00692_ _00693_ VGND VGND VPWR VPWR _00694_ sky130_fd_sc_hd__and4bb_2
XFILLER_0_36_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11581_ _00515_ _01671_ VGND VGND VPWR VPWR _01674_ sky130_fd_sc_hd__nor2_4
XFILLER_0_147_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10532_ _04646_ _04438_ _08757_ _05246_ VGND VGND VPWR VPWR _00625_ sky130_fd_sc_hd__nand4_2
X_13320_ _03426_ _03427_ _03254_ _03256_ VGND VGND VPWR VPWR _03430_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_91_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_135_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10463_ _00554_ _00539_ _00540_ VGND VGND VPWR VPWR _00556_ sky130_fd_sc_hd__or3_1
XFILLER_0_51_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13251_ _03353_ _03354_ VGND VGND VPWR VPWR _03355_ sky130_fd_sc_hd__or2_4
XFILLER_0_122_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12202_ _02230_ _02282_ net129 _02294_ VGND VGND VPWR VPWR _02295_ sky130_fd_sc_hd__a211oi_4
X_13182_ _07058_ _00502_ VGND VGND VPWR VPWR _03282_ sky130_fd_sc_hd__nand2_1
X_10394_ _00484_ _00485_ _00482_ _00483_ VGND VGND VPWR VPWR _00487_ sky130_fd_sc_hd__o211ai_4
X_12133_ _02190_ _02192_ VGND VGND VPWR VPWR _02226_ sky130_fd_sc_hd__nand2_1
X_17990_ _08512_ _08513_ _08514_ VGND VGND VPWR VPWR _08516_ sky130_fd_sc_hd__a21o_1
X_12064_ _02070_ _02153_ _02148_ _02152_ VGND VGND VPWR VPWR _02157_ sky130_fd_sc_hd__a211oi_1
X_16941_ _02973_ _07370_ _07372_ _06484_ VGND VGND VPWR VPWR _07373_ sky130_fd_sc_hd__o211a_1
X_11015_ _07799_ _05715_ VGND VGND VPWR VPWR _01108_ sky130_fd_sc_hd__and2_4
X_16872_ _07200_ _07296_ VGND VGND VPWR VPWR _07298_ sky130_fd_sc_hd__or2_1
X_18611_ net283 _09157_ _09165_ _09162_ VGND VGND VPWR VPWR _00026_ sky130_fd_sc_hd__o211a_1
X_15823_ _06153_ _06160_ VGND VGND VPWR VPWR _06161_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_126_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18542_ net24 _09110_ _09111_ VGND VGND VPWR VPWR _09113_ sky130_fd_sc_hd__nor3_2
X_15754_ _06061_ _06063_ VGND VGND VPWR VPWR _06086_ sky130_fd_sc_hd__or2b_1
XFILLER_0_99_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12966_ _03054_ _03058_ _03050_ VGND VGND VPWR VPWR _03059_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14705_ _04943_ _04944_ VGND VGND VPWR VPWR _04945_ sky130_fd_sc_hd__nor2_2
XFILLER_0_87_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11917_ _01924_ _01923_ VGND VGND VPWR VPWR _02010_ sky130_fd_sc_hd__nand2_1
X_18473_ _08999_ _09002_ VGND VGND VPWR VPWR _09039_ sky130_fd_sc_hd__nand2_1
X_15685_ _06010_ _06011_ VGND VGND VPWR VPWR _06012_ sky130_fd_sc_hd__or2_1
XTAP_2660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12897_ _02985_ _02987_ _02988_ _02989_ VGND VGND VPWR VPWR _02990_ sky130_fd_sc_hd__or4_1
XTAP_2671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_900 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17424_ _07821_ _07786_ _07899_ VGND VGND VPWR VPWR _07900_ sky130_fd_sc_hd__o21ba_2
XTAP_2682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14636_ _03006_ _00716_ VGND VGND VPWR VPWR _04869_ sky130_fd_sc_hd__nand2_1
XFILLER_0_51_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11848_ _01938_ _01939_ _01940_ VGND VGND VPWR VPWR _01941_ sky130_fd_sc_hd__or3_1
XTAP_1970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17355_ _07091_ _06753_ _07780_ VGND VGND VPWR VPWR _07824_ sky130_fd_sc_hd__and3_1
XFILLER_0_144_106 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14567_ _04776_ _04664_ _04793_ VGND VGND VPWR VPWR _04794_ sky130_fd_sc_hd__a21oi_4
X_11779_ _01844_ _01871_ VGND VGND VPWR VPWR _01872_ sky130_fd_sc_hd__or2b_1
XFILLER_0_55_465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16306_ _06427_ _06429_ _06682_ VGND VGND VPWR VPWR _06683_ sky130_fd_sc_hd__a21oi_1
X_13518_ _03622_ _03623_ _03646_ VGND VGND VPWR VPWR _03647_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_125_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17286_ _07747_ _07748_ VGND VGND VPWR VPWR _07749_ sky130_fd_sc_hd__nand2_1
X_14498_ _04716_ _04717_ VGND VGND VPWR VPWR _04718_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_70_424 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16237_ _03117_ _03035_ _03121_ _06590_ _06607_ VGND VGND VPWR VPWR _06608_ sky130_fd_sc_hd__o311a_1
XFILLER_0_140_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_695 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13449_ _03570_ _03157_ _02983_ VGND VGND VPWR VPWR _03571_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16168_ ApproximateM_inst.lob_16.lob1.genblk1\[7\].genblk1.mux.sel sel_op\[0\] VGND
+ VGND VPWR VPWR _06533_ sky130_fd_sc_hd__or2b_1
XFILLER_0_140_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15119_ _05310_ _05395_ VGND VGND VPWR VPWR _05396_ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16099_ _06415_ _06416_ _06421_ _06457_ VGND VGND VPWR VPWR _06458_ sky130_fd_sc_hd__a31o_1
X_09611_ ApproximateM_inst.lob_16.lob2.genblk1\[10\].genblk1.mux.sel VGND VGND VPWR
+ VPWR _05279_ sky130_fd_sc_hd__buf_4
X_18809_ _01417_ net53 _09301_ VGND VGND VPWR VPWR _09316_ sky130_fd_sc_hd__mux2_1
X_09542_ _04438_ _04460_ _04482_ _04515_ VGND VGND VPWR VPWR _04526_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_78_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09473_ ApproximateM_inst.lob_16.lob2.genblk2.mux_final.sel VGND VGND VPWR VPWR _03771_
+ sky130_fd_sc_hd__buf_6
XFILLER_0_65_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_108_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_129_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_150_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_132_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09809_ _07080_ _07406_ _07112_ _07047_ VGND VGND VPWR VPWR _07428_ sky130_fd_sc_hd__a22o_1
X_12820_ _01492_ _01494_ _02911_ _02912_ VGND VGND VPWR VPWR _02913_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_69_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12751_ _02633_ _02671_ _02842_ _02843_ _02590_ VGND VGND VPWR VPWR _02844_ sky130_fd_sc_hd__o32a_4
XTAP_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11702_ _01764_ _01792_ _01794_ VGND VGND VPWR VPWR _01795_ sky130_fd_sc_hd__o21ai_2
X_15470_ _05674_ _05776_ _05777_ VGND VGND VPWR VPWR _05778_ sky130_fd_sc_hd__nor3_1
XTAP_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12682_ _02762_ _02773_ _02774_ VGND VGND VPWR VPWR _02775_ sky130_fd_sc_hd__a21o_1
XFILLER_0_49_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14421_ _04632_ _04633_ VGND VGND VPWR VPWR _04634_ sky130_fd_sc_hd__nor2_1
XTAP_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11633_ _01722_ _01723_ _01724_ VGND VGND VPWR VPWR _01726_ sky130_fd_sc_hd__a21o_1
XFILLER_0_65_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_112_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17140_ _07485_ _07491_ VGND VGND VPWR VPWR _07589_ sky130_fd_sc_hd__or2_1
XFILLER_0_64_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14352_ _03921_ _04557_ VGND VGND VPWR VPWR _04559_ sky130_fd_sc_hd__nor2_1
X_11564_ _01082_ _01081_ ApproximateM_inst.lob_16.lob1.genblk1\[14\].genblk1.mux.sel
+ ApproximateM_inst.lob_16.lob1.genblk1\[13\].genblk1.mux.sel VGND VGND VPWR VPWR
+ _01657_ sky130_fd_sc_hd__and4_1
XFILLER_0_64_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13303_ _06040_ _06051_ _07733_ VGND VGND VPWR VPWR _03412_ sky130_fd_sc_hd__and3_1
X_10515_ _00604_ _00605_ _00606_ VGND VGND VPWR VPWR _00608_ sky130_fd_sc_hd__a21o_1
X_17071_ _07512_ _07513_ VGND VGND VPWR VPWR _07514_ sky130_fd_sc_hd__and2b_1
XFILLER_0_150_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14283_ _04309_ _04473_ _04483_ VGND VGND VPWR VPWR _04484_ sky130_fd_sc_hd__o21ai_1
X_11495_ _01571_ _01570_ VGND VGND VPWR VPWR _01588_ sky130_fd_sc_hd__and2b_1
XFILLER_0_134_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16022_ _04034_ VGND VGND VPWR VPWR _06374_ sky130_fd_sc_hd__clkbuf_4
X_10446_ _00384_ _00393_ VGND VGND VPWR VPWR _00539_ sky130_fd_sc_hd__and2b_1
X_13234_ _00690_ _00692_ _03335_ _03336_ VGND VGND VPWR VPWR _03337_ sky130_fd_sc_hd__a211o_2
XFILLER_0_122_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_676 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10377_ _05366_ _05704_ _05606_ _05410_ VGND VGND VPWR VPWR _00470_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13165_ _03240_ _03241_ _03261_ _03262_ VGND VGND VPWR VPWR _03264_ sky130_fd_sc_hd__and4_2
X_12116_ _09219_ _02205_ _02208_ VGND VGND VPWR VPWR _02209_ sky130_fd_sc_hd__a21oi_1
X_17973_ _08449_ _08400_ _08495_ VGND VGND VPWR VPWR _08498_ sky130_fd_sc_hd__or3_1
X_13096_ _01863_ _03188_ _03022_ VGND VGND VPWR VPWR _03189_ sky130_fd_sc_hd__o21a_1
X_12047_ _02059_ _09354_ _02139_ VGND VGND VPWR VPWR _02140_ sky130_fd_sc_hd__nand3_1
X_16924_ _06673_ VGND VGND VPWR VPWR _07355_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_137_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16855_ _02776_ _02834_ _02968_ VGND VGND VPWR VPWR _07280_ sky130_fd_sc_hd__a21oi_1
X_15806_ _03910_ _03924_ _02981_ VGND VGND VPWR VPWR _06143_ sky130_fd_sc_hd__mux2_1
X_16786_ _07107_ _07202_ VGND VGND VPWR VPWR _07204_ sky130_fd_sc_hd__and2_1
X_13998_ _04024_ _04041_ _04042_ VGND VGND VPWR VPWR _04172_ sky130_fd_sc_hd__or3_1
XFILLER_0_87_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18525_ _06421_ _09082_ _09083_ _09090_ _09094_ VGND VGND VPWR VPWR _09095_ sky130_fd_sc_hd__a311o_1
XFILLER_0_99_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15737_ _05994_ _06067_ VGND VGND VPWR VPWR _06068_ sky130_fd_sc_hd__nor2_1
XFILLER_0_88_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12949_ _03025_ _03041_ _01674_ VGND VGND VPWR VPWR _03042_ sky130_fd_sc_hd__a21o_1
XFILLER_0_153_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_141_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18456_ _08980_ _08982_ _08979_ VGND VGND VPWR VPWR _09021_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_8_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15668_ _02994_ _05652_ _05992_ VGND VGND VPWR VPWR _05993_ sky130_fd_sc_hd__and3_1
XTAP_2490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_180 _02646_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17407_ _07731_ _07767_ _07880_ VGND VGND VPWR VPWR _07881_ sky130_fd_sc_hd__o21ai_1
X_14619_ _04841_ _04843_ _04848_ VGND VGND VPWR VPWR _04850_ sky130_fd_sc_hd__a21o_1
XFILLER_0_117_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18387_ _08909_ _08910_ VGND VGND VPWR VPWR _08946_ sky130_fd_sc_hd__or2b_1
XFILLER_0_55_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15599_ _05916_ _05917_ VGND VGND VPWR VPWR _05918_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17338_ _04853_ _06370_ _06371_ VGND VGND VPWR VPWR _07806_ sky130_fd_sc_hd__nand3_1
XFILLER_0_16_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_126_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17269_ _07718_ _07728_ VGND VGND VPWR VPWR _07730_ sky130_fd_sc_hd__or2_1
XFILLER_0_70_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19008_ clknet_4_5_0_clk _09375_ VGND VGND VPWR VPWR salida\[61\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_192 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_140_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09525_ ApproximateM_inst.lob_16.lob2.genblk1\[13\].genblk1.mux.sel VGND VGND VPWR
+ VPWR _04340_ sky130_fd_sc_hd__buf_4
XFILLER_0_149_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09456_ _03574_ _03432_ VGND VGND VPWR VPWR _03585_ sky130_fd_sc_hd__and2_1
XFILLER_0_66_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_80 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_148_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_108_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_571 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_722 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_632 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10300_ _00385_ _00392_ VGND VGND VPWR VPWR _00393_ sky130_fd_sc_hd__xor2_1
X_11280_ _01368_ _01369_ _01238_ _01273_ VGND VGND VPWR VPWR _01373_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_120_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10231_ _00321_ _00323_ VGND VGND VPWR VPWR _00324_ sky130_fd_sc_hd__nor2_1
XFILLER_0_104_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_120_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10162_ _00184_ _00183_ _03618_ _00171_ VGND VGND VPWR VPWR _00255_ sky130_fd_sc_hd__and4_1
X_14970_ _05231_ _05232_ VGND VGND VPWR VPWR _05233_ sky130_fd_sc_hd__nor2_1
X_10093_ _00170_ _00172_ _00182_ _00185_ VGND VGND VPWR VPWR _00186_ sky130_fd_sc_hd__and4_1
X_13921_ _04087_ VGND VGND VPWR VPWR _09381_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16640_ _07031_ _07044_ VGND VGND VPWR VPWR _07045_ sky130_fd_sc_hd__xnor2_1
X_13852_ _04010_ _04011_ VGND VGND VPWR VPWR _04013_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_88_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12803_ _01483_ _01469_ _01484_ VGND VGND VPWR VPWR _02896_ sky130_fd_sc_hd__or3_1
XFILLER_0_97_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16571_ _06527_ _06877_ _06969_ VGND VGND VPWR VPWR _06970_ sky130_fd_sc_hd__and3_1
X_13783_ _03755_ _03757_ _03756_ VGND VGND VPWR VPWR _03937_ sky130_fd_sc_hd__a21bo_1
X_10995_ _07973_ _08746_ _06613_ _07984_ VGND VGND VPWR VPWR _01088_ sky130_fd_sc_hd__a22o_1
XFILLER_0_29_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18310_ _08785_ _08791_ _08861_ VGND VGND VPWR VPWR _08863_ sky130_fd_sc_hd__and3_1
XTAP_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15522_ _05833_ VGND VGND VPWR VPWR _05835_ sky130_fd_sc_hd__inv_2
XFILLER_0_97_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12734_ _02803_ _02819_ VGND VGND VPWR VPWR _02827_ sky130_fd_sc_hd__xor2_1
XFILLER_0_32_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18241_ _07608_ _07861_ _08638_ VGND VGND VPWR VPWR _08788_ sky130_fd_sc_hd__or3_1
XFILLER_0_154_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15453_ _03006_ _03044_ VGND VGND VPWR VPWR _05760_ sky130_fd_sc_hd__nand2_1
XTAP_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_368 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12665_ _02721_ _02755_ VGND VGND VPWR VPWR _02758_ sky130_fd_sc_hd__and2_1
XTAP_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_700 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14404_ _04614_ _01575_ _07537_ _04615_ VGND VGND VPWR VPWR _04616_ sky130_fd_sc_hd__and4b_1
X_11616_ _01166_ _01177_ _01176_ VGND VGND VPWR VPWR _01709_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_93_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18172_ _08629_ _08711_ _08698_ VGND VGND VPWR VPWR _08714_ sky130_fd_sc_hd__and3_1
X_15384_ _05677_ _05684_ VGND VGND VPWR VPWR _05685_ sky130_fd_sc_hd__or2_1
X_12596_ _02647_ _02686_ VGND VGND VPWR VPWR _02689_ sky130_fd_sc_hd__and2_1
X_17123_ _00787_ _06331_ _06365_ _07084_ _07571_ VGND VGND VPWR VPWR _07572_ sky130_fd_sc_hd__a311oi_1
XFILLER_0_142_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14335_ _04538_ _04539_ _04426_ _04385_ VGND VGND VPWR VPWR _04541_ sky130_fd_sc_hd__o211a_1
X_11547_ _01621_ _01638_ _01639_ VGND VGND VPWR VPWR _01640_ sky130_fd_sc_hd__nor3_4
X_17054_ _07494_ _07495_ VGND VGND VPWR VPWR _07496_ sky130_fd_sc_hd__or2_1
X_14266_ _00644_ _04125_ _04130_ VGND VGND VPWR VPWR _04465_ sky130_fd_sc_hd__and3_1
XFILLER_0_12_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11478_ _00806_ _05290_ _00949_ _03421_ VGND VGND VPWR VPWR _01571_ sky130_fd_sc_hd__and4_1
XFILLER_0_111_816 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_150_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16005_ _02533_ _00214_ VGND VGND VPWR VPWR _06355_ sky130_fd_sc_hd__or2_2
XFILLER_0_150_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13217_ _01356_ _00213_ _00728_ _00727_ VGND VGND VPWR VPWR _03319_ sky130_fd_sc_hd__a31o_1
X_10429_ _07635_ _00193_ VGND VGND VPWR VPWR _00522_ sky130_fd_sc_hd__nand2_1
X_14197_ _04387_ _04388_ _04389_ VGND VGND VPWR VPWR _04390_ sky130_fd_sc_hd__nor3_1
XFILLER_0_122_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13148_ _05747_ _09311_ VGND VGND VPWR VPWR _03246_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13079_ _02685_ _03170_ _03023_ VGND VGND VPWR VPWR _03171_ sky130_fd_sc_hd__o21ai_1
X_17956_ _08477_ _08478_ VGND VGND VPWR VPWR _08479_ sky130_fd_sc_hd__and2_1
X_16907_ _06665_ _07332_ _07335_ VGND VGND VPWR VPWR _07336_ sky130_fd_sc_hd__or3_4
X_17887_ _08292_ _08348_ _08402_ VGND VGND VPWR VPWR _08404_ sky130_fd_sc_hd__nor3_1
XFILLER_0_79_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16838_ _07259_ _07260_ VGND VGND VPWR VPWR _07261_ sky130_fd_sc_hd__or2_1
XFILLER_0_88_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16769_ _03916_ _06503_ _07185_ _06645_ VGND VGND VPWR VPWR _07186_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_87_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18508_ _06303_ _06416_ VGND VGND VPWR VPWR _09076_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18439_ _06277_ _09000_ _04995_ _07592_ _09001_ VGND VGND VPWR VPWR _09002_ sky130_fd_sc_hd__o311a_1
XFILLER_0_29_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_120 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09508_ _03410_ VGND VGND VPWR VPWR _04154_ sky130_fd_sc_hd__buf_4
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10780_ cla_inst.in2\[23\] _00129_ ApproximateM_inst.lob_16.lob1.genblk1\[2\].genblk1.mux.sel
+ cla_inst.in2\[24\] VGND VGND VPWR VPWR _00873_ sky130_fd_sc_hd__a22o_1
XFILLER_0_137_702 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09439_ _03388_ VGND VGND VPWR VPWR _03399_ sky130_fd_sc_hd__clkbuf_4
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12450_ _02491_ _02497_ _02496_ VGND VGND VPWR VPWR _02543_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_35_744 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11401_ _01452_ _01453_ _01492_ _01493_ VGND VGND VPWR VPWR _01494_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_152_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12381_ _05747_ _00193_ _02473_ _02424_ VGND VGND VPWR VPWR _02474_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_105_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_80 _07766_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_91 _08880_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14120_ _04303_ _04304_ VGND VGND VPWR VPWR _04305_ sky130_fd_sc_hd__or2_1
X_11332_ _00169_ _00146_ _00872_ _00873_ VGND VGND VPWR VPWR _01425_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_105_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_698 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14051_ _04089_ _04090_ _04228_ _04229_ VGND VGND VPWR VPWR _04230_ sky130_fd_sc_hd__a211oi_2
X_11263_ _09353_ VGND VGND VPWR VPWR _01356_ sky130_fd_sc_hd__clkbuf_8
X_13002_ _00167_ _03094_ _02505_ VGND VGND VPWR VPWR _03095_ sky130_fd_sc_hd__mux2_1
X_10214_ _08605_ _08626_ VGND VGND VPWR VPWR _00307_ sky130_fd_sc_hd__nand2_1
X_11194_ _01278_ _01275_ _01276_ VGND VGND VPWR VPWR _01287_ sky130_fd_sc_hd__and3_1
X_17810_ _08318_ _08319_ VGND VGND VPWR VPWR _08320_ sky130_fd_sc_hd__nand2_1
X_10145_ _09349_ _00181_ _00197_ _00109_ VGND VGND VPWR VPWR _00238_ sky130_fd_sc_hd__a22o_1
X_18790_ _09250_ VGND VGND VPWR VPWR _09301_ sky130_fd_sc_hd__clkbuf_4
X_17741_ _06462_ _08242_ _08244_ VGND VGND VPWR VPWR _08245_ sky130_fd_sc_hd__or3_1
X_14953_ _02986_ _09311_ VGND VGND VPWR VPWR _05215_ sky130_fd_sc_hd__nand2_1
X_10076_ cla_inst.in2\[22\] VGND VGND VPWR VPWR _00169_ sky130_fd_sc_hd__buf_2
X_13904_ _03900_ _03901_ _04069_ VGND VGND VPWR VPWR _04070_ sky130_fd_sc_hd__a21o_1
XFILLER_0_89_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17672_ _08054_ _08061_ _08168_ VGND VGND VPWR VPWR _08170_ sky130_fd_sc_hd__a21bo_1
X_14884_ _05034_ VGND VGND VPWR VPWR _05140_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16623_ _07613_ _06541_ _07026_ VGND VGND VPWR VPWR _07027_ sky130_fd_sc_hd__and3_1
X_13835_ _03989_ _03992_ _03986_ VGND VGND VPWR VPWR _03994_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_69_140 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16554_ _06427_ _06651_ _06951_ VGND VGND VPWR VPWR _06952_ sky130_fd_sc_hd__or3_1
XFILLER_0_97_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13766_ _03913_ _03918_ VGND VGND VPWR VPWR _03919_ sky130_fd_sc_hd__nor2_1
X_10978_ _00990_ _00996_ VGND VGND VPWR VPWR _01071_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_128_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15505_ _00107_ _07744_ _05814_ _05815_ VGND VGND VPWR VPWR _05816_ sky130_fd_sc_hd__and4_1
XFILLER_0_85_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12717_ _02489_ _02779_ _02809_ VGND VGND VPWR VPWR _02810_ sky130_fd_sc_hd__or3b_1
X_16485_ _06567_ _06570_ _06807_ _00357_ VGND VGND VPWR VPWR _06877_ sky130_fd_sc_hd__o211a_1
X_13697_ _03841_ _03842_ VGND VGND VPWR VPWR _03843_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_57_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18224_ _08762_ _08765_ _08769_ _08770_ VGND VGND VPWR VPWR _08771_ sky130_fd_sc_hd__and4b_1
X_15436_ _02996_ _00495_ _00339_ _02993_ VGND VGND VPWR VPWR _05741_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_72_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12648_ _02701_ _02703_ _02702_ VGND VGND VPWR VPWR _02741_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_143_716 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_127_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18155_ _08665_ _08666_ VGND VGND VPWR VPWR _08695_ sky130_fd_sc_hd__and2_1
XFILLER_0_4_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15367_ _05653_ _05585_ _05664_ VGND VGND VPWR VPWR _05666_ sky130_fd_sc_hd__and3_1
XFILLER_0_142_226 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12579_ _02644_ _02645_ _02651_ VGND VGND VPWR VPWR _02672_ sky130_fd_sc_hd__nand3_1
XFILLER_0_81_883 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17106_ _07324_ _07326_ _07436_ _07438_ VGND VGND VPWR VPWR _07553_ sky130_fd_sc_hd__o31ai_2
X_14318_ _04516_ _04521_ VGND VGND VPWR VPWR _04522_ sky130_fd_sc_hd__xnor2_1
X_18086_ _07313_ _07410_ _07486_ _07593_ VGND VGND VPWR VPWR _08620_ sky130_fd_sc_hd__or4_1
XFILLER_0_13_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15298_ _00591_ _03154_ VGND VGND VPWR VPWR _05591_ sky130_fd_sc_hd__nand2_2
XFILLER_0_1_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17037_ _06425_ _06437_ _07469_ _07473_ _07477_ VGND VGND VPWR VPWR _07478_ sky130_fd_sc_hd__o311a_1
X_14249_ _04442_ _04443_ _04444_ VGND VGND VPWR VPWR _04446_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09790_ ApproximateM_inst.lob_16.lob2.genblk1\[4\].genblk1.mux.sel VGND VGND VPWR
+ VPWR _07221_ sky130_fd_sc_hd__buf_4
XTAP_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18988_ clknet_4_6_0_clk _09384_ VGND VGND VPWR VPWR salida\[41\] sky130_fd_sc_hd__dfxtp_1
XTAP_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17939_ _07042_ _08260_ VGND VGND VPWR VPWR _08460_ sky130_fd_sc_hd__nor2_1
XFILLER_0_84_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_419 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_368 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_146_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_755 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_552 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_134_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_141_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09988_ _09271_ _09279_ VGND VGND VPWR VPWR _09295_ sky130_fd_sc_hd__or2_1
X_11950_ _02028_ _02041_ VGND VGND VPWR VPWR _02043_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_87_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwb_buttons_leds_154 VGND VGND VPWR VPWR wb_buttons_leds_154/HI led_enb[3] sky130_fd_sc_hd__conb_1
X_10901_ _05638_ _05028_ _04569_ _00992_ VGND VGND VPWR VPWR _00994_ sky130_fd_sc_hd__a22o_1
XFILLER_0_98_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11881_ _01971_ _01972_ _01960_ _01968_ VGND VGND VPWR VPWR _01974_ sky130_fd_sc_hd__o211a_1
X_13620_ _03755_ _03756_ _03757_ VGND VGND VPWR VPWR _03758_ sky130_fd_sc_hd__nand3_2
X_10832_ _00918_ _00919_ _00924_ VGND VGND VPWR VPWR _00925_ sky130_fd_sc_hd__nor3b_2
XFILLER_0_104_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13551_ _00170_ _00715_ _03475_ _03474_ VGND VGND VPWR VPWR _03683_ sky130_fd_sc_hd__a31o_1
X_10763_ _00823_ _00854_ _08311_ _00855_ VGND VGND VPWR VPWR _00856_ sky130_fd_sc_hd__o211a_4
XFILLER_0_109_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12502_ _07036_ _07069_ _00130_ _00871_ VGND VGND VPWR VPWR _02595_ sky130_fd_sc_hd__nand4_2
XFILLER_0_125_705 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16270_ _06636_ _06643_ _03538_ VGND VGND VPWR VPWR _06644_ sky130_fd_sc_hd__o21a_1
X_13482_ _03603_ _03604_ _03605_ VGND VGND VPWR VPWR _03608_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_35_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10694_ _04427_ _03804_ VGND VGND VPWR VPWR _00787_ sky130_fd_sc_hd__nand2_4
XFILLER_0_70_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15221_ _05387_ _05505_ VGND VGND VPWR VPWR _05507_ sky130_fd_sc_hd__or2_1
X_12433_ _02524_ _02523_ _02525_ VGND VGND VPWR VPWR _02526_ sky130_fd_sc_hd__nor3_1
XFILLER_0_120_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15152_ _05326_ _05328_ VGND VGND VPWR VPWR _05432_ sky130_fd_sc_hd__and2_1
XFILLER_0_23_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12364_ _02385_ _02388_ _02387_ VGND VGND VPWR VPWR _02457_ sky130_fd_sc_hd__o21a_1
XFILLER_0_23_758 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14103_ _04103_ _04104_ _04102_ VGND VGND VPWR VPWR _04287_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_50_555 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11315_ net139 _01405_ _01306_ _01304_ VGND VGND VPWR VPWR _01408_ sky130_fd_sc_hd__o211a_1
X_15083_ _05354_ _05356_ VGND VGND VPWR VPWR _05357_ sky130_fd_sc_hd__or2_1
XFILLER_0_120_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12295_ _02282_ _02384_ _02352_ net323 VGND VGND VPWR VPWR _02388_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_120_443 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14034_ _04191_ _04210_ _04211_ VGND VGND VPWR VPWR _04212_ sky130_fd_sc_hd__or3_2
X_18911_ clknet_4_10_0_clk _00065_ VGND VGND VPWR VPWR cla_inst.in1\[29\] sky130_fd_sc_hd__dfxtp_1
X_11246_ _01241_ _01258_ VGND VGND VPWR VPWR _01339_ sky130_fd_sc_hd__and2_1
XFILLER_0_38_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18842_ clknet_4_0_0_clk net251 VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__dfxtp_1
X_11177_ _01252_ _01269_ VGND VGND VPWR VPWR _01270_ sky130_fd_sc_hd__xnor2_1
X_10128_ _00170_ _00206_ _00216_ _00219_ VGND VGND VPWR VPWR _00221_ sky130_fd_sc_hd__o2bb2a_1
X_18773_ _09288_ VGND VGND VPWR VPWR _00082_ sky130_fd_sc_hd__clkbuf_1
X_15985_ _07711_ _00357_ VGND VGND VPWR VPWR _06333_ sky130_fd_sc_hd__or2_2
X_10059_ _00149_ _00131_ _00127_ _00151_ VGND VGND VPWR VPWR _00152_ sky130_fd_sc_hd__a22o_1
X_14936_ _05194_ _05195_ VGND VGND VPWR VPWR _05197_ sky130_fd_sc_hd__nand2_1
X_17724_ _02467_ _08226_ _02326_ VGND VGND VPWR VPWR _08227_ sky130_fd_sc_hd__a21o_1
X_14867_ _05119_ _05120_ VGND VGND VPWR VPWR _05121_ sky130_fd_sc_hd__or2_1
X_17655_ _02977_ _06753_ _07859_ _08150_ _06762_ VGND VGND VPWR VPWR _08151_ sky130_fd_sc_hd__a32o_1
X_13818_ _03796_ _03798_ VGND VGND VPWR VPWR _03975_ sky130_fd_sc_hd__nand2_1
X_16606_ _03537_ _03197_ _04076_ _06680_ _07008_ VGND VGND VPWR VPWR _07009_ sky130_fd_sc_hd__a311o_1
X_17586_ _08066_ _08074_ _08075_ VGND VGND VPWR VPWR _08076_ sky130_fd_sc_hd__nor3_1
X_14798_ _05044_ _05043_ VGND VGND VPWR VPWR _05046_ sky130_fd_sc_hd__or2b_1
X_16537_ _06933_ VGND VGND VPWR VPWR _09413_ sky130_fd_sc_hd__inv_2
X_13749_ _03897_ _03899_ VGND VGND VPWR VPWR _03900_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_45_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16468_ _06425_ _06851_ _06853_ _06856_ _06858_ VGND VGND VPWR VPWR _06859_ sky130_fd_sc_hd__o311a_1
XFILLER_0_45_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_658 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15419_ _02991_ _08876_ _05721_ VGND VGND VPWR VPWR _05722_ sky130_fd_sc_hd__a21oi_1
X_18207_ _04900_ _08428_ _02994_ VGND VGND VPWR VPWR _08752_ sky130_fd_sc_hd__or3b_1
XFILLER_0_60_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16399_ _06780_ _06781_ _06782_ VGND VGND VPWR VPWR _06784_ sky130_fd_sc_hd__a21o_1
XFILLER_0_53_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18138_ _08609_ _08610_ _08607_ VGND VGND VPWR VPWR _08677_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_79_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold103 _00023_ VGND VGND VPWR VPWR net266 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold114 net114 VGND VGND VPWR VPWR net277 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18069_ _06394_ _06790_ _08601_ _04647_ VGND VGND VPWR VPWR _08602_ sky130_fd_sc_hd__a22o_1
XFILLER_0_110_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold125 _00028_ VGND VGND VPWR VPWR net288 sky130_fd_sc_hd__dlygate4sd3_1
Xhold136 net87 VGND VGND VPWR VPWR net299 sky130_fd_sc_hd__dlygate4sd3_1
Xhold147 net107 VGND VGND VPWR VPWR net310 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09911_ _06277_ _06288_ _06298_ VGND VGND VPWR VPWR _08539_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_22_791 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09842_ _07700_ VGND VGND VPWR VPWR _07788_ sky130_fd_sc_hd__clkbuf_4
XTAP_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09773_ ApproximateM_inst.lob_16.lob2.genblk1\[4\].genblk1.mux.sel VGND VGND VPWR
+ VPWR _07036_ sky130_fd_sc_hd__buf_4
XTAP_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_110 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_135_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_138_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_901 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_147_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_134_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11100_ _01167_ _01170_ VGND VGND VPWR VPWR _01193_ sky130_fd_sc_hd__nand2_1
X_12080_ _02164_ _02166_ VGND VGND VPWR VPWR _02173_ sky130_fd_sc_hd__xnor2_2
X_11031_ _05671_ _04580_ _01122_ _01123_ VGND VGND VPWR VPWR _01124_ sky130_fd_sc_hd__a31o_1
X_15770_ _06101_ _06102_ VGND VGND VPWR VPWR _06103_ sky130_fd_sc_hd__xor2_1
X_12982_ _07810_ _03074_ _03024_ VGND VGND VPWR VPWR _03075_ sky130_fd_sc_hd__o21ai_1
X_14721_ _04937_ _04936_ VGND VGND VPWR VPWR _04961_ sky130_fd_sc_hd__and2b_2
XFILLER_0_99_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11933_ _01968_ _02025_ VGND VGND VPWR VPWR _02026_ sky130_fd_sc_hd__nand2_1
XTAP_2820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17440_ _06374_ _06592_ _06551_ VGND VGND VPWR VPWR _07917_ sky130_fd_sc_hd__a21o_1
X_14652_ _00253_ _05975_ VGND VGND VPWR VPWR _04887_ sky130_fd_sc_hd__nand2_4
X_11864_ _01953_ _01956_ VGND VGND VPWR VPWR _01957_ sky130_fd_sc_hd__xor2_2
XFILLER_0_39_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13603_ _03738_ _03740_ VGND VGND VPWR VPWR _03741_ sky130_fd_sc_hd__nand2_1
X_10815_ _00906_ _00907_ VGND VGND VPWR VPWR _00908_ sky130_fd_sc_hd__nor2_2
X_17371_ _07723_ _07725_ _07721_ _07018_ VGND VGND VPWR VPWR _07841_ sky130_fd_sc_hd__o2bb2a_1
X_14583_ _04809_ _04811_ VGND VGND VPWR VPWR _04812_ sky130_fd_sc_hd__xnor2_2
X_11795_ _01844_ _01870_ net199 _01869_ VGND VGND VPWR VPWR _01888_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_67_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16322_ _02982_ _06500_ _06699_ _06466_ VGND VGND VPWR VPWR _06701_ sky130_fd_sc_hd__o211a_1
XFILLER_0_137_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13534_ _03661_ _03664_ VGND VGND VPWR VPWR _03665_ sky130_fd_sc_hd__xor2_1
X_10746_ _06019_ _08039_ _08049_ VGND VGND VPWR VPWR _00839_ sky130_fd_sc_hd__and3_1
XFILLER_0_82_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16253_ _06466_ VGND VGND VPWR VPWR _06626_ sky130_fd_sc_hd__clkbuf_4
X_13465_ _03366_ _05311_ _05028_ _03345_ VGND VGND VPWR VPWR _03589_ sky130_fd_sc_hd__a22oi_2
X_10677_ _04263_ _04253_ _04231_ VGND VGND VPWR VPWR _00770_ sky130_fd_sc_hd__a21o_1
XFILLER_0_35_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15204_ _05485_ _05488_ VGND VGND VPWR VPWR _05489_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_125_568 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_691 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12416_ _02500_ _02508_ VGND VGND VPWR VPWR _02509_ sky130_fd_sc_hd__nand2_1
XFILLER_0_113_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16184_ _06550_ VGND VGND VPWR VPWR _06551_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_106_760 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13396_ _03333_ _03335_ _03512_ _03513_ VGND VGND VPWR VPWR _03514_ sky130_fd_sc_hd__o211ai_4
X_15135_ _04950_ net117 VGND VGND VPWR VPWR _05414_ sky130_fd_sc_hd__nand2_2
XFILLER_0_49_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12347_ _02437_ _02438_ _02439_ VGND VGND VPWR VPWR _02440_ sky130_fd_sc_hd__or3_1
XFILLER_0_121_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15066_ _05335_ _05337_ VGND VGND VPWR VPWR _05338_ sky130_fd_sc_hd__or2_1
X_12278_ _07711_ _00247_ _02370_ VGND VGND VPWR VPWR _02371_ sky130_fd_sc_hd__and3_1
XFILLER_0_121_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14017_ _04028_ _04039_ VGND VGND VPWR VPWR _04193_ sky130_fd_sc_hd__nand2_1
XFILLER_0_120_284 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11229_ _00835_ _01321_ VGND VGND VPWR VPWR _01322_ sky130_fd_sc_hd__and2b_1
X_18825_ _09125_ _09328_ VGND VGND VPWR VPWR _09329_ sky130_fd_sc_hd__and2_1
XFILLER_0_65_34 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18756_ _09273_ _09274_ VGND VGND VPWR VPWR _09275_ sky130_fd_sc_hd__and2_1
X_15968_ _03920_ _05097_ VGND VGND VPWR VPWR _06316_ sky130_fd_sc_hd__nor2_1
X_17707_ _08206_ _08207_ VGND VGND VPWR VPWR _08208_ sky130_fd_sc_hd__nor2_1
X_14919_ _05176_ _05177_ VGND VGND VPWR VPWR _05178_ sky130_fd_sc_hd__and2_1
X_18687_ _09222_ VGND VGND VPWR VPWR _00053_ sky130_fd_sc_hd__clkbuf_1
X_15899_ _06211_ _06241_ VGND VGND VPWR VPWR _06242_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17638_ _08023_ _08027_ VGND VGND VPWR VPWR _08133_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17569_ _07944_ _08056_ VGND VGND VPWR VPWR _08057_ sky130_fd_sc_hd__nor2_1
XFILLER_0_19_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_496 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_128_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_128_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_719 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_842 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09825_ _07591_ VGND VGND VPWR VPWR _07602_ sky130_fd_sc_hd__clkbuf_8
X_09756_ _05551_ _05791_ _06841_ VGND VGND VPWR VPWR _06852_ sky130_fd_sc_hd__a21o_1
XTAP_2105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09687_ _06084_ _06094_ _05257_ _06040_ VGND VGND VPWR VPWR _06105_ sky130_fd_sc_hd__a22o_1
XTAP_2116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10600_ _00690_ _00691_ _00507_ _00528_ VGND VGND VPWR VPWR _00693_ sky130_fd_sc_hd__a211o_1
XFILLER_0_92_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11580_ _01106_ _01671_ _01672_ VGND VGND VPWR VPWR _01673_ sky130_fd_sc_hd__or3b_4
XFILLER_0_25_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10531_ _04373_ _05617_ _05246_ _04351_ VGND VGND VPWR VPWR _00624_ sky130_fd_sc_hd__a22o_1
XFILLER_0_64_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_107_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13250_ _00752_ _00754_ VGND VGND VPWR VPWR _03354_ sky130_fd_sc_hd__nor2_1
XFILLER_0_134_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10462_ _00539_ _00540_ _00554_ VGND VGND VPWR VPWR _00555_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12201_ _02287_ _02291_ _02292_ _02290_ VGND VGND VPWR VPWR _02294_ sky130_fd_sc_hd__o22a_1
XFILLER_0_60_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13181_ _00639_ _00642_ _00640_ VGND VGND VPWR VPWR _03280_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_33_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10393_ _00482_ _00483_ _00484_ _00485_ VGND VGND VPWR VPWR _00486_ sky130_fd_sc_hd__a211o_1
XFILLER_0_0_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12132_ _02223_ _02210_ _02221_ VGND VGND VPWR VPWR _02225_ sky130_fd_sc_hd__and3_1
XFILLER_0_102_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16940_ _02972_ _07371_ VGND VGND VPWR VPWR _07372_ sky130_fd_sc_hd__nand2_1
X_12063_ _02135_ _02155_ VGND VGND VPWR VPWR _02156_ sky130_fd_sc_hd__nand2_1
X_11014_ _01106_ _00514_ _06776_ _00309_ VGND VGND VPWR VPWR _01107_ sky130_fd_sc_hd__or4b_4
X_16871_ _07285_ _07295_ VGND VGND VPWR VPWR _07296_ sky130_fd_sc_hd__xnor2_1
X_18610_ salida\[22\] _09159_ _09160_ salida\[54\] _09163_ VGND VGND VPWR VPWR _09165_
+ sky130_fd_sc_hd__a221o_1
X_15822_ _06157_ _06158_ VGND VGND VPWR VPWR _06160_ sky130_fd_sc_hd__nor2_1
X_18541_ net13 net2 VGND VGND VPWR VPWR _09111_ sky130_fd_sc_hd__or2_2
XFILLER_0_87_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15753_ _04823_ _06081_ _06082_ _06085_ VGND VGND VPWR VPWR _09370_ sky130_fd_sc_hd__a31o_1
X_12965_ _03024_ _03057_ VGND VGND VPWR VPWR _03058_ sky130_fd_sc_hd__nand2_1
XFILLER_0_99_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14704_ _04814_ _04812_ VGND VGND VPWR VPWR _04944_ sky130_fd_sc_hd__and2b_1
X_11916_ _02007_ _02008_ VGND VGND VPWR VPWR _02009_ sky130_fd_sc_hd__or2_1
X_15684_ _05955_ _06009_ VGND VGND VPWR VPWR _06011_ sky130_fd_sc_hd__and2_1
X_18472_ _03108_ _04853_ _08150_ VGND VGND VPWR VPWR _09038_ sky130_fd_sc_hd__and3_1
X_12896_ _04099_ VGND VGND VPWR VPWR _02989_ sky130_fd_sc_hd__clkbuf_8
XTAP_2650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17423_ _07896_ _07898_ VGND VGND VPWR VPWR _07899_ sky130_fd_sc_hd__xnor2_1
X_14635_ _04865_ _04866_ _04737_ _04739_ VGND VGND VPWR VPWR _04868_ sky130_fd_sc_hd__a211o_4
XFILLER_0_68_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11847_ _01917_ _01918_ VGND VGND VPWR VPWR _01940_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_142_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14566_ _04791_ _04792_ VGND VGND VPWR VPWR _04793_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17354_ _07710_ _07716_ VGND VGND VPWR VPWR _07823_ sky130_fd_sc_hd__or2b_1
XFILLER_0_28_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11778_ net199 _01869_ _01844_ _01870_ VGND VGND VPWR VPWR _01871_ sky130_fd_sc_hd__a211o_1
XFILLER_0_126_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13517_ _03644_ _03645_ VGND VGND VPWR VPWR _03646_ sky130_fd_sc_hd__nor2_1
X_16305_ _06424_ _06430_ VGND VGND VPWR VPWR _06682_ sky130_fd_sc_hd__or2_1
X_10729_ _06149_ _06159_ _06170_ _05181_ VGND VGND VPWR VPWR _00822_ sky130_fd_sc_hd__a22o_1
X_17285_ _06581_ _07621_ _07742_ _07746_ VGND VGND VPWR VPWR _07748_ sky130_fd_sc_hd__a2bb2o_1
X_14497_ _04001_ _09248_ VGND VGND VPWR VPWR _04717_ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16236_ _06600_ _06604_ _06606_ VGND VGND VPWR VPWR _06607_ sky130_fd_sc_hd__and3_1
X_13448_ _03162_ VGND VGND VPWR VPWR _03570_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_152_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16167_ _00217_ _00909_ VGND VGND VPWR VPWR _06532_ sky130_fd_sc_hd__or2_1
X_13379_ _01356_ _00166_ _03326_ _03325_ VGND VGND VPWR VPWR _03495_ sky130_fd_sc_hd__a31o_1
X_15118_ _05392_ _05394_ VGND VGND VPWR VPWR _05395_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_62_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16098_ _06426_ _06453_ _06456_ VGND VGND VPWR VPWR _06457_ sky130_fd_sc_hd__o21ai_1
X_15049_ _05317_ _05318_ VGND VGND VPWR VPWR _05319_ sky130_fd_sc_hd__xnor2_1
X_09610_ _05235_ _05257_ VGND VGND VPWR VPWR _05268_ sky130_fd_sc_hd__nand2_1
X_18808_ _09315_ VGND VGND VPWR VPWR _00093_ sky130_fd_sc_hd__clkbuf_1
X_09541_ _04504_ VGND VGND VPWR VPWR _04515_ sky130_fd_sc_hd__buf_4
X_18739_ _03117_ net61 _09251_ VGND VGND VPWR VPWR _09261_ sky130_fd_sc_hd__mux2_1
X_09472_ _03728_ _03750_ VGND VGND VPWR VPWR _03760_ sky130_fd_sc_hd__nand2_4
XFILLER_0_148_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_148_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_116_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_132_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_131_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_132_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_112_560 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09808_ _07232_ _07254_ _07406_ _07102_ VGND VGND VPWR VPWR _07417_ sky130_fd_sc_hd__and4_1
X_09739_ _06646_ _06656_ VGND VGND VPWR VPWR _06667_ sky130_fd_sc_hd__xor2_1
XFILLER_0_96_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12750_ _02669_ _02670_ _02632_ VGND VGND VPWR VPWR _02843_ sky130_fd_sc_hd__o21a_1
XTAP_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11701_ _01251_ _01793_ VGND VGND VPWR VPWR _01794_ sky130_fd_sc_hd__nor2_1
XTAP_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12681_ _02768_ _02772_ _02739_ _02763_ VGND VGND VPWR VPWR _02774_ sky130_fd_sc_hd__o211a_1
XTAP_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14420_ _00195_ _00702_ _05845_ _00443_ VGND VGND VPWR VPWR _04633_ sky130_fd_sc_hd__and4_1
XTAP_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11632_ _01722_ _01723_ _01724_ VGND VGND VPWR VPWR _01725_ sky130_fd_sc_hd__nand3_1
XFILLER_0_139_479 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14351_ _03131_ _03178_ _03080_ VGND VGND VPWR VPWR _04557_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11563_ _01081_ ApproximateM_inst.lob_16.lob1.genblk1\[14\].genblk1.mux.sel ApproximateM_inst.lob_16.lob1.genblk1\[13\].genblk1.mux.sel
+ _01082_ VGND VGND VPWR VPWR _01656_ sky130_fd_sc_hd__a22o_1
XFILLER_0_80_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13302_ _03226_ _03234_ _03233_ VGND VGND VPWR VPWR _03411_ sky130_fd_sc_hd__a21o_1
X_10514_ _00604_ _00605_ _00606_ VGND VGND VPWR VPWR _00607_ sky130_fd_sc_hd__nand3_1
X_17070_ net334 _07124_ _07126_ _07511_ VGND VGND VPWR VPWR _07513_ sky130_fd_sc_hd__or4_1
X_14282_ _04480_ _04481_ VGND VGND VPWR VPWR _04483_ sky130_fd_sc_hd__and2_1
XFILLER_0_108_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11494_ _05224_ _04056_ VGND VGND VPWR VPWR _01587_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16021_ _06370_ _06371_ _04853_ VGND VGND VPWR VPWR _06372_ sky130_fd_sc_hd__a21bo_1
X_13233_ _03333_ _03334_ _03314_ VGND VGND VPWR VPWR _03336_ sky130_fd_sc_hd__o21a_1
X_10445_ _00396_ _00397_ _00415_ VGND VGND VPWR VPWR _00538_ sky130_fd_sc_hd__nand3_1
XFILLER_0_150_688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13164_ _03240_ _03241_ _03261_ _03262_ VGND VGND VPWR VPWR _03263_ sky130_fd_sc_hd__a22oi_2
X_10376_ _00299_ _00300_ VGND VGND VPWR VPWR _00469_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12115_ _08713_ _00131_ _02206_ _02207_ VGND VGND VPWR VPWR _02208_ sky130_fd_sc_hd__and4_1
X_17972_ _08449_ _08400_ _08495_ VGND VGND VPWR VPWR _08497_ sky130_fd_sc_hd__o21ai_1
X_13095_ _02505_ _01671_ VGND VGND VPWR VPWR _03188_ sky130_fd_sc_hd__nor2_1
X_12046_ _02088_ _02138_ VGND VGND VPWR VPWR _02139_ sky130_fd_sc_hd__and2_1
X_16923_ _02751_ _02836_ VGND VGND VPWR VPWR _07354_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16854_ _03198_ _04414_ _07266_ _07278_ VGND VGND VPWR VPWR _07279_ sky130_fd_sc_hd__a211o_1
X_15805_ _02976_ _04241_ _04415_ _03036_ VGND VGND VPWR VPWR _06142_ sky130_fd_sc_hd__a31o_1
X_13997_ _04041_ VGND VGND VPWR VPWR _04171_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16785_ _07107_ _07202_ VGND VGND VPWR VPWR _07203_ sky130_fd_sc_hd__nor2_1
X_18524_ _03201_ _09092_ _09093_ VGND VGND VPWR VPWR _09094_ sky130_fd_sc_hd__and3_1
X_12948_ _01695_ VGND VGND VPWR VPWR _03041_ sky130_fd_sc_hd__clkbuf_4
X_15736_ _06065_ _06066_ VGND VGND VPWR VPWR _06067_ sky130_fd_sc_hd__or2_1
XFILLER_0_87_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18455_ _09018_ _09019_ VGND VGND VPWR VPWR _09020_ sky130_fd_sc_hd__or2b_1
X_12879_ _07058_ VGND VGND VPWR VPWR _02972_ sky130_fd_sc_hd__buf_4
X_15667_ _02997_ _03154_ VGND VGND VPWR VPWR _05992_ sky130_fd_sc_hd__nand2_1
XANTENNA_170 _02646_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_181 _02646_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17406_ _07878_ _07879_ VGND VGND VPWR VPWR _07880_ sky130_fd_sc_hd__nor2_1
XFILLER_0_134_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14618_ _04841_ _04843_ _04848_ VGND VGND VPWR VPWR _04849_ sky130_fd_sc_hd__nand3_1
X_15598_ _02994_ _02997_ _04125_ _03153_ VGND VGND VPWR VPWR _05917_ sky130_fd_sc_hd__and4_1
X_18386_ _03068_ _06464_ _08924_ _08945_ VGND VGND VPWR VPWR _09405_ sky130_fd_sc_hd__o2bb2a_1
XTAP_1790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14549_ _01873_ _01112_ VGND VGND VPWR VPWR _04774_ sky130_fd_sc_hd__nand2_1
X_17337_ _07801_ _07802_ _07803_ VGND VGND VPWR VPWR _07805_ sky130_fd_sc_hd__a21o_1
XFILLER_0_16_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_756 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_114_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17268_ _07718_ _07728_ VGND VGND VPWR VPWR _07729_ sky130_fd_sc_hd__nand2_1
XFILLER_0_102_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_110 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19007_ clknet_4_7_0_clk _09374_ VGND VGND VPWR VPWR salida\[60\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16219_ _06586_ _06587_ _06513_ VGND VGND VPWR VPWR _06588_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_114_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17199_ _07652_ _07531_ _07653_ VGND VGND VPWR VPWR _07654_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_3_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09524_ _04023_ _04110_ _04165_ VGND VGND VPWR VPWR _04329_ sky130_fd_sc_hd__o21ba_2
XFILLER_0_66_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09455_ _03454_ VGND VGND VPWR VPWR _03574_ sky130_fd_sc_hd__buf_4
XFILLER_0_78_388 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_789 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_116_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10230_ _08865_ _00322_ _00317_ _00320_ VGND VGND VPWR VPWR _00323_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_14_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10161_ _00253_ _00212_ VGND VGND VPWR VPWR _00254_ sky130_fd_sc_hd__nand2_1
XFILLER_0_100_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10092_ _00183_ _00177_ _00146_ _00184_ VGND VGND VPWR VPWR _00185_ sky130_fd_sc_hd__a22o_1
XFILLER_0_100_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13920_ _04074_ _04086_ VGND VGND VPWR VPWR _04087_ sky130_fd_sc_hd__or2_1
X_13851_ _00170_ _04591_ VGND VGND VPWR VPWR _04011_ sky130_fd_sc_hd__nand2_1
XFILLER_0_69_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12802_ _00592_ _00881_ _01481_ _01479_ VGND VGND VPWR VPWR _02895_ sky130_fd_sc_hd__a31o_1
X_13782_ _03574_ _00459_ _03932_ _03933_ VGND VGND VPWR VPWR _03936_ sky130_fd_sc_hd__a22o_1
X_16570_ _06968_ VGND VGND VPWR VPWR _06969_ sky130_fd_sc_hd__clkbuf_4
X_10994_ _07036_ _07069_ _08746_ _06613_ VGND VGND VPWR VPWR _01087_ sky130_fd_sc_hd__nand4_1
XFILLER_0_97_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15521_ _02993_ _02996_ _00665_ _03071_ VGND VGND VPWR VPWR _05833_ sky130_fd_sc_hd__and4_1
X_12733_ _02823_ _02825_ VGND VGND VPWR VPWR _02826_ sky130_fd_sc_hd__and2_1
XTAP_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15452_ _05755_ _05756_ _05717_ _05718_ VGND VGND VPWR VPWR _05759_ sky130_fd_sc_hd__o211ai_2
XTAP_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18240_ _06368_ _07390_ _08700_ _08699_ VGND VGND VPWR VPWR _08787_ sky130_fd_sc_hd__a31o_1
XTAP_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12664_ _00845_ _00134_ _02720_ VGND VGND VPWR VPWR _02757_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_139_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14403_ _07504_ _03750_ _04012_ _00358_ VGND VGND VPWR VPWR _04615_ sky130_fd_sc_hd__a22o_1
XFILLER_0_53_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11615_ _01166_ _01176_ _01177_ VGND VGND VPWR VPWR _01708_ sky130_fd_sc_hd__or3_4
XFILLER_0_127_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15383_ _05681_ _05683_ VGND VGND VPWR VPWR _05684_ sky130_fd_sc_hd__xor2_1
XFILLER_0_5_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18171_ _08629_ _08698_ _08711_ VGND VGND VPWR VPWR _08712_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_143_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12595_ _07700_ _00194_ _02646_ VGND VGND VPWR VPWR _02688_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_154_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14334_ _04426_ _04385_ _04538_ _04539_ VGND VGND VPWR VPWR _04540_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_107_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17122_ _00787_ _06331_ _06365_ VGND VGND VPWR VPWR _07571_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_142_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11546_ _01619_ _01620_ _01605_ _01606_ VGND VGND VPWR VPWR _01639_ sky130_fd_sc_hd__o211a_1
XFILLER_0_53_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17053_ _07388_ _07492_ VGND VGND VPWR VPWR _07495_ sky130_fd_sc_hd__and2_1
X_14265_ _04287_ _04291_ _04292_ _04294_ _04286_ VGND VGND VPWR VPWR _04464_ sky130_fd_sc_hd__a32o_1
X_11477_ _06591_ _03476_ _00210_ _00806_ VGND VGND VPWR VPWR _01570_ sky130_fd_sc_hd__a22o_1
X_16004_ _06338_ _06350_ _06353_ _06339_ VGND VGND VPWR VPWR _06354_ sky130_fd_sc_hd__a211o_1
XFILLER_0_0_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13216_ _01503_ _00511_ _00684_ _00686_ VGND VGND VPWR VPWR _03318_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_110_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_828 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10428_ _00134_ _00359_ _00520_ VGND VGND VPWR VPWR _00521_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_20_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14196_ _04214_ _04216_ VGND VGND VPWR VPWR _04389_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13147_ _07744_ _03243_ _03244_ VGND VGND VPWR VPWR _03245_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_103_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10359_ _04427_ _06613_ _08049_ _04504_ VGND VGND VPWR VPWR _00452_ sky130_fd_sc_hd__a22o_1
XFILLER_0_148_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13078_ _03026_ _03169_ VGND VGND VPWR VPWR _03170_ sky130_fd_sc_hd__and2_1
X_17955_ _08475_ _08476_ _08352_ _08471_ VGND VGND VPWR VPWR _08478_ sky130_fd_sc_hd__o211ai_1
X_12029_ _02108_ _02121_ VGND VGND VPWR VPWR _02122_ sky130_fd_sc_hd__or2_1
X_16906_ _07333_ _07334_ VGND VGND VPWR VPWR _07335_ sky130_fd_sc_hd__xor2_1
X_17886_ _08292_ _08348_ _08402_ VGND VGND VPWR VPWR _08403_ sky130_fd_sc_hd__o21a_1
XFILLER_0_79_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16837_ _07168_ _07170_ _07165_ VGND VGND VPWR VPWR _07260_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_87_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16768_ _07183_ _07184_ _03920_ VGND VGND VPWR VPWR _07185_ sky130_fd_sc_hd__mux2_1
X_18507_ _03011_ _06512_ _03155_ VGND VGND VPWR VPWR _09075_ sky130_fd_sc_hd__a21boi_1
X_15719_ _06046_ _06047_ VGND VGND VPWR VPWR _06048_ sky130_fd_sc_hd__xnor2_1
X_16699_ _07108_ VGND VGND VPWR VPWR _07109_ sky130_fd_sc_hd__clkbuf_4
X_18438_ _09000_ _04995_ _06277_ VGND VGND VPWR VPWR _09001_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_146_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18369_ _08925_ _08926_ VGND VGND VPWR VPWR _08927_ sky130_fd_sc_hd__and2b_1
XFILLER_0_16_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_132 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09507_ _03914_ VGND VGND VPWR VPWR _04143_ sky130_fd_sc_hd__buf_4
XFILLER_0_149_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_336 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_109_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_714 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09438_ ApproximateM_inst.lob_16.lob1.genblk1\[10\].genblk1.mux.sel VGND VGND VPWR
+ VPWR _03388_ sky130_fd_sc_hd__buf_4
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_583 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11400_ _01490_ _01491_ _01415_ _01454_ VGND VGND VPWR VPWR _01493_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_124_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12380_ _02423_ VGND VGND VPWR VPWR _02473_ sky130_fd_sc_hd__inv_2
XANTENNA_70 _05845_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_81 _07810_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11331_ cla_inst.in2\[21\] _00223_ VGND VGND VPWR VPWR _01424_ sky130_fd_sc_hd__nand2_1
XANTENNA_92 _08880_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14050_ _04225_ _04226_ _04227_ VGND VGND VPWR VPWR _04229_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_132_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11262_ _01353_ _01354_ VGND VGND VPWR VPWR _01355_ sky130_fd_sc_hd__xor2_4
XFILLER_0_30_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13001_ _00214_ VGND VGND VPWR VPWR _03094_ sky130_fd_sc_hd__clkbuf_4
X_10213_ _08539_ _08594_ VGND VGND VPWR VPWR _00306_ sky130_fd_sc_hd__or2b_1
X_11193_ _01284_ _01285_ VGND VGND VPWR VPWR _01286_ sky130_fd_sc_hd__nand2_1
X_10144_ _00109_ _09349_ _00146_ _00197_ VGND VGND VPWR VPWR _00237_ sky130_fd_sc_hd__and4_1
XFILLER_0_100_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17740_ _03119_ _05621_ _06705_ _08243_ VGND VGND VPWR VPWR _08244_ sky130_fd_sc_hd__a2bb2o_1
X_14952_ _05211_ _05212_ VGND VGND VPWR VPWR _05214_ sky130_fd_sc_hd__nor2_1
X_10075_ _00164_ _00167_ VGND VGND VPWR VPWR _00168_ sky130_fd_sc_hd__nand2_2
X_13903_ _03900_ _03901_ _03738_ VGND VGND VPWR VPWR _04069_ sky130_fd_sc_hd__o21a_1
X_17671_ _08052_ _08053_ VGND VGND VPWR VPWR _08168_ sky130_fd_sc_hd__nand2_1
X_14883_ _05136_ _05138_ VGND VGND VPWR VPWR _05139_ sky130_fd_sc_hd__nor2_1
X_16622_ _07023_ _07024_ _06040_ VGND VGND VPWR VPWR _07026_ sky130_fd_sc_hd__o21a_2
X_13834_ _03986_ _03989_ _03992_ VGND VGND VPWR VPWR _03993_ sky130_fd_sc_hd__or3_2
XFILLER_0_43_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16553_ _06802_ _06806_ _03535_ VGND VGND VPWR VPWR _06951_ sky130_fd_sc_hd__a21o_2
X_13765_ _03164_ _03066_ VGND VGND VPWR VPWR _03918_ sky130_fd_sc_hd__nor2_2
X_10977_ _01044_ _01047_ VGND VGND VPWR VPWR _01070_ sky130_fd_sc_hd__nand2_1
XFILLER_0_69_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15504_ _03322_ _03321_ _08224_ _08158_ VGND VGND VPWR VPWR _05815_ sky130_fd_sc_hd__nand4_4
XFILLER_0_85_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12716_ _02785_ _02806_ _02808_ VGND VGND VPWR VPWR _02809_ sky130_fd_sc_hd__o21a_1
XFILLER_0_128_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13696_ _00169_ _04700_ VGND VGND VPWR VPWR _03842_ sky130_fd_sc_hd__nand2_1
X_16484_ _06563_ _06875_ VGND VGND VPWR VPWR _06876_ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18223_ _03198_ _06083_ _07184_ _08141_ VGND VGND VPWR VPWR _08770_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_127_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15435_ _05659_ _05658_ VGND VGND VPWR VPWR _05740_ sky130_fd_sc_hd__or2b_1
X_12647_ _02701_ _02702_ _02703_ VGND VGND VPWR VPWR _02740_ sky130_fd_sc_hd__and3_1
XFILLER_0_128_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15366_ _05653_ _05585_ _05664_ VGND VGND VPWR VPWR _05665_ sky130_fd_sc_hd__a21oi_1
X_18154_ _03052_ _06463_ _08672_ _08694_ VGND VGND VPWR VPWR _09401_ sky130_fd_sc_hd__a22oi_2
X_12578_ _02669_ _02670_ VGND VGND VPWR VPWR _02671_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_80_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_142_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17105_ _07549_ _07551_ VGND VGND VPWR VPWR _07552_ sky130_fd_sc_hd__xnor2_1
X_14317_ _04519_ _04520_ VGND VGND VPWR VPWR _04521_ sky130_fd_sc_hd__xnor2_1
X_11529_ _01185_ _01183_ _01184_ VGND VGND VPWR VPWR _01622_ sky130_fd_sc_hd__nand3_1
X_15297_ _05588_ _05589_ VGND VGND VPWR VPWR _05590_ sky130_fd_sc_hd__nand2_1
X_18085_ _07649_ _07489_ _07596_ _07664_ VGND VGND VPWR VPWR _08619_ sky130_fd_sc_hd__a22o_1
XFILLER_0_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14248_ _04442_ _04443_ _04444_ VGND VGND VPWR VPWR _04445_ sky130_fd_sc_hd__and3_2
X_17036_ _03920_ _07474_ _07476_ _06645_ VGND VGND VPWR VPWR _07477_ sky130_fd_sc_hd__a211o_1
XFILLER_0_68_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14179_ _04158_ _04368_ VGND VGND VPWR VPWR _04370_ sky130_fd_sc_hd__nand2_1
XTAP_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18987_ clknet_4_6_0_clk _09383_ VGND VGND VPWR VPWR salida\[40\] sky130_fd_sc_hd__dfxtp_1
XTAP_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17938_ _07130_ _07706_ VGND VGND VPWR VPWR _08459_ sky130_fd_sc_hd__nor2_1
XFILLER_0_30_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17869_ _07302_ _07741_ VGND VGND VPWR VPWR _08384_ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_483 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_656 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_767 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_564 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_895 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110_680 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09987_ _09271_ _09279_ VGND VGND VPWR VPWR _09287_ sky130_fd_sc_hd__nand2_1
XFILLER_0_99_715 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10900_ _00992_ _05638_ _04569_ VGND VGND VPWR VPWR _00993_ sky130_fd_sc_hd__and3_1
Xwb_buttons_leds_155 VGND VGND VPWR VPWR wb_buttons_leds_155/HI led_enb[4] sky130_fd_sc_hd__conb_1
X_11880_ _01960_ _01968_ net193 _01972_ VGND VGND VPWR VPWR _01973_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_86_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10831_ _00922_ _00923_ VGND VGND VPWR VPWR _00924_ sky130_fd_sc_hd__xnor2_1
X_13550_ _03680_ _03681_ VGND VGND VPWR VPWR _03682_ sky130_fd_sc_hd__xor2_2
XFILLER_0_13_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10762_ _08278_ _08289_ _08300_ _06938_ VGND VGND VPWR VPWR _00855_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_149_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12501_ _02550_ _02555_ _02554_ VGND VGND VPWR VPWR _02594_ sky130_fd_sc_hd__a21o_1
XFILLER_0_137_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13481_ _03603_ _03604_ _03605_ VGND VGND VPWR VPWR _03606_ sky130_fd_sc_hd__and3_2
X_10693_ _04635_ _03739_ VGND VGND VPWR VPWR _00786_ sky130_fd_sc_hd__nand2_4
XFILLER_0_152_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15220_ _05387_ _05505_ VGND VGND VPWR VPWR _05506_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12432_ _02456_ _02522_ _02515_ net122 VGND VGND VPWR VPWR _02525_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_81_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15151_ _05223_ _05329_ VGND VGND VPWR VPWR _05430_ sky130_fd_sc_hd__or2_1
XFILLER_0_63_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12363_ _02450_ _02454_ _02455_ VGND VGND VPWR VPWR _02456_ sky130_fd_sc_hd__or3_4
X_14102_ _04112_ _04113_ VGND VGND VPWR VPWR _04286_ sky130_fd_sc_hd__or2_2
X_11314_ _01304_ _01306_ _01405_ net139 VGND VGND VPWR VPWR _01407_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_133_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15082_ _09352_ _00309_ _05352_ _05353_ VGND VGND VPWR VPWR _05356_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_50_567 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_105_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12294_ _02263_ _02386_ VGND VGND VPWR VPWR _02387_ sky130_fd_sc_hd__xor2_1
XFILLER_0_31_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14033_ _04192_ _04193_ _04207_ VGND VGND VPWR VPWR _04211_ sky130_fd_sc_hd__and3_1
X_18910_ clknet_4_8_0_clk _00064_ VGND VGND VPWR VPWR cla_inst.in1\[28\] sky130_fd_sc_hd__dfxtp_4
XFILLER_0_31_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11245_ _01120_ _01144_ _01118_ VGND VGND VPWR VPWR _01338_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_120_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_120_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18841_ clknet_4_0_0_clk net260 VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__dfxtp_1
X_11176_ _01267_ _01268_ VGND VGND VPWR VPWR _01269_ sky130_fd_sc_hd__nor2_1
X_10127_ _00216_ _00219_ _00170_ _00206_ VGND VGND VPWR VPWR _00220_ sky130_fd_sc_hd__and4bb_1
X_18772_ _09273_ _09286_ VGND VGND VPWR VPWR _09288_ sky130_fd_sc_hd__and2_1
X_15984_ _06993_ _00108_ VGND VGND VPWR VPWR _06332_ sky130_fd_sc_hd__or2_1
X_17723_ _02849_ _02846_ VGND VGND VPWR VPWR _08226_ sky130_fd_sc_hd__or2b_1
X_10058_ cla_inst.in2\[27\] VGND VGND VPWR VPWR _00151_ sky130_fd_sc_hd__clkbuf_4
X_14935_ _05194_ _05195_ VGND VGND VPWR VPWR _05196_ sky130_fd_sc_hd__or2_1
XFILLER_0_89_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17654_ _07825_ VGND VGND VPWR VPWR _08150_ sky130_fd_sc_hd__clkbuf_4
X_14866_ _04986_ _04990_ _05118_ VGND VGND VPWR VPWR _05120_ sky130_fd_sc_hd__and3_1
XFILLER_0_58_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16605_ _06345_ _06545_ _07007_ _03169_ VGND VGND VPWR VPWR _07008_ sky130_fd_sc_hd__a22o_1
X_13817_ _03972_ _03973_ VGND VGND VPWR VPWR _03974_ sky130_fd_sc_hd__xnor2_2
X_17585_ _08067_ _07947_ _08073_ VGND VGND VPWR VPWR _08075_ sky130_fd_sc_hd__nor3_1
X_14797_ _05043_ _05044_ VGND VGND VPWR VPWR _05045_ sky130_fd_sc_hd__or2b_1
X_16536_ _06904_ _06907_ _06932_ _06463_ _03086_ VGND VGND VPWR VPWR _06933_ sky130_fd_sc_hd__a32o_2
X_13748_ _03368_ _03693_ _03692_ _03898_ VGND VGND VPWR VPWR _03899_ sky130_fd_sc_hd__a31o_1
XFILLER_0_57_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16467_ _06349_ _06338_ _06348_ _06598_ _06857_ VGND VGND VPWR VPWR _06858_ sky130_fd_sc_hd__a311o_1
X_13679_ _03817_ _03820_ _03822_ VGND VGND VPWR VPWR _03823_ sky130_fd_sc_hd__or3_2
XFILLER_0_73_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18206_ _02994_ _06511_ _06776_ VGND VGND VPWR VPWR _08751_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_143_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15418_ _09350_ _07015_ VGND VGND VPWR VPWR _05721_ sky130_fd_sc_hd__and2_1
XFILLER_0_26_553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16398_ _06780_ _06781_ _06782_ VGND VGND VPWR VPWR _06783_ sky130_fd_sc_hd__nand3_1
XFILLER_0_143_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18137_ _03052_ _08428_ _02997_ VGND VGND VPWR VPWR _08676_ sky130_fd_sc_hd__or3b_1
X_15349_ _05644_ _05645_ VGND VGND VPWR VPWR _05646_ sky130_fd_sc_hd__nor2_1
XFILLER_0_53_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold104 net102 VGND VGND VPWR VPWR net267 sky130_fd_sc_hd__dlygate4sd3_1
Xhold115 _00013_ VGND VGND VPWR VPWR net278 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18068_ _02998_ _06920_ _06921_ VGND VGND VPWR VPWR _08601_ sky130_fd_sc_hd__a21o_1
Xhold126 net90 VGND VGND VPWR VPWR net289 sky130_fd_sc_hd__dlygate4sd3_1
Xhold137 _00017_ VGND VGND VPWR VPWR net300 sky130_fd_sc_hd__dlygate4sd3_1
Xhold148 net105 VGND VGND VPWR VPWR net311 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09910_ _08496_ _08507_ _08518_ VGND VGND VPWR VPWR _08529_ sky130_fd_sc_hd__and3_2
X_17019_ _02968_ _07457_ VGND VGND VPWR VPWR _07458_ sky130_fd_sc_hd__or2_1
XFILLER_0_1_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09841_ _07711_ _07744_ _07766_ VGND VGND VPWR VPWR _07777_ sky130_fd_sc_hd__nand3_1
XTAP_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09772_ _07015_ VGND VGND VPWR VPWR _07025_ sky130_fd_sc_hd__clkbuf_8
XTAP_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_280 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_134_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_383 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_761 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_731 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11030_ _00992_ _08039_ _04449_ _04471_ VGND VGND VPWR VPWR _01123_ sky130_fd_sc_hd__and4_1
X_12981_ _03025_ _03073_ VGND VGND VPWR VPWR _03074_ sky130_fd_sc_hd__and2_1
X_14720_ _04953_ _04954_ _04956_ _03125_ _04960_ VGND VGND VPWR VPWR _09357_ sky130_fd_sc_hd__a221o_1
X_11932_ _01965_ _01966_ _01967_ _01961_ VGND VGND VPWR VPWR _02025_ sky130_fd_sc_hd__o31ai_1
XTAP_2810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14651_ _04764_ _04765_ VGND VGND VPWR VPWR _04885_ sky130_fd_sc_hd__nand2_1
X_11863_ _01954_ _01955_ VGND VGND VPWR VPWR _01956_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_39_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13602_ _03736_ _03737_ VGND VGND VPWR VPWR _03740_ sky130_fd_sc_hd__nand2_1
X_10814_ _00761_ _00905_ VGND VGND VPWR VPWR _00907_ sky130_fd_sc_hd__and2_1
X_17370_ _07823_ _07839_ VGND VGND VPWR VPWR _07840_ sky130_fd_sc_hd__xor2_1
X_14582_ _04678_ _04681_ VGND VGND VPWR VPWR _04811_ sky130_fd_sc_hd__nor2_1
X_11794_ _01881_ _01884_ _01885_ _01886_ VGND VGND VPWR VPWR _01887_ sky130_fd_sc_hd__a211o_2
XFILLER_0_94_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16321_ _03047_ _06489_ VGND VGND VPWR VPWR _06699_ sky130_fd_sc_hd__or2_1
X_13533_ _02972_ _03456_ _03663_ VGND VGND VPWR VPWR _03664_ sky130_fd_sc_hd__and3_1
X_10745_ _08039_ net230 net222 _06019_ VGND VGND VPWR VPWR _00838_ sky130_fd_sc_hd__a22o_1
XFILLER_0_55_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_851 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13464_ _03454_ _05377_ VGND VGND VPWR VPWR _03588_ sky130_fd_sc_hd__nand2_8
X_16252_ _03048_ _06623_ VGND VGND VPWR VPWR _06625_ sky130_fd_sc_hd__or2_1
XFILLER_0_42_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10676_ _04263_ _04231_ _04253_ VGND VGND VPWR VPWR _00769_ sky130_fd_sc_hd__nand3_1
X_15203_ _05370_ _05487_ VGND VGND VPWR VPWR _05488_ sky130_fd_sc_hd__nor2_1
X_12415_ _02501_ _02507_ VGND VGND VPWR VPWR _02508_ sky130_fd_sc_hd__or2b_1
X_13395_ _03510_ _03511_ _03471_ _03472_ VGND VGND VPWR VPWR _03513_ sky130_fd_sc_hd__a211o_1
X_16183_ _06459_ _03292_ _03217_ VGND VGND VPWR VPWR _06550_ sky130_fd_sc_hd__and3b_1
XFILLER_0_62_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15134_ _05198_ _05201_ _05302_ _05412_ VGND VGND VPWR VPWR _05413_ sky130_fd_sc_hd__o31a_1
X_12346_ _02371_ _02436_ VGND VGND VPWR VPWR _02439_ sky130_fd_sc_hd__nor2b_1
XFILLER_0_23_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_121_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15065_ _00362_ _00461_ _05336_ _05332_ VGND VGND VPWR VPWR _05337_ sky130_fd_sc_hd__o2bb2a_1
X_12277_ _00120_ _00398_ VGND VGND VPWR VPWR _02370_ sky130_fd_sc_hd__and2_2
X_14016_ _03823_ _04038_ VGND VGND VPWR VPWR _04192_ sky130_fd_sc_hd__or2_1
XFILLER_0_121_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11228_ _06971_ _05704_ _00833_ _00834_ VGND VGND VPWR VPWR _01321_ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18824_ _06200_ net59 _09250_ VGND VGND VPWR VPWR _09328_ sky130_fd_sc_hd__mux2_1
X_11159_ _01231_ _01233_ VGND VGND VPWR VPWR _01252_ sky130_fd_sc_hd__nor2_1
XFILLER_0_65_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18755_ _02476_ net66 _09251_ VGND VGND VPWR VPWR _09274_ sky130_fd_sc_hd__mux2_1
X_15967_ _06314_ _03930_ VGND VGND VPWR VPWR _06315_ sky130_fd_sc_hd__and2_4
X_17706_ _08203_ _08205_ VGND VGND VPWR VPWR _08207_ sky130_fd_sc_hd__nor2_1
X_14918_ _00591_ _03142_ _05175_ VGND VGND VPWR VPWR _05177_ sky130_fd_sc_hd__a21o_1
X_18686_ _09209_ _09221_ VGND VGND VPWR VPWR _09222_ sky130_fd_sc_hd__and2_1
X_15898_ _06238_ _06240_ VGND VGND VPWR VPWR _06241_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_81_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17637_ _08129_ _08131_ VGND VGND VPWR VPWR _08132_ sky130_fd_sc_hd__and2_1
X_14849_ _03596_ _07755_ cla_inst.in1\[27\] _03629_ VGND VGND VPWR VPWR _05101_ sky130_fd_sc_hd__a22o_1
X_17568_ _06969_ _07596_ VGND VGND VPWR VPWR _08056_ sky130_fd_sc_hd__nand2_1
XFILLER_0_147_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_129_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16519_ _06616_ _06621_ _03099_ VGND VGND VPWR VPWR _06914_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17499_ _07207_ net146 _07664_ _06947_ VGND VGND VPWR VPWR _07981_ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_723 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_854 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09824_ _07581_ VGND VGND VPWR VPWR _07591_ sky130_fd_sc_hd__clkbuf_8
X_09755_ _05540_ _05442_ VGND VGND VPWR VPWR _06841_ sky130_fd_sc_hd__and2b_1
X_09686_ _06062_ VGND VGND VPWR VPWR _06094_ sky130_fd_sc_hd__buf_4
XTAP_2106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10530_ _04984_ _00443_ _00441_ _00440_ _04132_ VGND VGND VPWR VPWR _00623_ sky130_fd_sc_hd__a32o_1
XFILLER_0_64_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10461_ _00542_ _00553_ VGND VGND VPWR VPWR _00554_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_10_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12200_ _02287_ _02290_ _02291_ _02292_ VGND VGND VPWR VPWR _02293_ sky130_fd_sc_hd__nor4_1
XFILLER_0_33_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13180_ _00669_ _00670_ VGND VGND VPWR VPWR _03279_ sky130_fd_sc_hd__nand2_1
X_10392_ _00316_ _00324_ VGND VGND VPWR VPWR _00485_ sky130_fd_sc_hd__and2_1
XFILLER_0_103_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12131_ _02210_ _02221_ _02223_ VGND VGND VPWR VPWR _02224_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_20_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12062_ _02049_ _02107_ _02134_ VGND VGND VPWR VPWR _02155_ sky130_fd_sc_hd__or3_1
X_11013_ _01105_ VGND VGND VPWR VPWR _01106_ sky130_fd_sc_hd__buf_4
X_16870_ _07287_ _07294_ VGND VGND VPWR VPWR _07295_ sky130_fd_sc_hd__xnor2_2
X_15821_ _03016_ _03154_ _06154_ _06156_ VGND VGND VPWR VPWR _06158_ sky130_fd_sc_hd__a22oi_1
X_18540_ net28 _09109_ net27 VGND VGND VPWR VPWR _09110_ sky130_fd_sc_hd__or3b_2
X_15752_ _04264_ _05623_ _06083_ _03124_ VGND VGND VPWR VPWR _06085_ sky130_fd_sc_hd__a22o_1
X_12964_ _03027_ _03056_ _01114_ VGND VGND VPWR VPWR _03057_ sky130_fd_sc_hd__a21o_1
X_14703_ _04811_ _04809_ VGND VGND VPWR VPWR _04943_ sky130_fd_sc_hd__and2b_1
X_11915_ _01928_ _01931_ VGND VGND VPWR VPWR _02008_ sky130_fd_sc_hd__xnor2_1
X_18471_ _09007_ VGND VGND VPWR VPWR _09036_ sky130_fd_sc_hd__inv_2
X_15683_ _05955_ _06009_ VGND VGND VPWR VPWR _06010_ sky130_fd_sc_hd__nor2_1
XTAP_2640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12895_ _01520_ VGND VGND VPWR VPWR _02988_ sky130_fd_sc_hd__clkbuf_8
XTAP_2651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17422_ _06750_ _07780_ _07778_ _07776_ VGND VGND VPWR VPWR _07898_ sky130_fd_sc_hd__a31oi_2
X_14634_ _04737_ _04739_ _04865_ _04866_ VGND VGND VPWR VPWR _04867_ sky130_fd_sc_hd__o211ai_4
XTAP_2673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11846_ _01936_ _01937_ net341 _01932_ VGND VGND VPWR VPWR _01939_ sky130_fd_sc_hd__a211oi_1
XTAP_2684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17353_ _07705_ _07717_ VGND VGND VPWR VPWR _07822_ sky130_fd_sc_hd__or2b_1
X_14565_ _04778_ _04779_ _04790_ VGND VGND VPWR VPWR _04792_ sky130_fd_sc_hd__or3_1
X_11777_ _01843_ _01842_ _01841_ _01828_ VGND VGND VPWR VPWR _01870_ sky130_fd_sc_hd__o211a_1
XTAP_1994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16304_ _02981_ _06592_ _06550_ VGND VGND VPWR VPWR _06681_ sky130_fd_sc_hd__a21o_1
X_13516_ _03642_ _03643_ _03422_ _03424_ VGND VGND VPWR VPWR _03645_ sky130_fd_sc_hd__o211a_1
X_10728_ _00797_ _00819_ _00820_ VGND VGND VPWR VPWR _00821_ sky130_fd_sc_hd__nor3_2
XFILLER_0_82_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17284_ _06581_ _07621_ _07742_ _07746_ VGND VGND VPWR VPWR _07747_ sky130_fd_sc_hd__or4bb_2
X_14496_ _04714_ _04715_ VGND VGND VPWR VPWR _04716_ sky130_fd_sc_hd__nor2_1
XFILLER_0_36_670 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_126_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16235_ _02806_ _02968_ _06605_ VGND VGND VPWR VPWR _06606_ sky130_fd_sc_hd__or3b_1
XFILLER_0_36_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10659_ _00585_ _00599_ _00750_ _00751_ VGND VGND VPWR VPWR _00752_ sky130_fd_sc_hd__o211a_2
XFILLER_0_42_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13447_ _03567_ _03568_ _03098_ VGND VGND VPWR VPWR _03569_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13378_ _03319_ _03329_ _03493_ VGND VGND VPWR VPWR _03494_ sky130_fd_sc_hd__a21o_1
XFILLER_0_23_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16166_ _00211_ _06529_ _06530_ VGND VGND VPWR VPWR _06531_ sky130_fd_sc_hd__or3_2
XFILLER_0_140_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15117_ _05243_ _05287_ _05393_ VGND VGND VPWR VPWR _05394_ sky130_fd_sc_hd__o21ba_1
X_12329_ _02419_ _02421_ VGND VGND VPWR VPWR _02422_ sky130_fd_sc_hd__or2_1
XFILLER_0_50_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16097_ _03038_ _06454_ _06455_ _03120_ VGND VGND VPWR VPWR _06456_ sky130_fd_sc_hd__o22a_1
X_15048_ _02987_ _00513_ VGND VGND VPWR VPWR _05318_ sky130_fd_sc_hd__nand2_1
X_18807_ _09298_ _09314_ VGND VGND VPWR VPWR _09315_ sky130_fd_sc_hd__and2_1
X_16999_ _07316_ _07320_ _07315_ VGND VGND VPWR VPWR _07436_ sky130_fd_sc_hd__o21ba_1
X_09540_ _04493_ VGND VGND VPWR VPWR _04504_ sky130_fd_sc_hd__buf_6
X_18738_ _09260_ VGND VGND VPWR VPWR _00071_ sky130_fd_sc_hd__buf_1
X_09471_ _03739_ VGND VGND VPWR VPWR _03750_ sky130_fd_sc_hd__buf_6
X_18669_ net36 _03101_ _09193_ VGND VGND VPWR VPWR _09210_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_116_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_506 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_117_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_132_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_143_196 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_112_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_140_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09807_ cla_inst.in1\[26\] VGND VGND VPWR VPWR _07406_ sky130_fd_sc_hd__clkbuf_4
X_09738_ _05235_ _05257_ _05421_ _05344_ VGND VGND VPWR VPWR _06656_ sky130_fd_sc_hd__a31o_1
X_09669_ _05410_ _05366_ _05497_ VGND VGND VPWR VPWR _05910_ sky130_fd_sc_hd__and3_1
XTAP_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11700_ _01226_ _01250_ VGND VGND VPWR VPWR _01793_ sky130_fd_sc_hd__nor2_1
XTAP_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12680_ _02739_ _02763_ _02768_ _02772_ VGND VGND VPWR VPWR _02773_ sky130_fd_sc_hd__a211o_1
XFILLER_0_38_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11631_ _01685_ _01686_ _01684_ VGND VGND VPWR VPWR _01724_ sky130_fd_sc_hd__a21bo_1
XTAP_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11562_ _01646_ _01654_ VGND VGND VPWR VPWR _01655_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_65_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14350_ _03125_ _04414_ _04419_ _03199_ _04556_ VGND VGND VPWR VPWR _09384_ sky130_fd_sc_hd__a221o_1
XFILLER_0_80_724 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_108_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10513_ _03465_ _04460_ VGND VGND VPWR VPWR _00606_ sky130_fd_sc_hd__and2_1
X_13301_ _03406_ _03407_ _03224_ _03375_ VGND VGND VPWR VPWR _03409_ sky130_fd_sc_hd__a211o_2
XFILLER_0_64_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14281_ _04477_ _04479_ _04474_ VGND VGND VPWR VPWR _04481_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_80_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11493_ _01581_ _01584_ _01583_ VGND VGND VPWR VPWR _01586_ sky130_fd_sc_hd__a21o_1
XFILLER_0_134_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13232_ _03314_ _03333_ _03334_ VGND VGND VPWR VPWR _03335_ sky130_fd_sc_hd__nor3_4
X_16020_ _02200_ _03311_ VGND VGND VPWR VPWR _06371_ sky130_fd_sc_hd__or2_1
X_10444_ net186 _00375_ _00535_ _00536_ VGND VGND VPWR VPWR _00537_ sky130_fd_sc_hd__o211a_2
XFILLER_0_134_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13163_ _03258_ _03259_ _00651_ _00653_ VGND VGND VPWR VPWR _03262_ sky130_fd_sc_hd__o211ai_2
X_10375_ _00292_ _00298_ VGND VGND VPWR VPWR _00468_ sky130_fd_sc_hd__or2b_1
XFILLER_0_0_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12114_ _05301_ _09212_ _09188_ _05279_ VGND VGND VPWR VPWR _02207_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13094_ _02125_ _03186_ _03022_ VGND VGND VPWR VPWR _03187_ sky130_fd_sc_hd__o21a_1
X_17971_ _08484_ _08494_ VGND VGND VPWR VPWR _08495_ sky130_fd_sc_hd__xnor2_1
X_12045_ _02083_ _02087_ VGND VGND VPWR VPWR _02138_ sky130_fd_sc_hd__nand2_1
X_16922_ _02751_ _02836_ VGND VGND VPWR VPWR _07353_ sky130_fd_sc_hd__or2_1
X_16853_ _06462_ _07271_ _07273_ _07277_ VGND VGND VPWR VPWR _07278_ sky130_fd_sc_hd__or4_1
XFILLER_0_46_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15804_ _06137_ _06139_ VGND VGND VPWR VPWR _06141_ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16784_ _07200_ _07201_ VGND VGND VPWR VPWR _07202_ sky130_fd_sc_hd__nand2_1
X_13996_ _04166_ _04167_ _04168_ VGND VGND VPWR VPWR _04170_ sky130_fd_sc_hd__a21oi_1
X_18523_ _02949_ _09061_ _02956_ VGND VGND VPWR VPWR _09093_ sky130_fd_sc_hd__o21ai_1
X_15735_ _06023_ _06064_ VGND VGND VPWR VPWR _06066_ sky130_fd_sc_hd__and2_1
X_12947_ _03022_ VGND VGND VPWR VPWR _03040_ sky130_fd_sc_hd__clkbuf_4
X_18454_ _03073_ _08428_ _03013_ VGND VGND VPWR VPWR _09019_ sky130_fd_sc_hd__or3b_1
X_15666_ _05989_ _05990_ VGND VGND VPWR VPWR _05991_ sky130_fd_sc_hd__nand2_1
XTAP_2470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12878_ _00759_ _02964_ _02970_ VGND VGND VPWR VPWR _02971_ sky130_fd_sc_hd__o21ai_2
XANTENNA_160 _08762_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_171 _02646_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17405_ _07854_ _07877_ VGND VGND VPWR VPWR _07879_ sky130_fd_sc_hd__and2_1
XTAP_2492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14617_ _04846_ _04847_ VGND VGND VPWR VPWR _04848_ sky130_fd_sc_hd__xnor2_1
X_18385_ _07256_ _08929_ _08931_ _08944_ VGND VGND VPWR VPWR _08945_ sky130_fd_sc_hd__a31o_1
X_11829_ ApproximateM_inst.lob_16.lob2.genblk1\[8\].genblk1.mux.sel _03607_ VGND VGND
+ VPWR VPWR _01922_ sky130_fd_sc_hd__and2_1
X_15597_ _02997_ _04125_ _03153_ _02994_ VGND VGND VPWR VPWR _05916_ sky130_fd_sc_hd__a22oi_1
XTAP_1780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17336_ _07801_ _07802_ _07803_ VGND VGND VPWR VPWR _07804_ sky130_fd_sc_hd__nand3_1
XFILLER_0_127_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14548_ _04771_ _04772_ VGND VGND VPWR VPWR _04773_ sky130_fd_sc_hd__nor2_1
X_17267_ _07719_ _07727_ VGND VGND VPWR VPWR _07728_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_125_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14479_ _03125_ _04559_ _04563_ _03199_ _04697_ VGND VGND VPWR VPWR _09385_ sky130_fd_sc_hd__a221o_1
XFILLER_0_71_768 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_114_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19006_ clknet_4_5_0_clk _09373_ VGND VGND VPWR VPWR salida\[59\] sky130_fd_sc_hd__dfxtp_1
X_16218_ _01106_ _07646_ _06585_ VGND VGND VPWR VPWR _06587_ sky130_fd_sc_hd__or3_1
XFILLER_0_140_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17198_ _06581_ _07516_ _07512_ _07513_ VGND VGND VPWR VPWR _07653_ sky130_fd_sc_hd__o31a_1
X_16149_ _06511_ VGND VGND VPWR VPWR _06512_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_122_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09523_ _03968_ _03979_ _04307_ VGND VGND VPWR VPWR _04318_ sky130_fd_sc_hd__nand3_4
XFILLER_0_78_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09454_ _03443_ _03542_ _03487_ VGND VGND VPWR VPWR _03563_ sky130_fd_sc_hd__a21o_1
XFILLER_0_148_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_105_826 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10160_ _00169_ VGND VGND VPWR VPWR _00253_ sky130_fd_sc_hd__buf_4
X_10091_ cla_inst.in2\[24\] VGND VGND VPWR VPWR _00184_ sky130_fd_sc_hd__clkbuf_4
X_13850_ _04008_ _04009_ VGND VGND VPWR VPWR _04010_ sky130_fd_sc_hd__nor2_1
XFILLER_0_16_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12801_ _02892_ _02888_ _02889_ _02893_ VGND VGND VPWR VPWR _02894_ sky130_fd_sc_hd__o22ai_4
X_13781_ _03574_ _00459_ _03932_ _03933_ VGND VGND VPWR VPWR _03934_ sky130_fd_sc_hd__nand4_2
X_10993_ _06471_ _00993_ _00991_ _00995_ VGND VGND VPWR VPWR _01086_ sky130_fd_sc_hd__o2bb2a_1
XTAP_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15520_ _02996_ _03153_ _03071_ _02993_ VGND VGND VPWR VPWR _05832_ sky130_fd_sc_hd__a22o_1
XTAP_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12732_ _02818_ _02824_ VGND VGND VPWR VPWR _02825_ sky130_fd_sc_hd__nor2_1
XFILLER_0_139_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15451_ _05717_ _05718_ _05755_ _05756_ VGND VGND VPWR VPWR _05757_ sky130_fd_sc_hd__a211o_1
XTAP_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12663_ _02721_ _02755_ VGND VGND VPWR VPWR _02756_ sky130_fd_sc_hd__nor2_1
XFILLER_0_84_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14402_ _00358_ _07504_ _03750_ _04012_ VGND VGND VPWR VPWR _04614_ sky130_fd_sc_hd__and4_1
XTAP_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11614_ _01642_ _01704_ _01705_ _01706_ VGND VGND VPWR VPWR _01707_ sky130_fd_sc_hd__nor4_2
X_18170_ _08709_ _08710_ VGND VGND VPWR VPWR _08711_ sky130_fd_sc_hd__nand2_1
X_15382_ _03015_ _01112_ VGND VGND VPWR VPWR _05683_ sky130_fd_sc_hd__nand2_1
X_12594_ _02647_ _02686_ VGND VGND VPWR VPWR _02687_ sky130_fd_sc_hd__nor2_1
X_17121_ _07565_ _07566_ _07567_ VGND VGND VPWR VPWR _07569_ sky130_fd_sc_hd__a21o_1
XFILLER_0_25_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14333_ _04489_ _04490_ _04535_ _04536_ VGND VGND VPWR VPWR _04539_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_52_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11545_ _01636_ _01637_ VGND VGND VPWR VPWR _01638_ sky130_fd_sc_hd__nand2_1
XFILLER_0_107_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17052_ _07388_ _07492_ VGND VGND VPWR VPWR _07494_ sky130_fd_sc_hd__nor2_1
X_14264_ _04305_ _04306_ VGND VGND VPWR VPWR _04463_ sky130_fd_sc_hd__or2b_1
X_11476_ _01565_ _01567_ _01566_ VGND VGND VPWR VPWR _01569_ sky130_fd_sc_hd__a21o_1
X_16003_ _06341_ _06345_ _06352_ VGND VGND VPWR VPWR _06353_ sky130_fd_sc_hd__and3_1
X_13215_ _00724_ _00731_ _03316_ VGND VGND VPWR VPWR _03317_ sky130_fd_sc_hd__a21o_1
X_10427_ _07504_ _00131_ _09219_ _00358_ VGND VGND VPWR VPWR _00520_ sky130_fd_sc_hd__a22o_1
X_14195_ _04385_ _04386_ _04169_ net120 VGND VGND VPWR VPWR _04388_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_104_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13146_ _06051_ _00498_ _07384_ _06029_ VGND VGND VPWR VPWR _03244_ sky130_fd_sc_hd__a22o_1
X_10358_ _04351_ _00294_ _05246_ _05322_ VGND VGND VPWR VPWR _00451_ sky130_fd_sc_hd__nand4_2
XFILLER_0_0_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13077_ _00878_ VGND VGND VPWR VPWR _03169_ sky130_fd_sc_hd__clkbuf_4
X_17954_ _08352_ _08471_ _08475_ _08476_ VGND VGND VPWR VPWR _08477_ sky130_fd_sc_hd__a211o_1
X_10289_ _00241_ _00235_ VGND VGND VPWR VPWR _00382_ sky130_fd_sc_hd__and2b_1
X_12028_ _02111_ _02119_ _02120_ VGND VGND VPWR VPWR _02121_ sky130_fd_sc_hd__a21oi_1
X_16905_ _07220_ _07222_ _07219_ VGND VGND VPWR VPWR _07334_ sky130_fd_sc_hd__o21ai_2
X_17885_ _08400_ _08401_ VGND VGND VPWR VPWR _08402_ sky130_fd_sc_hd__nor2_1
X_16836_ _07257_ _07258_ VGND VGND VPWR VPWR _07259_ sky130_fd_sc_hd__nor2_1
XFILLER_0_73_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16767_ _02979_ _06494_ VGND VGND VPWR VPWR _07184_ sky130_fd_sc_hd__or2_1
X_13979_ _03005_ _00213_ VGND VGND VPWR VPWR _04151_ sky130_fd_sc_hd__nand2_1
X_18506_ _09044_ _09047_ _09073_ _06649_ VGND VGND VPWR VPWR _09074_ sky130_fd_sc_hd__o31a_1
X_15718_ _05972_ _05982_ _05980_ VGND VGND VPWR VPWR _06047_ sky130_fd_sc_hd__a21oi_1
X_16698_ _02533_ _07104_ _07105_ VGND VGND VPWR VPWR _07108_ sky130_fd_sc_hd__and3_2
X_18437_ _06374_ _03311_ VGND VGND VPWR VPWR _09000_ sky130_fd_sc_hd__nand2_1
X_15649_ _01359_ _03071_ _05900_ _05898_ VGND VGND VPWR VPWR _05972_ sky130_fd_sc_hd__a31o_1
XFILLER_0_118_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_145_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18368_ _03068_ _08428_ _02992_ VGND VGND VPWR VPWR _08926_ sky130_fd_sc_hd__or3b_1
XFILLER_0_71_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17319_ _07783_ _07784_ VGND VGND VPWR VPWR _07785_ sky130_fd_sc_hd__xor2_1
XFILLER_0_16_448 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_126_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18299_ _07314_ _08260_ _08777_ _04023_ VGND VGND VPWR VPWR _08851_ sky130_fd_sc_hd__or4b_1
XFILLER_0_71_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_144 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_141_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09506_ _04121_ VGND VGND VPWR VPWR _04132_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_67_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09437_ net172 VGND VGND VPWR VPWR _03377_ sky130_fd_sc_hd__buf_6
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_60 _04406_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_71 _05845_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11330_ cla_inst.in2\[21\] _00193_ _01349_ VGND VGND VPWR VPWR _01423_ sky130_fd_sc_hd__and3_1
XANTENNA_82 _07810_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_93 _08880_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11261_ _00163_ _00223_ VGND VGND VPWR VPWR _01354_ sky130_fd_sc_hd__nand2_2
X_10212_ _08529_ _08659_ _00303_ _00304_ VGND VGND VPWR VPWR _00305_ sky130_fd_sc_hd__o211a_1
X_13000_ _03040_ _03092_ VGND VGND VPWR VPWR _03093_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11192_ _01283_ _01280_ VGND VGND VPWR VPWR _01285_ sky130_fd_sc_hd__or2b_1
X_10143_ _00106_ _00194_ VGND VGND VPWR VPWR _00236_ sky130_fd_sc_hd__nand2_1
XFILLER_0_100_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14951_ _02984_ _01520_ _09256_ _00498_ VGND VGND VPWR VPWR _05212_ sky130_fd_sc_hd__and4_2
X_10074_ _00166_ VGND VGND VPWR VPWR _00167_ sky130_fd_sc_hd__buf_4
X_13902_ _04065_ _04066_ VGND VGND VPWR VPWR _04068_ sky130_fd_sc_hd__nand2_1
X_17670_ _08165_ _08166_ VGND VGND VPWR VPWR _08167_ sky130_fd_sc_hd__nor2_1
X_14882_ _05100_ _05013_ _05135_ VGND VGND VPWR VPWR _05138_ sky130_fd_sc_hd__nor3_1
X_16621_ _04132_ _03184_ _03313_ net150 VGND VGND VPWR VPWR _07024_ sky130_fd_sc_hd__a211oi_2
X_13833_ _07537_ _00247_ _03988_ _03991_ VGND VGND VPWR VPWR _03992_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_43_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16552_ _06945_ _06948_ VGND VGND VPWR VPWR _06950_ sky130_fd_sc_hd__nand2_1
XFILLER_0_69_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13764_ _03054_ _03058_ _03070_ _03075_ _03050_ _03061_ VGND VGND VPWR VPWR _03917_
+ sky130_fd_sc_hd__mux4_1
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10976_ _01040_ _01043_ VGND VGND VPWR VPWR _01069_ sky130_fd_sc_hd__nand2_1
XFILLER_0_85_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15503_ _03321_ _07384_ _08158_ _03322_ VGND VGND VPWR VPWR _05814_ sky130_fd_sc_hd__a22o_1
XFILLER_0_57_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_123 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12715_ _02783_ _02784_ _02807_ VGND VGND VPWR VPWR _02808_ sky130_fd_sc_hd__a21oi_1
X_16483_ _06874_ VGND VGND VPWR VPWR _06875_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_57_359 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13695_ _03839_ _03840_ VGND VGND VPWR VPWR _03841_ sky130_fd_sc_hd__or2_1
XFILLER_0_128_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18222_ _06776_ _08766_ _08767_ _06721_ VGND VGND VPWR VPWR _08769_ sky130_fd_sc_hd__o211a_1
X_15434_ _05737_ _05738_ VGND VGND VPWR VPWR _05739_ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_84_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12646_ _02733_ _02737_ _02738_ VGND VGND VPWR VPWR _02739_ sky130_fd_sc_hd__nand3_2
XFILLER_0_25_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18153_ _02969_ _08674_ _08693_ VGND VGND VPWR VPWR _08694_ sky130_fd_sc_hd__o21a_1
XFILLER_0_143_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15365_ _05662_ _05663_ VGND VGND VPWR VPWR _05664_ sky130_fd_sc_hd__nand2_1
XFILLER_0_25_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12577_ _02592_ _02631_ VGND VGND VPWR VPWR _02670_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_136_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_779 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17104_ _07432_ _07433_ _07550_ VGND VGND VPWR VPWR _07551_ sky130_fd_sc_hd__o21ai_1
X_14316_ _00107_ _04591_ VGND VGND VPWR VPWR _04520_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11528_ _01605_ _01606_ _01619_ _01620_ VGND VGND VPWR VPWR _01621_ sky130_fd_sc_hd__a211oi_4
X_18084_ _08541_ _08542_ _08543_ _08537_ VGND VGND VPWR VPWR _08618_ sky130_fd_sc_hd__or4b_1
X_15296_ _05575_ _05576_ _05587_ VGND VGND VPWR VPWR _05589_ sky130_fd_sc_hd__nand3_1
XFILLER_0_150_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17035_ _02973_ _07475_ VGND VGND VPWR VPWR _07476_ sky130_fd_sc_hd__nor2_1
X_14247_ _04275_ _04281_ _04273_ VGND VGND VPWR VPWR _04444_ sky130_fd_sc_hd__a21o_1
X_11459_ _03717_ _00177_ VGND VGND VPWR VPWR _01552_ sky130_fd_sc_hd__and2_1
XFILLER_0_110_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14178_ _04158_ _04368_ VGND VGND VPWR VPWR _04369_ sky130_fd_sc_hd__or2_1
XTAP_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13129_ _03221_ _03222_ _03223_ VGND VGND VPWR VPWR _03225_ sky130_fd_sc_hd__a21oi_2
XTAP_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18986_ clknet_4_1_0_clk _09382_ VGND VGND VPWR VPWR salida\[39\] sky130_fd_sc_hd__dfxtp_1
XTAP_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17937_ _08456_ _08457_ VGND VGND VPWR VPWR _08458_ sky130_fd_sc_hd__xor2_1
XFILLER_0_84_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17868_ _07303_ _07621_ VGND VGND VPWR VPWR _08383_ sky130_fd_sc_hd__nor2_1
XFILLER_0_108_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16819_ _07231_ _07239_ VGND VGND VPWR VPWR _07240_ sky130_fd_sc_hd__xor2_1
X_17799_ _07038_ _07859_ _08306_ VGND VGND VPWR VPWR _08308_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_76_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_624 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_495 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_715 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_668 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_146_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09986_ _07700_ _07733_ _07766_ VGND VGND VPWR VPWR _09279_ sky130_fd_sc_hd__and3_1
XFILLER_0_110_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwb_buttons_leds_156 VGND VGND VPWR VPWR wb_buttons_leds_156/HI led_enb[5] sky130_fd_sc_hd__conb_1
X_10830_ _03717_ _03476_ VGND VGND VPWR VPWR _00923_ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10761_ _00824_ _00852_ _00853_ VGND VGND VPWR VPWR _00854_ sky130_fd_sc_hd__and3_2
XFILLER_0_82_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12500_ _02576_ _02577_ VGND VGND VPWR VPWR _02593_ sky130_fd_sc_hd__xnor2_1
X_13480_ _03383_ _03389_ _03382_ VGND VGND VPWR VPWR _03605_ sky130_fd_sc_hd__a21bo_1
X_10692_ _00783_ _00784_ VGND VGND VPWR VPWR _00785_ sky130_fd_sc_hd__or2_1
X_12431_ _02439_ _02518_ VGND VGND VPWR VPWR _02524_ sky130_fd_sc_hd__nand2_1
XFILLER_0_125_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_118_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_124_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15150_ _05345_ _05346_ VGND VGND VPWR VPWR _05429_ sky130_fd_sc_hd__nor2_1
XFILLER_0_62_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12362_ net128 _02449_ _02416_ _02448_ VGND VGND VPWR VPWR _02455_ sky130_fd_sc_hd__o211a_1
X_14101_ _04267_ _04268_ _04282_ VGND VGND VPWR VPWR _04284_ sky130_fd_sc_hd__nor3_1
XFILLER_0_105_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11313_ _01396_ _01404_ _01397_ _01398_ VGND VGND VPWR VPWR _01406_ sky130_fd_sc_hd__nor4_1
X_15081_ _05352_ _05353_ _00106_ _00309_ VGND VGND VPWR VPWR _05354_ sky130_fd_sc_hd__and4bb_1
X_12293_ _02378_ _02380_ VGND VGND VPWR VPWR _02386_ sky130_fd_sc_hd__nor2_1
XFILLER_0_132_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14032_ _04208_ VGND VGND VPWR VPWR _04210_ sky130_fd_sc_hd__inv_2
X_11244_ _01079_ _01147_ _01335_ _01336_ VGND VGND VPWR VPWR _01337_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_31_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_120_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11175_ _01141_ _01266_ VGND VGND VPWR VPWR _01268_ sky130_fd_sc_hd__and2_1
X_18840_ clknet_4_1_0_clk net312 VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__dfxtp_1
X_10126_ _00175_ _00218_ _00178_ _00173_ VGND VGND VPWR VPWR _00219_ sky130_fd_sc_hd__a22oi_1
X_18771_ _02200_ net40 _09276_ VGND VGND VPWR VPWR _09286_ sky130_fd_sc_hd__mux2_1
X_15983_ _02347_ _00558_ VGND VGND VPWR VPWR _06331_ sky130_fd_sc_hd__or2_1
X_17722_ _06516_ _08222_ _08223_ VGND VGND VPWR VPWR _08225_ sky130_fd_sc_hd__and3_1
X_10057_ _00148_ _00149_ _00131_ _00127_ VGND VGND VPWR VPWR _00150_ sky130_fd_sc_hd__nand4_2
X_14934_ _05069_ _05071_ VGND VGND VPWR VPWR _05195_ sky130_fd_sc_hd__and2_1
XFILLER_0_89_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17653_ _08065_ _08078_ VGND VGND VPWR VPWR _08149_ sky130_fd_sc_hd__nor2_1
X_14865_ _04986_ _04990_ _05118_ VGND VGND VPWR VPWR _05119_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_86_900 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16604_ _02728_ _06592_ _06551_ VGND VGND VPWR VPWR _07007_ sky130_fd_sc_hd__a21o_1
X_13816_ _05224_ _09256_ VGND VGND VPWR VPWR _03973_ sky130_fd_sc_hd__nand2_1
XFILLER_0_58_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17584_ _08067_ _07947_ _08073_ VGND VGND VPWR VPWR _08074_ sky130_fd_sc_hd__o21a_1
X_14796_ _04887_ _04888_ _04889_ VGND VGND VPWR VPWR _05044_ sky130_fd_sc_hd__o21ba_1
X_16535_ _06836_ _06911_ _06912_ _06931_ VGND VGND VPWR VPWR _06932_ sky130_fd_sc_hd__o31a_1
X_13747_ _03687_ _03688_ _03691_ VGND VGND VPWR VPWR _03898_ sky130_fd_sc_hd__and3_1
X_10959_ _00941_ _00954_ _00953_ VGND VGND VPWR VPWR _01052_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_70_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16466_ _06349_ _06348_ _06338_ VGND VGND VPWR VPWR _06857_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_6_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13678_ _07526_ _00165_ _03819_ _03821_ VGND VGND VPWR VPWR _03822_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_45_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18205_ _08748_ _08749_ VGND VGND VPWR VPWR _08750_ sky130_fd_sc_hd__and2b_1
X_15417_ _05449_ _01112_ _05678_ _05680_ VGND VGND VPWR VPWR _05720_ sky130_fd_sc_hd__a31o_1
X_12629_ _02686_ _02721_ VGND VGND VPWR VPWR _02722_ sky130_fd_sc_hd__and2_1
X_16397_ _06674_ _06675_ _06672_ VGND VGND VPWR VPWR _06782_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_115_228 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18136_ _02997_ _06512_ _03052_ VGND VGND VPWR VPWR _08675_ sky130_fd_sc_hd__a21boi_1
X_15348_ _05563_ _05630_ _05643_ VGND VGND VPWR VPWR _05645_ sky130_fd_sc_hd__nor3_1
XFILLER_0_85_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_112_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_250 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18067_ _04647_ _06445_ VGND VGND VPWR VPWR _08600_ sky130_fd_sc_hd__or2_1
Xhold105 _00031_ VGND VGND VPWR VPWR net268 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15279_ _05567_ _05569_ VGND VGND VPWR VPWR _05570_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_79_78 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold116 net95 VGND VGND VPWR VPWR net279 sky130_fd_sc_hd__dlygate4sd3_1
Xhold127 _00020_ VGND VGND VPWR VPWR net290 sky130_fd_sc_hd__dlygate4sd3_1
Xhold138 net94 VGND VGND VPWR VPWR net301 sky130_fd_sc_hd__dlygate4sd3_1
Xhold149 _00006_ VGND VGND VPWR VPWR net312 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17018_ _07455_ _07456_ VGND VGND VPWR VPWR _07457_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09840_ ApproximateM_inst.lob_16.lob2.mux.sel _07755_ VGND VGND VPWR VPWR _07766_
+ sky130_fd_sc_hd__and2_4
XTAP_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09771_ _07004_ VGND VGND VPWR VPWR _07015_ sky130_fd_sc_hd__buf_4
XTAP_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18969_ clknet_4_5_0_clk _09400_ VGND VGND VPWR VPWR salida\[22\] sky130_fd_sc_hd__dfxtp_1
XTAP_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_386 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_151_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_395 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_130_743 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09969_ _09037_ _09048_ _09145_ VGND VGND VPWR VPWR _09152_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_99_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12980_ _03072_ VGND VGND VPWR VPWR _03073_ sky130_fd_sc_hd__buf_4
X_11931_ _02023_ VGND VGND VPWR VPWR _02024_ sky130_fd_sc_hd__inv_2
XTAP_2800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14650_ _04603_ _04752_ VGND VGND VPWR VPWR _04884_ sky130_fd_sc_hd__and2b_1
X_11862_ _01847_ _01846_ VGND VGND VPWR VPWR _01955_ sky130_fd_sc_hd__and2b_1
XFILLER_0_86_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13601_ _03736_ _03737_ VGND VGND VPWR VPWR _03738_ sky130_fd_sc_hd__or2_1
X_10813_ _00761_ _00905_ VGND VGND VPWR VPWR _00906_ sky130_fd_sc_hd__nor2_1
X_14581_ _04807_ _04808_ VGND VGND VPWR VPWR _04809_ sky130_fd_sc_hd__xor2_2
XFILLER_0_83_903 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11793_ _01601_ _01602_ _01603_ _01564_ VGND VGND VPWR VPWR _01886_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_55_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16320_ _03061_ _06696_ _06697_ VGND VGND VPWR VPWR _06698_ sky130_fd_sc_hd__a21bo_1
X_13532_ _03453_ _03457_ VGND VGND VPWR VPWR _03663_ sky130_fd_sc_hd__or2b_1
X_10744_ _07352_ _06722_ _07951_ _07995_ VGND VGND VPWR VPWR _00837_ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16251_ _03026_ _03041_ _01696_ VGND VGND VPWR VPWR _06623_ sky130_fd_sc_hd__a21o_1
X_13463_ _03393_ _03394_ _03405_ VGND VGND VPWR VPWR _03587_ sky130_fd_sc_hd__nor3_1
XFILLER_0_36_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10675_ _00766_ _00767_ VGND VGND VPWR VPWR _00768_ sky130_fd_sc_hd__xor2_2
XFILLER_0_152_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15202_ _01505_ _00322_ _05371_ VGND VGND VPWR VPWR _05487_ sky130_fd_sc_hd__and3_1
XFILLER_0_153_868 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12414_ _02503_ _02504_ _02506_ VGND VGND VPWR VPWR _02507_ sky130_fd_sc_hd__and3_1
X_16182_ _03200_ _06547_ _06477_ VGND VGND VPWR VPWR _06549_ sky130_fd_sc_hd__o21a_1
X_13394_ _03471_ _03472_ _03510_ _03511_ VGND VGND VPWR VPWR _03512_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_50_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15133_ _05196_ _05299_ _05300_ VGND VGND VPWR VPWR _05412_ sky130_fd_sc_hd__o21ba_1
X_12345_ _00846_ _00248_ _02370_ VGND VGND VPWR VPWR _02438_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_133_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_105_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15064_ _05334_ VGND VGND VPWR VPWR _05336_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12276_ _02353_ _02367_ VGND VGND VPWR VPWR _02369_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_120_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_120_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14015_ _04189_ _04190_ VGND VGND VPWR VPWR _04191_ sky130_fd_sc_hd__xor2_4
X_11227_ _05050_ _01009_ _01008_ _01011_ VGND VGND VPWR VPWR _01320_ sky130_fd_sc_hd__o2bb2a_1
X_18823_ _09327_ VGND VGND VPWR VPWR _00098_ sky130_fd_sc_hd__buf_1
X_11158_ _01226_ _01250_ VGND VGND VPWR VPWR _01251_ sky130_fd_sc_hd__and2_1
X_10109_ _00188_ _00201_ VGND VGND VPWR VPWR _00202_ sky130_fd_sc_hd__and2b_1
X_11089_ _08713_ _00715_ _01054_ _01055_ VGND VGND VPWR VPWR _01182_ sky130_fd_sc_hd__a22o_2
X_18754_ _09125_ VGND VGND VPWR VPWR _09273_ sky130_fd_sc_hd__buf_2
X_15966_ _06299_ _06301_ _06312_ VGND VGND VPWR VPWR _06314_ sky130_fd_sc_hd__a21o_1
XFILLER_0_65_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17705_ _08203_ _08205_ VGND VGND VPWR VPWR _08206_ sky130_fd_sc_hd__and2_1
X_14917_ _00591_ _03142_ _05175_ VGND VGND VPWR VPWR _05176_ sky130_fd_sc_hd__nand3_1
X_18685_ net43 _03111_ _09193_ VGND VGND VPWR VPWR _09221_ sky130_fd_sc_hd__mux2_1
X_15897_ _06194_ _06195_ _06197_ _06239_ VGND VGND VPWR VPWR _06240_ sky130_fd_sc_hd__a31oi_2
X_14848_ _04862_ _04969_ _04997_ _04998_ VGND VGND VPWR VPWR _05100_ sky130_fd_sc_hd__o211a_1
X_17636_ _08130_ VGND VGND VPWR VPWR _08131_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17567_ _06961_ _07487_ _07593_ _07018_ VGND VGND VPWR VPWR _08055_ sky130_fd_sc_hd__o22a_1
XFILLER_0_147_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14779_ _05019_ _05023_ _05024_ VGND VGND VPWR VPWR _05025_ sky130_fd_sc_hd__and3_1
XFILLER_0_81_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16518_ _02981_ _06611_ VGND VGND VPWR VPWR _06913_ sky130_fd_sc_hd__or2_2
XFILLER_0_14_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17498_ _07302_ _07115_ _07218_ _07313_ VGND VGND VPWR VPWR _07980_ sky130_fd_sc_hd__or4_1
XFILLER_0_144_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16449_ _03535_ _06673_ _01264_ VGND VGND VPWR VPWR _06838_ sky130_fd_sc_hd__o21a_1
XFILLER_0_6_735 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_143_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18119_ _08488_ _08556_ _08559_ VGND VGND VPWR VPWR _08656_ sky130_fd_sc_hd__and3_1
XFILLER_0_41_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09823_ ApproximateM_inst.lob_16.lob1.mux.sel VGND VGND VPWR VPWR _07581_ sky130_fd_sc_hd__clkbuf_4
X_09754_ _06558_ _06569_ _06808_ VGND VGND VPWR VPWR _06830_ sky130_fd_sc_hd__nand3_1
X_09685_ _05649_ VGND VGND VPWR VPWR _06084_ sky130_fd_sc_hd__buf_4
XTAP_2107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_744 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_147_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_119_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10460_ _00543_ _00552_ VGND VGND VPWR VPWR _00553_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_150_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10391_ _00314_ _00315_ VGND VGND VPWR VPWR _00484_ sky130_fd_sc_hd__and2_1
XFILLER_0_33_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12130_ _02187_ _02222_ VGND VGND VPWR VPWR _02223_ sky130_fd_sc_hd__nand2_1
XFILLER_0_102_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_798 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12061_ _02148_ _02152_ _02070_ _02153_ VGND VGND VPWR VPWR _02154_ sky130_fd_sc_hd__o211a_1
XFILLER_0_3_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11012_ ApproximateM_inst.lob_16.lob2.genblk1\[1\].genblk1.mux.sel VGND VGND VPWR
+ VPWR _01105_ sky130_fd_sc_hd__inv_2
X_15820_ _03016_ _03154_ _06154_ _06156_ VGND VGND VPWR VPWR _06157_ sky130_fd_sc_hd__and4_1
X_15751_ _04256_ _04261_ _03537_ VGND VGND VPWR VPWR _06083_ sky130_fd_sc_hd__mux2_1
X_12963_ _03055_ VGND VGND VPWR VPWR _03056_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_87_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_99_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14702_ _04939_ _04940_ VGND VGND VPWR VPWR _04942_ sky130_fd_sc_hd__or2_4
X_11914_ _02001_ _02004_ _02006_ VGND VGND VPWR VPWR _02007_ sky130_fd_sc_hd__o21ai_1
X_18470_ _03073_ _06464_ _09017_ _09035_ VGND VGND VPWR VPWR _09407_ sky130_fd_sc_hd__o2bb2a_1
X_15682_ _06006_ _06007_ VGND VGND VPWR VPWR _06009_ sky130_fd_sc_hd__or2_1
XTAP_2630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12894_ _02986_ VGND VGND VPWR VPWR _02987_ sky130_fd_sc_hd__buf_4
XTAP_2641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17421_ _07893_ _07895_ VGND VGND VPWR VPWR _07896_ sky130_fd_sc_hd__xor2_1
XTAP_2652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14633_ _04862_ _04863_ _04730_ _04833_ VGND VGND VPWR VPWR _04866_ sky130_fd_sc_hd__o211ai_4
XTAP_2663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11845_ net341 _01932_ _01936_ _01937_ VGND VGND VPWR VPWR _01938_ sky130_fd_sc_hd__o211a_1
XTAP_2674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17352_ _07783_ _07784_ VGND VGND VPWR VPWR _07821_ sky130_fd_sc_hd__and2b_1
XFILLER_0_28_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14564_ _04778_ _04779_ _04790_ VGND VGND VPWR VPWR _04791_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_55_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11776_ _01861_ _01865_ _01867_ _01868_ VGND VGND VPWR VPWR _01869_ sky130_fd_sc_hd__or4_4
XTAP_1984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16303_ _06461_ VGND VGND VPWR VPWR _06680_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_126_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13515_ _03422_ _03424_ _03642_ _03643_ VGND VGND VPWR VPWR _03644_ sky130_fd_sc_hd__a211oi_4
X_10727_ _00795_ _00796_ _00779_ _00794_ VGND VGND VPWR VPWR _00820_ sky130_fd_sc_hd__o211a_1
X_17283_ _07038_ _07665_ _07745_ _06527_ VGND VGND VPWR VPWR _07746_ sky130_fd_sc_hd__a22o_1
X_14495_ _03859_ _03793_ cla_inst.in1\[28\] _07374_ VGND VGND VPWR VPWR _04715_ sky130_fd_sc_hd__and4_1
XFILLER_0_43_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16234_ _03161_ _03029_ _02805_ VGND VGND VPWR VPWR _06605_ sky130_fd_sc_hd__a21o_1
XFILLER_0_152_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13446_ _03145_ _03151_ _03089_ VGND VGND VPWR VPWR _03568_ sky130_fd_sc_hd__mux2_1
X_10658_ _00747_ _00748_ _00749_ VGND VGND VPWR VPWR _00751_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_152_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_125_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16165_ ApproximateM_inst.lob_16.lob1.genblk1\[12\].genblk1.mux.sel net208 ApproximateM_inst.lob_16.lob1.genblk1\[10\].genblk1.mux.sel
+ ApproximateM_inst.lob_16.lob1.genblk1\[9\].genblk1.mux.sel VGND VGND VPWR VPWR _06530_
+ sky130_fd_sc_hd__or4_4
X_13377_ _03320_ _03328_ VGND VGND VPWR VPWR _03493_ sky130_fd_sc_hd__and2b_1
XFILLER_0_11_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10589_ _00680_ _00681_ _07537_ _00194_ VGND VGND VPWR VPWR _00682_ sky130_fd_sc_hd__and4bb_1
X_15116_ _05240_ _05242_ VGND VGND VPWR VPWR _05393_ sky130_fd_sc_hd__and2b_1
X_12328_ _02419_ _02420_ _00832_ _03618_ VGND VGND VPWR VPWR _02421_ sky130_fd_sc_hd__and4bb_1
X_16096_ _05419_ _05422_ _02974_ VGND VGND VPWR VPWR _06455_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15047_ _05315_ _05316_ VGND VGND VPWR VPWR _05317_ sky130_fd_sc_hd__nor2_1
X_12259_ _02228_ _02350_ _02351_ VGND VGND VPWR VPWR _02352_ sky130_fd_sc_hd__and3_1
X_18806_ _01359_ net52 _09301_ VGND VGND VPWR VPWR _09314_ sky130_fd_sc_hd__mux2_1
X_16998_ _07324_ _07326_ VGND VGND VPWR VPWR _07435_ sky130_fd_sc_hd__nor2_1
X_18737_ _09245_ _09259_ VGND VGND VPWR VPWR _09260_ sky130_fd_sc_hd__and2_1
X_15949_ _03121_ _06295_ VGND VGND VPWR VPWR _06296_ sky130_fd_sc_hd__nand2_1
X_09470_ ApproximateM_inst.lob_16.lob1.genblk1\[13\].genblk1.mux.sel VGND VGND VPWR
+ VPWR _03739_ sky130_fd_sc_hd__buf_6
X_18668_ _09125_ VGND VGND VPWR VPWR _09209_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_25_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17619_ _07999_ _08007_ _07997_ VGND VGND VPWR VPWR _08112_ sky130_fd_sc_hd__a21o_1
X_18599_ salida\[19\] _09141_ _09142_ salida\[51\] _09146_ VGND VGND VPWR VPWR _09156_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_58_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_571 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_144_676 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_332 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_104_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_112_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09806_ _07363_ _07384_ VGND VGND VPWR VPWR _07395_ sky130_fd_sc_hd__nand2_1
X_09737_ _06580_ _06635_ VGND VGND VPWR VPWR _06646_ sky130_fd_sc_hd__xnor2_1
X_09668_ _05366_ _05497_ _04580_ _05410_ VGND VGND VPWR VPWR _05899_ sky130_fd_sc_hd__a22o_1
XTAP_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09599_ _04941_ _04952_ _04962_ VGND VGND VPWR VPWR _05148_ sky130_fd_sc_hd__a21o_1
XTAP_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11630_ _01215_ _01214_ _01209_ VGND VGND VPWR VPWR _01723_ sky130_fd_sc_hd__a21o_1
XTAP_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11561_ _01652_ _01653_ VGND VGND VPWR VPWR _01654_ sky130_fd_sc_hd__and2b_1
XFILLER_0_108_835 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13300_ _03224_ net135 _03406_ _03407_ VGND VGND VPWR VPWR _03408_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_107_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10512_ _03651_ _03662_ _04580_ _04482_ VGND VGND VPWR VPWR _00605_ sky130_fd_sc_hd__nand4_2
XFILLER_0_52_427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_736 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_134_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14280_ _04474_ _04477_ _04479_ VGND VGND VPWR VPWR _04480_ sky130_fd_sc_hd__or3_2
X_11492_ _01581_ _01583_ _01584_ VGND VGND VPWR VPWR _01585_ sky130_fd_sc_hd__nand3_4
XFILLER_0_80_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13231_ _03315_ _00735_ _03332_ VGND VGND VPWR VPWR _03334_ sky130_fd_sc_hd__and3_1
XFILLER_0_122_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10443_ _00532_ _00533_ _00534_ _00491_ VGND VGND VPWR VPWR _00536_ sky130_fd_sc_hd__a22o_1
X_13162_ _00651_ _00653_ _03258_ _03259_ VGND VGND VPWR VPWR _03261_ sky130_fd_sc_hd__a211o_1
X_10374_ _00291_ _00431_ _00465_ _00466_ VGND VGND VPWR VPWR _00467_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_103_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12113_ _00127_ _02205_ VGND VGND VPWR VPWR _02206_ sky130_fd_sc_hd__nand2_1
X_13093_ _02505_ _01862_ VGND VGND VPWR VPWR _03186_ sky130_fd_sc_hd__nor2_1
X_17970_ _08391_ _08493_ VGND VGND VPWR VPWR _08494_ sky130_fd_sc_hd__xor2_1
X_12044_ _02073_ _02076_ _02075_ VGND VGND VPWR VPWR _02137_ sky130_fd_sc_hd__o21ai_1
X_16921_ _07349_ _07350_ VGND VGND VPWR VPWR _07351_ sky130_fd_sc_hd__nor2_2
X_16852_ _06357_ _07274_ _07275_ _00167_ VGND VGND VPWR VPWR _07277_ sky130_fd_sc_hd__a2bb2o_1
X_15803_ _06137_ _06139_ VGND VGND VPWR VPWR _06140_ sky130_fd_sc_hd__or2_1
X_16783_ _06937_ _07143_ _07198_ VGND VGND VPWR VPWR _07201_ sky130_fd_sc_hd__o21ai_1
X_13995_ _04166_ _04167_ _04168_ VGND VGND VPWR VPWR _04169_ sky130_fd_sc_hd__and3_4
XFILLER_0_99_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15734_ _06023_ _06064_ VGND VGND VPWR VPWR _06065_ sky130_fd_sc_hd__nor2_1
X_18522_ _02949_ _02956_ _09061_ VGND VGND VPWR VPWR _09092_ sky130_fd_sc_hd__or3_1
XFILLER_0_99_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12946_ _03038_ VGND VGND VPWR VPWR _03039_ sky130_fd_sc_hd__clkbuf_4
X_15665_ _05970_ _05971_ _05988_ VGND VGND VPWR VPWR _05990_ sky130_fd_sc_hd__or3_1
X_18453_ _03013_ _06512_ _03073_ VGND VGND VPWR VPWR _09018_ sky130_fd_sc_hd__a21boi_1
X_12877_ _00759_ _02964_ _02969_ VGND VGND VPWR VPWR _02970_ sky130_fd_sc_hd__a21oi_1
XANTENNA_150 _08762_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_161 _08762_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17404_ _07854_ _07877_ VGND VGND VPWR VPWR _07878_ sky130_fd_sc_hd__nor2_1
X_14616_ _04001_ _00502_ VGND VGND VPWR VPWR _04847_ sky130_fd_sc_hd__nand2_1
XANTENNA_172 _02646_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18384_ _04238_ _08934_ _08943_ VGND VGND VPWR VPWR _08944_ sky130_fd_sc_hd__o21ai_1
X_11828_ _01831_ _01830_ _01829_ VGND VGND VPWR VPWR _01921_ sky130_fd_sc_hd__a21oi_1
X_15596_ _05838_ _05839_ VGND VGND VPWR VPWR _05915_ sky130_fd_sc_hd__nand2_1
XTAP_1770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17335_ _07681_ _07682_ _07680_ VGND VGND VPWR VPWR _07803_ sky130_fd_sc_hd__a21bo_1
X_14547_ _04639_ _04641_ _04770_ VGND VGND VPWR VPWR _04772_ sky130_fd_sc_hd__nor3_1
X_11759_ _01849_ _01851_ VGND VGND VPWR VPWR _01852_ sky130_fd_sc_hd__or2_4
XFILLER_0_43_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17266_ _07720_ _07726_ VGND VGND VPWR VPWR _07727_ sky130_fd_sc_hd__xor2_1
X_14478_ _04695_ _04696_ VGND VGND VPWR VPWR _04697_ sky130_fd_sc_hd__nor2_1
XFILLER_0_153_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16217_ _01106_ _06585_ _07646_ VGND VGND VPWR VPWR _06586_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_113_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19005_ clknet_4_7_0_clk _09372_ VGND VGND VPWR VPWR salida\[58\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13429_ _03096_ _03103_ _03047_ VGND VGND VPWR VPWR _03550_ sky130_fd_sc_hd__mux2_1
X_17197_ _07651_ VGND VGND VPWR VPWR _07652_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_140_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16148_ _06510_ VGND VGND VPWR VPWR _06511_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_12_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_122_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16079_ _00167_ _00214_ _06435_ VGND VGND VPWR VPWR _06436_ sky130_fd_sc_hd__and3_1
XFILLER_0_11_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput1 buttons VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__buf_4
X_09522_ _04187_ _04285_ _04296_ VGND VGND VPWR VPWR _04307_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_79_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09453_ _03443_ _03487_ _03542_ VGND VGND VPWR VPWR _03553_ sky130_fd_sc_hd__nand3_1
XPHY_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_117_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10090_ _00174_ VGND VGND VPWR VPWR _00183_ sky130_fd_sc_hd__buf_2
XFILLER_0_100_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12800_ _02869_ _02880_ _02879_ VGND VGND VPWR VPWR _02893_ sky130_fd_sc_hd__a21o_1
X_13780_ _03531_ _03509_ _08746_ _08049_ VGND VGND VPWR VPWR _03933_ sky130_fd_sc_hd__nand4_2
X_10992_ _07058_ _07091_ _00460_ _05856_ _01084_ VGND VGND VPWR VPWR _01085_ sky130_fd_sc_hd__a41o_1
XFILLER_0_69_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12731_ _02814_ _02817_ VGND VGND VPWR VPWR _02824_ sky130_fd_sc_hd__and2_1
XTAP_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15450_ _05739_ _05754_ VGND VGND VPWR VPWR _05756_ sky130_fd_sc_hd__nor2_1
XFILLER_0_32_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12662_ _07788_ _00120_ _00132_ _09219_ VGND VGND VPWR VPWR _02755_ sky130_fd_sc_hd__and4_1
XTAP_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14401_ _03005_ _00399_ VGND VGND VPWR VPWR _04612_ sky130_fd_sc_hd__nand2_1
XTAP_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11613_ _01640_ _01641_ _01564_ _01604_ VGND VGND VPWR VPWR _01706_ sky130_fd_sc_hd__o211a_1
XFILLER_0_139_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15381_ _05679_ _05680_ VGND VGND VPWR VPWR _05681_ sky130_fd_sc_hd__nor2_1
XFILLER_0_38_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12593_ ApproximateM_inst.lob_16.lob2.genblk1\[1\].genblk1.mux.sel _00180_ _02685_
+ VGND VGND VPWR VPWR _02686_ sky130_fd_sc_hd__and3_1
XFILLER_0_92_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17120_ _07565_ _07566_ _07567_ VGND VGND VPWR VPWR _07568_ sky130_fd_sc_hd__nand3_1
X_14332_ _04489_ _04490_ _04535_ _04536_ VGND VGND VPWR VPWR _04538_ sky130_fd_sc_hd__and4_2
X_11544_ _01633_ _01634_ _01635_ VGND VGND VPWR VPWR _01637_ sky130_fd_sc_hd__a21o_1
XFILLER_0_80_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17051_ _07485_ _07491_ VGND VGND VPWR VPWR _07492_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_150_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14263_ _04283_ _04429_ _04459_ VGND VGND VPWR VPWR _04462_ sky130_fd_sc_hd__or3_2
XFILLER_0_123_635 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11475_ _01565_ _01566_ _01567_ VGND VGND VPWR VPWR _01568_ sky130_fd_sc_hd__nand3_1
XFILLER_0_40_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16002_ _07058_ _00193_ _06346_ _02358_ _02215_ VGND VGND VPWR VPWR _06352_ sky130_fd_sc_hd__a311o_1
XFILLER_0_122_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13214_ _00725_ _00730_ VGND VGND VPWR VPWR _03316_ sky130_fd_sc_hd__and2_1
XFILLER_0_122_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10426_ _00512_ _00518_ VGND VGND VPWR VPWR _00519_ sky130_fd_sc_hd__xor2_1
XFILLER_0_104_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14194_ _04169_ net120 _04385_ _04386_ VGND VGND VPWR VPWR _04387_ sky130_fd_sc_hd__o211a_4
XFILLER_0_104_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13145_ _06029_ _06051_ _07384_ VGND VGND VPWR VPWR _03243_ sky130_fd_sc_hd__and3_1
XFILLER_0_103_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10357_ _00447_ _00448_ _00449_ VGND VGND VPWR VPWR _00450_ sky130_fd_sc_hd__and3_2
XTAP_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13076_ _03023_ _03167_ VGND VGND VPWR VPWR _03168_ sky130_fd_sc_hd__nand2_1
X_17953_ _07106_ _07621_ _08472_ _08473_ VGND VGND VPWR VPWR _08476_ sky130_fd_sc_hd__o22a_1
X_10288_ _00233_ _00243_ VGND VGND VPWR VPWR _00381_ sky130_fd_sc_hd__or2_1
X_12027_ _02115_ net187 VGND VGND VPWR VPWR _02120_ sky130_fd_sc_hd__and2b_1
X_16904_ _07224_ _07226_ VGND VGND VPWR VPWR _07333_ sky130_fd_sc_hd__nand2_1
X_17884_ _08380_ _08399_ VGND VGND VPWR VPWR _08401_ sky130_fd_sc_hd__nor2_1
X_16835_ _02476_ _02099_ _06510_ VGND VGND VPWR VPWR _07258_ sky130_fd_sc_hd__and3_1
X_13978_ _03965_ _03978_ VGND VGND VPWR VPWR _04150_ sky130_fd_sc_hd__and2b_1
XFILLER_0_87_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16766_ _03912_ _06474_ VGND VGND VPWR VPWR _07183_ sky130_fd_sc_hd__nor2_1
XFILLER_0_87_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18505_ _03108_ _08150_ _09072_ _09042_ _09041_ VGND VGND VPWR VPWR _09073_ sky130_fd_sc_hd__a32o_1
X_15717_ _05966_ _06045_ VGND VGND VPWR VPWR _06046_ sky130_fd_sc_hd__xnor2_1
X_12929_ _03002_ _03021_ VGND VGND VPWR VPWR _03022_ sky130_fd_sc_hd__nor2_2
X_16697_ _06563_ _06937_ _06961_ _07106_ VGND VGND VPWR VPWR _07107_ sky130_fd_sc_hd__or4_1
XFILLER_0_87_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18436_ _08950_ _08952_ _08949_ VGND VGND VPWR VPWR _08999_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_8_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15648_ _05909_ _05908_ VGND VGND VPWR VPWR _05971_ sky130_fd_sc_hd__and2b_1
XTAP_2290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15579_ _00112_ _07384_ VGND VGND VPWR VPWR _05896_ sky130_fd_sc_hd__and2_1
X_18367_ _02992_ _06512_ _03068_ VGND VGND VPWR VPWR _08925_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_84_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_75 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_145_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17318_ _07647_ _07660_ _07645_ VGND VGND VPWR VPWR _07784_ sky130_fd_sc_hd__a21o_1
XFILLER_0_28_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18298_ _02200_ _07780_ _08150_ _07650_ VGND VGND VPWR VPWR _08850_ sky130_fd_sc_hd__a22o_1
XFILLER_0_154_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_114_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17249_ _02059_ _07592_ VGND VGND VPWR VPWR _07708_ sky130_fd_sc_hd__and2_2
XFILLER_0_12_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09505_ _03771_ VGND VGND VPWR VPWR _04121_ sky130_fd_sc_hd__buf_6
XFILLER_0_94_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09436_ cla_inst.in2\[17\] VGND VGND VPWR VPWR _03366_ sky130_fd_sc_hd__buf_8
XFILLER_0_94_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_658 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_50 _03432_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_61 _04406_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_72 _06326_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_83 _08345_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_94 _08880_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_443 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11260_ _01351_ _01352_ VGND VGND VPWR VPWR _01353_ sky130_fd_sc_hd__nor2_2
X_10211_ _00291_ _00302_ _00301_ VGND VGND VPWR VPWR _00304_ sky130_fd_sc_hd__o21ai_1
X_11191_ _01280_ _01283_ VGND VGND VPWR VPWR _01284_ sky130_fd_sc_hd__or2b_1
X_10142_ _00150_ _00153_ VGND VGND VPWR VPWR _00235_ sky130_fd_sc_hd__nand2_1
X_10073_ _00165_ VGND VGND VPWR VPWR _00166_ sky130_fd_sc_hd__buf_8
X_14950_ _01520_ _00502_ _07733_ _02984_ VGND VGND VPWR VPWR _05211_ sky130_fd_sc_hd__a22oi_4
X_13901_ _04062_ _04064_ VGND VGND VPWR VPWR _04066_ sky130_fd_sc_hd__nand2_1
X_14881_ _05100_ _05013_ _05135_ VGND VGND VPWR VPWR _05136_ sky130_fd_sc_hd__o21a_1
X_13832_ _03987_ VGND VGND VPWR VPWR _03991_ sky130_fd_sc_hd__inv_2
X_16620_ _06812_ _03003_ net211 VGND VGND VPWR VPWR _07023_ sky130_fd_sc_hd__nor3_1
XFILLER_0_69_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16551_ _06571_ _06874_ _06947_ _06542_ VGND VGND VPWR VPWR _06948_ sky130_fd_sc_hd__a2bb2o_1
X_13763_ _03913_ VGND VGND VPWR VPWR _03916_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_57_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10975_ _01062_ _01067_ VGND VGND VPWR VPWR _01068_ sky130_fd_sc_hd__and2_1
XFILLER_0_85_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15502_ _03014_ _01317_ _05762_ _05761_ VGND VGND VPWR VPWR _05813_ sky130_fd_sc_hd__a31o_1
X_12714_ _02785_ _02806_ VGND VGND VPWR VPWR _02807_ sky130_fd_sc_hd__and2_1
X_16482_ _06869_ _06872_ _05736_ VGND VGND VPWR VPWR _06874_ sky130_fd_sc_hd__a21bo_2
X_13694_ cla_inst.in2\[24\] _00174_ _04471_ _03739_ VGND VGND VPWR VPWR _03840_ sky130_fd_sc_hd__and4_1
XFILLER_0_84_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15433_ _05719_ _05644_ _05735_ VGND VGND VPWR VPWR _05738_ sky130_fd_sc_hd__nor3_1
X_18221_ _06399_ _06546_ VGND VGND VPWR VPWR _08767_ sky130_fd_sc_hd__nand2_1
XFILLER_0_128_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12645_ _02700_ _02732_ _02731_ VGND VGND VPWR VPWR _02738_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_150_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15364_ _02999_ _03153_ _05661_ VGND VGND VPWR VPWR _05663_ sky130_fd_sc_hd__a21o_1
X_18152_ _06836_ _08678_ _08680_ _08685_ _08691_ VGND VGND VPWR VPWR _08693_ sky130_fd_sc_hd__o311a_1
XFILLER_0_65_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12576_ _02634_ _02668_ VGND VGND VPWR VPWR _02669_ sky130_fd_sc_hd__nand2_1
X_14315_ _04517_ _04518_ VGND VGND VPWR VPWR _04519_ sky130_fd_sc_hd__nor2_1
X_17103_ _07434_ _07441_ VGND VGND VPWR VPWR _07550_ sky130_fd_sc_hd__or2_1
XFILLER_0_136_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11527_ _01610_ _01618_ _01617_ VGND VGND VPWR VPWR _01620_ sky130_fd_sc_hd__o21a_1
X_18083_ _08459_ _08460_ _08540_ VGND VGND VPWR VPWR _08617_ sky130_fd_sc_hd__nand3_1
X_15295_ _05575_ _05576_ _05587_ VGND VGND VPWR VPWR _05588_ sky130_fd_sc_hd__a21o_1
XFILLER_0_135_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17034_ _06739_ _06733_ _02978_ VGND VGND VPWR VPWR _07475_ sky130_fd_sc_hd__mux2_1
X_14246_ _04434_ _04435_ _04441_ VGND VGND VPWR VPWR _04443_ sky130_fd_sc_hd__a21o_1
XFILLER_0_151_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11458_ _01518_ _01523_ VGND VGND VPWR VPWR _01551_ sky130_fd_sc_hd__and2_1
XFILLER_0_40_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10409_ cla_inst.in1\[30\] VGND VGND VPWR VPWR _00502_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_110_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14177_ _04359_ _04367_ VGND VGND VPWR VPWR _04368_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_21_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11389_ _01474_ _01481_ VGND VGND VPWR VPWR _01482_ sky130_fd_sc_hd__xnor2_4
XTAP_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13128_ _03221_ _03222_ _03223_ VGND VGND VPWR VPWR _03224_ sky130_fd_sc_hd__and3_4
XTAP_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18985_ clknet_4_0_0_clk _09381_ VGND VGND VPWR VPWR salida\[38\] sky130_fd_sc_hd__dfxtp_1
XTAP_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13059_ _08180_ _03150_ _03023_ VGND VGND VPWR VPWR _03151_ sky130_fd_sc_hd__o21ai_1
X_17936_ _07664_ net145 VGND VGND VPWR VPWR _08457_ sky130_fd_sc_hd__nand2_1
X_17867_ _08285_ _08280_ VGND VGND VPWR VPWR _08382_ sky130_fd_sc_hd__and2b_1
XFILLER_0_108_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16818_ _07237_ _07238_ VGND VGND VPWR VPWR _07239_ sky130_fd_sc_hd__or2_1
X_17798_ _07038_ _07859_ _08306_ VGND VGND VPWR VPWR _08307_ sky130_fd_sc_hd__and3_1
XFILLER_0_16_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16749_ _07162_ _02831_ _07163_ VGND VGND VPWR VPWR _07164_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_76_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18419_ _08979_ _08980_ VGND VGND VPWR VPWR _08981_ sky130_fd_sc_hd__and2_1
XFILLER_0_91_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_141_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09985_ _07788_ _09248_ _09263_ VGND VGND VPWR VPWR _09271_ sky130_fd_sc_hd__nand3_1
XFILLER_0_149_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwb_buttons_leds_157 VGND VGND VPWR VPWR wb_buttons_leds_157/HI led_enb[6] sky130_fd_sc_hd__conb_1
X_10760_ _06181_ _00822_ _00797_ _00821_ VGND VGND VPWR VPWR _00853_ sky130_fd_sc_hd__a211o_1
XFILLER_0_94_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09419_ sel_op\[2\] VGND VGND VPWR VPWR _03184_ sky130_fd_sc_hd__buf_4
XFILLER_0_94_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10691_ _04722_ _00782_ _00780_ VGND VGND VPWR VPWR _00784_ sky130_fd_sc_hd__and3_1
XFILLER_0_94_499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12430_ _02515_ net122 _02456_ _02522_ VGND VGND VPWR VPWR _02523_ sky130_fd_sc_hd__o211a_1
XFILLER_0_47_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12361_ _02452_ _02453_ VGND VGND VPWR VPWR _02454_ sky130_fd_sc_hd__nand2_1
XFILLER_0_117_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14100_ _04267_ _04268_ _04282_ VGND VGND VPWR VPWR _04283_ sky130_fd_sc_hd__o21a_2
X_11312_ _01396_ _01397_ _01398_ _01404_ VGND VGND VPWR VPWR _01405_ sky130_fd_sc_hd__o31a_1
X_15080_ _00151_ _00125_ _05964_ _06062_ VGND VGND VPWR VPWR _05353_ sky130_fd_sc_hd__and4_1
X_12292_ _02352_ net323 _02282_ _02384_ VGND VGND VPWR VPWR _02385_ sky130_fd_sc_hd__o211a_1
XFILLER_0_133_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14031_ _04192_ _04193_ _04207_ VGND VGND VPWR VPWR _04208_ sky130_fd_sc_hd__a21o_1
X_11243_ _01332_ _01333_ _01334_ _01312_ VGND VGND VPWR VPWR _01336_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_30_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11174_ _01141_ _01266_ VGND VGND VPWR VPWR _01267_ sky130_fd_sc_hd__nor2_1
XFILLER_0_101_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10125_ _00217_ VGND VGND VPWR VPWR _00218_ sky130_fd_sc_hd__clkbuf_8
X_18770_ _09285_ VGND VGND VPWR VPWR _00081_ sky130_fd_sc_hd__buf_1
X_15982_ _02992_ _03068_ VGND VGND VPWR VPWR _06330_ sky130_fd_sc_hd__nand2_1
X_17721_ _08220_ _08221_ _08218_ VGND VGND VPWR VPWR _08223_ sky130_fd_sc_hd__o21ai_1
X_10056_ cla_inst.in2\[26\] VGND VGND VPWR VPWR _00149_ sky130_fd_sc_hd__clkbuf_4
X_14933_ _05190_ _05193_ VGND VGND VPWR VPWR _05194_ sky130_fd_sc_hd__xor2_1
X_17652_ _08147_ VGND VGND VPWR VPWR _09394_ sky130_fd_sc_hd__inv_2
X_14864_ _05116_ _05117_ VGND VGND VPWR VPWR _05118_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_89_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16603_ _03169_ _06432_ VGND VGND VPWR VPWR _07006_ sky130_fd_sc_hd__or2_1
X_13815_ _03970_ _03971_ VGND VGND VPWR VPWR _03972_ sky130_fd_sc_hd__nor2_1
XFILLER_0_86_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14795_ _05041_ _05042_ VGND VGND VPWR VPWR _05043_ sky130_fd_sc_hd__xnor2_1
X_17583_ _08070_ _08072_ VGND VGND VPWR VPWR _08073_ sky130_fd_sc_hd__xor2_1
X_13746_ _03895_ _03896_ VGND VGND VPWR VPWR _03897_ sky130_fd_sc_hd__xnor2_4
X_16534_ _02975_ _03120_ _03927_ _06919_ _06930_ VGND VGND VPWR VPWR _06931_ sky130_fd_sc_hd__o311a_1
XFILLER_0_58_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10958_ _00941_ _00953_ _00954_ VGND VGND VPWR VPWR _01051_ sky130_fd_sc_hd__or3_4
XFILLER_0_70_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13677_ _03818_ VGND VGND VPWR VPWR _03821_ sky130_fd_sc_hd__inv_2
X_16465_ _06680_ _06855_ VGND VGND VPWR VPWR _06856_ sky130_fd_sc_hd__nor2_1
XFILLER_0_38_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10889_ ApproximateM_inst.lob_16.lob2.genblk1\[10\].genblk1.mux.sel _05290_ ApproximateM_inst.lob_16.lob1.genblk1\[14\].genblk1.mux.sel
+ ApproximateM_inst.lob_16.lob1.genblk1\[13\].genblk1.mux.sel VGND VGND VPWR VPWR
+ _00982_ sky130_fd_sc_hd__and4_1
XFILLER_0_26_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18204_ _08745_ _08747_ _08741_ VGND VGND VPWR VPWR _08749_ sky130_fd_sc_hd__a21o_1
X_15416_ _05545_ _05642_ VGND VGND VPWR VPWR _05719_ sky130_fd_sc_hd__and2b_1
X_12628_ _07700_ _00131_ _02720_ VGND VGND VPWR VPWR _02721_ sky130_fd_sc_hd__nand3_1
XFILLER_0_143_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16396_ _02780_ _01248_ _06673_ VGND VGND VPWR VPWR _06781_ sky130_fd_sc_hd__or3_1
XFILLER_0_109_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_538 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15347_ _05563_ _05630_ _05643_ VGND VGND VPWR VPWR _05644_ sky130_fd_sc_hd__o21a_1
XFILLER_0_5_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18135_ _01998_ _08673_ VGND VGND VPWR VPWR _08674_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_124_730 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12559_ _02644_ _02645_ _02651_ VGND VGND VPWR VPWR _02652_ sky130_fd_sc_hd__and3_1
XFILLER_0_81_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15278_ _05463_ _05471_ _05568_ VGND VGND VPWR VPWR _05569_ sky130_fd_sc_hd__a21oi_1
X_18066_ _04647_ _06445_ VGND VGND VPWR VPWR _08599_ sky130_fd_sc_hd__nand2_1
Xhold106 net101 VGND VGND VPWR VPWR net269 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold117 _00024_ VGND VGND VPWR VPWR net280 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold128 net89 VGND VGND VPWR VPWR net291 sky130_fd_sc_hd__dlygate4sd3_1
X_14229_ _04387_ _04388_ _04389_ VGND VGND VPWR VPWR _04424_ sky130_fd_sc_hd__or3_4
Xhold139 _00005_ VGND VGND VPWR VPWR net302 sky130_fd_sc_hd__dlygate4sd3_1
X_17017_ _02840_ _07353_ VGND VGND VPWR VPWR _07456_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09770_ cla_inst.in1\[26\] VGND VGND VPWR VPWR _07004_ sky130_fd_sc_hd__clkbuf_4
XTAP_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18968_ clknet_4_4_0_clk _09399_ VGND VGND VPWR VPWR salida\[21\] sky130_fd_sc_hd__dfxtp_1
XTAP_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17919_ _04337_ _06389_ _06390_ _08438_ VGND VGND VPWR VPWR _08439_ sky130_fd_sc_hd__a31o_1
XFILLER_0_119_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18899_ clknet_4_12_0_clk _00053_ VGND VGND VPWR VPWR cla_inst.in1\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_96_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_700 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_147_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_875 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_90 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09968_ _09070_ _09137_ VGND VGND VPWR VPWR _09145_ sky130_fd_sc_hd__xnor2_2
X_09899_ _04395_ VGND VGND VPWR VPWR _08409_ sky130_fd_sc_hd__buf_6
X_11930_ _02016_ _02021_ _02022_ VGND VGND VPWR VPWR _02023_ sky130_fd_sc_hd__o21a_1
XTAP_2801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11861_ _00832_ _04482_ VGND VGND VPWR VPWR _01954_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13600_ _03523_ _03525_ VGND VGND VPWR VPWR _03737_ sky130_fd_sc_hd__nor2_2
X_10812_ _00900_ _00904_ VGND VGND VPWR VPWR _00905_ sky130_fd_sc_hd__nor2_1
X_14580_ _04672_ _04674_ VGND VGND VPWR VPWR _04808_ sky130_fd_sc_hd__nand2_2
X_11792_ _01564_ _01601_ _01602_ _01603_ VGND VGND VPWR VPWR _01885_ sky130_fd_sc_hd__and4_1
XFILLER_0_138_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13531_ _08865_ _00665_ _03413_ _03412_ _00495_ VGND VGND VPWR VPWR _03661_ sky130_fd_sc_hd__a32o_1
XFILLER_0_83_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_308 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10743_ _07058_ _07091_ _05975_ _06094_ _00835_ VGND VGND VPWR VPWR _00836_ sky130_fd_sc_hd__a41o_1
XFILLER_0_55_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16250_ _03027_ _03111_ _01674_ VGND VGND VPWR VPWR _06622_ sky130_fd_sc_hd__a21o_1
X_13462_ _03434_ _03435_ _03466_ VGND VGND VPWR VPWR _03586_ sky130_fd_sc_hd__nor3_1
XFILLER_0_152_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10674_ _03728_ _04143_ VGND VGND VPWR VPWR _00767_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15201_ _05483_ _05484_ VGND VGND VPWR VPWR _05485_ sky130_fd_sc_hd__xnor2_2
X_12413_ _02505_ _00247_ _00166_ _00845_ VGND VGND VPWR VPWR _02506_ sky130_fd_sc_hd__a22o_1
XFILLER_0_23_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16181_ _06419_ _06459_ VGND VGND VPWR VPWR _06547_ sky130_fd_sc_hd__nor2_2
X_13393_ _03507_ _03508_ _03490_ VGND VGND VPWR VPWR _03511_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_3_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15132_ _02959_ _02962_ _04403_ _05409_ VGND VGND VPWR VPWR _05411_ sky130_fd_sc_hd__a211o_4
X_12344_ _02436_ _02371_ VGND VGND VPWR VPWR _02437_ sky130_fd_sc_hd__and2b_1
XFILLER_0_121_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15063_ _05332_ _00461_ _00362_ _05334_ VGND VGND VPWR VPWR _05335_ sky130_fd_sc_hd__and4b_1
XFILLER_0_50_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_120_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12275_ _02353_ _02367_ VGND VGND VPWR VPWR _02368_ sky130_fd_sc_hd__or2_1
XFILLER_0_121_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14014_ _00164_ _01695_ VGND VGND VPWR VPWR _04190_ sky130_fd_sc_hd__nand2_2
X_11226_ _07058_ _07091_ _06094_ _00460_ _01089_ VGND VGND VPWR VPWR _01319_ sky130_fd_sc_hd__a41o_1
XFILLER_0_120_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18822_ _09125_ _09325_ VGND VGND VPWR VPWR _09327_ sky130_fd_sc_hd__and2_1
XFILLER_0_4_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11157_ _01247_ _01249_ VGND VGND VPWR VPWR _01250_ sky130_fd_sc_hd__xnor2_4
X_10108_ _00190_ _00192_ _00193_ _00132_ _00200_ VGND VGND VPWR VPWR _00201_ sky130_fd_sc_hd__a41o_1
X_18753_ _09272_ VGND VGND VPWR VPWR _00076_ sky130_fd_sc_hd__clkbuf_1
X_11088_ _01166_ net144 _01179_ _01180_ VGND VGND VPWR VPWR _01181_ sky130_fd_sc_hd__o211ai_4
X_15965_ _06299_ _06301_ _06312_ VGND VGND VPWR VPWR _06313_ sky130_fd_sc_hd__nand3_1
X_17704_ _08083_ _08098_ _08204_ VGND VGND VPWR VPWR _08205_ sky130_fd_sc_hd__a21o_1
X_14916_ _05173_ _05174_ VGND VGND VPWR VPWR _05175_ sky130_fd_sc_hd__xnor2_1
X_10039_ _00131_ VGND VGND VPWR VPWR _00132_ sky130_fd_sc_hd__clkbuf_8
X_18684_ net42 _09189_ _09220_ VGND VGND VPWR VPWR _00052_ sky130_fd_sc_hd__o21a_1
X_15896_ _06195_ _06199_ VGND VGND VPWR VPWR _06239_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_59_901 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17635_ _01866_ _06510_ _02988_ VGND VGND VPWR VPWR _08130_ sky130_fd_sc_hd__and3b_1
X_14847_ _03539_ _04241_ _04079_ _05098_ VGND VGND VPWR VPWR _05099_ sky130_fd_sc_hd__a31o_1
XFILLER_0_58_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17566_ _08052_ _08053_ VGND VGND VPWR VPWR _08054_ sky130_fd_sc_hd__xor2_1
X_14778_ _09353_ _04336_ _05020_ _05021_ VGND VGND VPWR VPWR _05024_ sky130_fd_sc_hd__a22o_1
XFILLER_0_19_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_904 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_129_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16517_ _06908_ _06909_ _06910_ VGND VGND VPWR VPWR _06912_ sky130_fd_sc_hd__nor3_1
X_13729_ _03875_ _03876_ _03856_ VGND VGND VPWR VPWR _03878_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_46_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17497_ _07977_ _07978_ VGND VGND VPWR VPWR _07979_ sky130_fd_sc_hd__and2b_1
XFILLER_0_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_128_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16448_ _01264_ _06673_ VGND VGND VPWR VPWR _06837_ sky130_fd_sc_hd__nor2_1
XFILLER_0_144_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_300 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16379_ _06758_ _06761_ _00134_ VGND VGND VPWR VPWR _06762_ sky130_fd_sc_hd__o21a_2
XFILLER_0_53_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18118_ _08556_ _08559_ _08488_ VGND VGND VPWR VPWR _08655_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_5_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18049_ _08391_ _08493_ _08579_ VGND VGND VPWR VPWR _08580_ sky130_fd_sc_hd__o21a_1
XFILLER_0_111_243 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_112_799 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09822_ _07559_ VGND VGND VPWR VPWR _07570_ sky130_fd_sc_hd__buf_4
X_09753_ _06558_ _06569_ _06808_ VGND VGND VPWR VPWR _06819_ sky130_fd_sc_hd__a21o_2
X_09684_ _06040_ _06051_ _06062_ _05257_ VGND VGND VPWR VPWR _06073_ sky130_fd_sc_hd__and4_1
XFILLER_0_146_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_527 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10390_ _00468_ _00469_ _00481_ VGND VGND VPWR VPWR _00483_ sky130_fd_sc_hd__nand3_2
XFILLER_0_60_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_563 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12060_ _02052_ _02068_ _02069_ VGND VGND VPWR VPWR _02153_ sky130_fd_sc_hd__o21ai_1
X_11011_ _01093_ _01103_ VGND VGND VPWR VPWR _01104_ sky130_fd_sc_hd__xor2_1
X_12962_ _00119_ VGND VGND VPWR VPWR _03055_ sky130_fd_sc_hd__clkbuf_4
X_15750_ _06074_ _06080_ VGND VGND VPWR VPWR _06082_ sky130_fd_sc_hd__nand2_1
X_14701_ _04938_ _04832_ VGND VGND VPWR VPWR _04940_ sky130_fd_sc_hd__and2b_1
X_11913_ _01911_ _02005_ VGND VGND VPWR VPWR _02006_ sky130_fd_sc_hd__xnor2_1
X_12893_ _03574_ VGND VGND VPWR VPWR _02986_ sky130_fd_sc_hd__clkbuf_8
X_15681_ _06004_ _06005_ _05956_ VGND VGND VPWR VPWR _06007_ sky130_fd_sc_hd__o21a_1
XTAP_2620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17420_ _07771_ _07782_ _07894_ VGND VGND VPWR VPWR _07895_ sky130_fd_sc_hd__a21bo_1
X_14632_ _04730_ _04833_ _04862_ _04863_ VGND VGND VPWR VPWR _04865_ sky130_fd_sc_hd__a211o_1
XFILLER_0_68_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11844_ _01933_ _01934_ _01935_ VGND VGND VPWR VPWR _01937_ sky130_fd_sc_hd__nand3_1
XTAP_2664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14563_ _04619_ _04789_ VGND VGND VPWR VPWR _04790_ sky130_fd_sc_hd__xor2_1
XTAP_1963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17351_ _07796_ _07800_ _07819_ _06723_ _02045_ VGND VGND VPWR VPWR _09391_ sky130_fd_sc_hd__o32a_1
X_11775_ _01675_ _01864_ VGND VGND VPWR VPWR _01868_ sky130_fd_sc_hd__nor2_1
XTAP_1974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16302_ _03077_ _03029_ _02809_ VGND VGND VPWR VPWR _06679_ sky130_fd_sc_hd__a21o_1
XTAP_1996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13514_ _03639_ _03641_ _03624_ VGND VGND VPWR VPWR _03643_ sky130_fd_sc_hd__a21oi_2
X_10726_ _00817_ _00818_ VGND VGND VPWR VPWR _00819_ sky130_fd_sc_hd__nand2_1
X_14494_ _03793_ _07722_ _08169_ _03859_ VGND VGND VPWR VPWR _04714_ sky130_fd_sc_hd__a22oi_1
X_17282_ _02045_ _07743_ VGND VGND VPWR VPWR _07745_ sky130_fd_sc_hd__nor2_4
XFILLER_0_125_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_153_622 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16233_ _06462_ _06603_ VGND VGND VPWR VPWR _06604_ sky130_fd_sc_hd__nor2_1
X_13445_ _03090_ _03137_ _03566_ VGND VGND VPWR VPWR _03567_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_125_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10657_ _00747_ _00748_ _00749_ VGND VGND VPWR VPWR _00750_ sky130_fd_sc_hd__or3_4
XFILLER_0_35_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_141_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13376_ _03317_ _03331_ VGND VGND VPWR VPWR _03492_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16164_ _06528_ VGND VGND VPWR VPWR _06529_ sky130_fd_sc_hd__buf_4
X_10588_ _00358_ _07504_ _00147_ _00131_ VGND VGND VPWR VPWR _00681_ sky130_fd_sc_hd__and4_1
XFILLER_0_50_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15115_ _05390_ _05391_ VGND VGND VPWR VPWR _05392_ sky130_fd_sc_hd__nor2_1
X_12327_ _07069_ _00774_ _00909_ _07036_ VGND VGND VPWR VPWR _02420_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_133_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16095_ _03921_ _05420_ VGND VGND VPWR VPWR _06454_ sky130_fd_sc_hd__or2_1
XFILLER_0_121_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15046_ _02984_ _02988_ _00509_ _09248_ VGND VGND VPWR VPWR _05316_ sky130_fd_sc_hd__and4_2
X_12258_ _02224_ _02225_ _02227_ VGND VGND VPWR VPWR _02351_ sky130_fd_sc_hd__o21ai_1
X_11209_ _01300_ _01301_ VGND VGND VPWR VPWR _01302_ sky130_fd_sc_hd__xor2_2
X_12189_ _02231_ _02279_ _02280_ _02281_ VGND VGND VPWR VPWR _02282_ sky130_fd_sc_hd__or4_4
X_18805_ _09313_ VGND VGND VPWR VPWR _00092_ sky130_fd_sc_hd__buf_1
X_16997_ _07432_ _07433_ VGND VGND VPWR VPWR _07434_ sky130_fd_sc_hd__xnor2_1
X_18736_ _04241_ net60 _09251_ VGND VGND VPWR VPWR _09259_ sky130_fd_sc_hd__mux2_1
X_15948_ _03921_ _06292_ _06294_ VGND VGND VPWR VPWR _06295_ sky130_fd_sc_hd__a21o_1
X_18667_ net66 _09189_ _09208_ VGND VGND VPWR VPWR _00045_ sky130_fd_sc_hd__o21a_1
XFILLER_0_78_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15879_ _06219_ _06220_ VGND VGND VPWR VPWR _06221_ sky130_fd_sc_hd__and2_1
XFILLER_0_59_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17618_ _08103_ _08110_ VGND VGND VPWR VPWR _08111_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_116_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18598_ net255 _09140_ _09155_ _09144_ VGND VGND VPWR VPWR _00022_ sky130_fd_sc_hd__o211a_1
XFILLER_0_47_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17549_ _03536_ _06483_ VGND VGND VPWR VPWR _08036_ sky130_fd_sc_hd__nand2_2
XFILLER_0_129_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_447 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09805_ _07374_ VGND VGND VPWR VPWR _07384_ sky130_fd_sc_hd__buf_4
XFILLER_0_5_94 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09736_ _06602_ _06624_ VGND VGND VPWR VPWR _06635_ sky130_fd_sc_hd__and2b_1
X_09667_ _05878_ VGND VGND VPWR VPWR _05888_ sky130_fd_sc_hd__buf_4
XFILLER_0_69_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_416 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09598_ _05115_ _05126_ VGND VGND VPWR VPWR _05137_ sky130_fd_sc_hd__xnor2_2
XTAP_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11560_ _01649_ _01651_ _01650_ VGND VGND VPWR VPWR _01653_ sky130_fd_sc_hd__a21o_1
XFILLER_0_107_302 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_108_847 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10511_ _03596_ _00439_ _04395_ _03629_ VGND VGND VPWR VPWR _00604_ sky130_fd_sc_hd__a22o_1
XFILLER_0_18_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11491_ _01573_ _01574_ _01580_ VGND VGND VPWR VPWR _01584_ sky130_fd_sc_hd__a21o_1
XFILLER_0_52_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13230_ _03315_ _00735_ _03332_ VGND VGND VPWR VPWR _03333_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_107_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10442_ _00491_ _00532_ _00533_ _00534_ VGND VGND VPWR VPWR _00535_ sky130_fd_sc_hd__nand4_4
XFILLER_0_17_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13161_ _03256_ _03257_ _03242_ VGND VGND VPWR VPWR _03259_ sky130_fd_sc_hd__a21oi_1
X_10373_ _00450_ _00464_ _00463_ VGND VGND VPWR VPWR _00466_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_103_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12112_ _05399_ _05355_ _07548_ VGND VGND VPWR VPWR _02205_ sky130_fd_sc_hd__and3_1
X_13092_ _01677_ _03180_ _03183_ VGND VGND VPWR VPWR _03185_ sky130_fd_sc_hd__o21ai_1
X_12043_ _02073_ _02075_ _02076_ VGND VGND VPWR VPWR _02136_ sky130_fd_sc_hd__or3_1
X_16920_ _07347_ _07348_ _06649_ VGND VGND VPWR VPWR _07350_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_46_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16851_ _02476_ _06920_ _06921_ VGND VGND VPWR VPWR _07275_ sky130_fd_sc_hd__a21o_1
X_15802_ _06071_ _06082_ VGND VGND VPWR VPWR _06139_ sky130_fd_sc_hd__nand2_1
X_16782_ _06937_ _07143_ _07198_ VGND VGND VPWR VPWR _07200_ sky130_fd_sc_hd__or3_1
X_13994_ _03984_ _04002_ VGND VGND VPWR VPWR _04168_ sky130_fd_sc_hd__or2_1
X_18521_ _06543_ _06453_ _09084_ _09089_ VGND VGND VPWR VPWR _09090_ sky130_fd_sc_hd__a31o_1
X_15733_ _06061_ _06063_ VGND VGND VPWR VPWR _06064_ sky130_fd_sc_hd__xor2_1
X_12945_ _03036_ _03037_ VGND VGND VPWR VPWR _03038_ sky130_fd_sc_hd__nand2_1
XFILLER_0_62_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18452_ _06649_ _09014_ _09015_ VGND VGND VPWR VPWR _09017_ sky130_fd_sc_hd__and3_1
X_15664_ _05970_ _05971_ _05988_ VGND VGND VPWR VPWR _05989_ sky130_fd_sc_hd__o21ai_2
XTAP_2450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_140 _06765_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12876_ _02968_ VGND VGND VPWR VPWR _02969_ sky130_fd_sc_hd__buf_8
XTAP_2461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_151 _08762_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17403_ _07855_ _07876_ VGND VGND VPWR VPWR _07877_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_56_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_162 _08934_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14615_ _04844_ _04845_ VGND VGND VPWR VPWR _04846_ sky130_fd_sc_hd__nor2_1
XFILLER_0_96_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_173 _02646_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18383_ _06426_ _06449_ _08935_ _08939_ _08942_ VGND VGND VPWR VPWR _08943_ sky130_fd_sc_hd__o311a_1
X_11827_ _01831_ _01829_ _01830_ VGND VGND VPWR VPWR _01920_ sky130_fd_sc_hd__and3_1
XTAP_2494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15595_ _05912_ _05913_ VGND VGND VPWR VPWR _05914_ sky130_fd_sc_hd__nor2_1
XFILLER_0_55_200 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17334_ _03311_ _07355_ _02200_ VGND VGND VPWR VPWR _07802_ sky130_fd_sc_hd__or3b_1
X_14546_ _04639_ _04641_ _04770_ VGND VGND VPWR VPWR _04771_ sky130_fd_sc_hd__o21a_1
X_11758_ _01849_ _01850_ ApproximateM_inst.lob_16.lob2.genblk1\[5\].genblk1.mux.sel
+ _03914_ VGND VGND VPWR VPWR _01851_ sky130_fd_sc_hd__and4b_1
XFILLER_0_83_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10709_ _06138_ _00800_ _00799_ VGND VGND VPWR VPWR _00802_ sky130_fd_sc_hd__a21o_1
XFILLER_0_43_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17265_ _07724_ _07725_ VGND VGND VPWR VPWR _07726_ sky130_fd_sc_hd__xnor2_1
X_14477_ _04691_ _04694_ _02969_ VGND VGND VPWR VPWR _04696_ sky130_fd_sc_hd__a21o_1
X_11689_ _01771_ _01780_ _01779_ VGND VGND VPWR VPWR _01782_ sky130_fd_sc_hd__o21a_1
XFILLER_0_55_299 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_126_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19004_ clknet_4_7_0_clk _09371_ VGND VGND VPWR VPWR salida\[57\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16216_ op_code\[0\] op_code\[3\] op_code\[2\] op_code\[1\] VGND VGND VPWR VPWR _06585_
+ sky130_fd_sc_hd__or4bb_1
XFILLER_0_11_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13428_ _03088_ _03093_ _03047_ VGND VGND VPWR VPWR _03549_ sky130_fd_sc_hd__mux2_1
X_17196_ _07510_ _07529_ VGND VGND VPWR VPWR _07651_ sky130_fd_sc_hd__nor2_1
XFILLER_0_141_636 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13359_ _00183_ _04864_ _04143_ _00184_ VGND VGND VPWR VPWR _03473_ sky130_fd_sc_hd__a22oi_1
X_16147_ _06509_ VGND VGND VPWR VPWR _06510_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_122_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16078_ _02214_ _06434_ VGND VGND VPWR VPWR _06435_ sky130_fd_sc_hd__nor2_1
XFILLER_0_121_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15029_ _05296_ _05297_ VGND VGND VPWR VPWR _05298_ sky130_fd_sc_hd__or2_1
Xinput2 i_wb_addr[0] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_1
X_09521_ _04198_ _04209_ _04274_ VGND VGND VPWR VPWR _04296_ sky130_fd_sc_hd__nand3_1
XFILLER_0_79_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18719_ _09125_ VGND VGND VPWR VPWR _09245_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_36_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09452_ _03509_ _03410_ _03432_ _03531_ VGND VGND VPWR VPWR _03542_ sky130_fd_sc_hd__a22o_1
XPHY_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_870 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_137_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_734 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_136_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_144_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_117_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_112_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09719_ _06384_ _06439_ VGND VGND VPWR VPWR _06450_ sky130_fd_sc_hd__xnor2_2
X_10991_ ApproximateM_inst.lob_16.lob2.genblk1\[2\].genblk1.mux.sel _05617_ _01080_
+ _01083_ VGND VGND VPWR VPWR _01084_ sky130_fd_sc_hd__and4_1
XTAP_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12730_ _02807_ _02822_ VGND VGND VPWR VPWR _02823_ sky130_fd_sc_hd__and2_1
XTAP_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12661_ _02713_ _02715_ VGND VGND VPWR VPWR _02754_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_139_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14400_ _04463_ _04466_ VGND VGND VPWR VPWR _04611_ sky130_fd_sc_hd__nor2_1
XTAP_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11612_ _01702_ _01703_ _01669_ _01681_ VGND VGND VPWR VPWR _01705_ sky130_fd_sc_hd__o211a_1
XFILLER_0_127_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15380_ _03009_ _07668_ _01139_ _01223_ VGND VGND VPWR VPWR _05680_ sky130_fd_sc_hd__and4_1
XFILLER_0_38_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12592_ ApproximateM_inst.lob_16.lob2.mux.sel net185 VGND VGND VPWR VPWR _02685_
+ sky130_fd_sc_hd__and2_2
XFILLER_0_80_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14331_ _04533_ _04534_ _04491_ _04378_ VGND VGND VPWR VPWR _04536_ sky130_fd_sc_hd__a211o_1
X_11543_ _01633_ _01634_ _01635_ VGND VGND VPWR VPWR _01636_ sky130_fd_sc_hd__nand3_1
XFILLER_0_93_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_123_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14262_ _04283_ _04429_ _04459_ VGND VGND VPWR VPWR _04461_ sky130_fd_sc_hd__o21ai_4
X_17050_ _07488_ _07490_ VGND VGND VPWR VPWR _07491_ sky130_fd_sc_hd__nand2_1
X_11474_ _05464_ _04056_ _00563_ _05508_ VGND VGND VPWR VPWR _01567_ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_647 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13213_ _00733_ VGND VGND VPWR VPWR _03315_ sky130_fd_sc_hd__inv_2
X_16001_ _06342_ _06347_ _06348_ _06349_ VGND VGND VPWR VPWR _06350_ sky130_fd_sc_hd__and4b_1
XFILLER_0_21_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10425_ _07853_ _00513_ _00517_ _00353_ VGND VGND VPWR VPWR _00518_ sky130_fd_sc_hd__a31oi_2
X_14193_ _04382_ _04383_ _04334_ VGND VGND VPWR VPWR _04386_ sky130_fd_sc_hd__a21o_1
XFILLER_0_150_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13144_ _00622_ _00629_ _00628_ VGND VGND VPWR VPWR _03242_ sky130_fd_sc_hd__a21o_1
X_10356_ _00286_ _00287_ _00281_ VGND VGND VPWR VPWR _00449_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_131_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13075_ _03166_ _01248_ _03028_ VGND VGND VPWR VPWR _03167_ sky130_fd_sc_hd__mux2_1
X_17952_ _08472_ _08473_ _07109_ _07623_ VGND VGND VPWR VPWR _08475_ sky130_fd_sc_hd__and4bb_1
X_10287_ _00234_ _00242_ VGND VGND VPWR VPWR _00380_ sky130_fd_sc_hd__nand2_1
XFILLER_0_57_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12026_ _02115_ _02118_ VGND VGND VPWR VPWR _02119_ sky130_fd_sc_hd__xnor2_1
X_16903_ _07126_ VGND VGND VPWR VPWR _07332_ sky130_fd_sc_hd__clkbuf_4
X_17883_ _08380_ _08399_ VGND VGND VPWR VPWR _08400_ sky130_fd_sc_hd__and2_1
X_16834_ _02476_ _06510_ _02099_ VGND VGND VPWR VPWR _07257_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_88_612 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16765_ _06680_ _07175_ _07177_ _07181_ VGND VGND VPWR VPWR _07182_ sky130_fd_sc_hd__or4b_2
X_13977_ _03967_ _03977_ VGND VGND VPWR VPWR _04149_ sky130_fd_sc_hd__and2b_1
XFILLER_0_88_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18504_ _04853_ _09039_ VGND VGND VPWR VPWR _09072_ sky130_fd_sc_hd__nand2_1
X_15716_ _06035_ _06044_ VGND VGND VPWR VPWR _06045_ sky130_fd_sc_hd__xor2_1
X_12928_ _03003_ net212 _03017_ _03020_ VGND VGND VPWR VPWR _03021_ sky130_fd_sc_hd__or4_4
XFILLER_0_87_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16696_ _02533_ _07104_ _07105_ VGND VGND VPWR VPWR _07106_ sky130_fd_sc_hd__nand3_4
XFILLER_0_76_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18435_ _06408_ _06463_ _08998_ VGND VGND VPWR VPWR _09406_ sky130_fd_sc_hd__a21oi_1
X_15647_ _05855_ _05907_ VGND VGND VPWR VPWR _05970_ sky130_fd_sc_hd__and2b_1
XTAP_2280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12859_ _02942_ _02947_ VGND VGND VPWR VPWR _02952_ sky130_fd_sc_hd__or2b_1
XTAP_2291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_222 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18366_ _06649_ _08922_ _08923_ VGND VGND VPWR VPWR _08924_ sky130_fd_sc_hd__and3_1
X_15578_ _05449_ _00119_ _05850_ _05849_ VGND VGND VPWR VPWR _05895_ sky130_fd_sc_hd__a31o_1
XTAP_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17317_ _07771_ _07782_ VGND VGND VPWR VPWR _07783_ sky130_fd_sc_hd__xnor2_1
X_14529_ _04750_ _04751_ VGND VGND VPWR VPWR _04752_ sky130_fd_sc_hd__and2_1
XFILLER_0_56_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18297_ _07665_ _07650_ _07708_ _08150_ _08848_ VGND VGND VPWR VPWR _08849_ sky130_fd_sc_hd__a41o_1
XFILLER_0_43_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17248_ _06562_ _06756_ _07410_ _07706_ VGND VGND VPWR VPWR _07707_ sky130_fd_sc_hd__or4_4
XFILLER_0_114_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17179_ _07631_ VGND VGND VPWR VPWR _07632_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09504_ _04034_ _04045_ _04067_ _04099_ VGND VGND VPWR VPWR _04110_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_154_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_149_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09435_ _03345_ VGND VGND VPWR VPWR _03356_ sky130_fd_sc_hd__clkbuf_4
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_40 _01697_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_299 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_51 _03432_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_62 _04406_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_73 _06482_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_84 _08615_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_105_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_95 _08880_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10210_ _00291_ _00301_ _00302_ VGND VGND VPWR VPWR _00303_ sky130_fd_sc_hd__or3_4
X_11190_ _01281_ _01282_ VGND VGND VPWR VPWR _01283_ sky130_fd_sc_hd__xnor2_1
X_10141_ _07690_ _07842_ _07864_ _07831_ VGND VGND VPWR VPWR _00234_ sky130_fd_sc_hd__a31o_1
XFILLER_0_101_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10072_ _03673_ VGND VGND VPWR VPWR _00165_ sky130_fd_sc_hd__buf_6
XFILLER_0_100_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13900_ _04062_ _04064_ VGND VGND VPWR VPWR _04065_ sky130_fd_sc_hd__or2_1
X_14880_ _05123_ _05134_ VGND VGND VPWR VPWR _05135_ sky130_fd_sc_hd__xnor2_1
X_13831_ _03987_ _04154_ _07526_ _03988_ VGND VGND VPWR VPWR _03989_ sky130_fd_sc_hd__and4b_1
X_16550_ _06946_ VGND VGND VPWR VPWR _06947_ sky130_fd_sc_hd__clkbuf_4
X_10974_ _01063_ _01066_ VGND VGND VPWR VPWR _01067_ sky130_fd_sc_hd__xor2_2
X_13762_ _03908_ _03911_ _03913_ VGND VGND VPWR VPWR _03915_ sky130_fd_sc_hd__mux2_1
X_15501_ _01356_ _09059_ _05724_ _05723_ VGND VGND VPWR VPWR _05811_ sky130_fd_sc_hd__a31o_1
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12713_ _07788_ _07613_ _02805_ VGND VGND VPWR VPWR _02806_ sky130_fd_sc_hd__and3_1
X_16481_ _03184_ _06575_ _06871_ VGND VGND VPWR VPWR _06872_ sky130_fd_sc_hd__a21o_1
X_13693_ _00174_ _04395_ _04657_ _00184_ VGND VGND VPWR VPWR _03839_ sky130_fd_sc_hd__a22oi_1
X_18220_ _02994_ _06593_ _06594_ VGND VGND VPWR VPWR _08766_ sky130_fd_sc_hd__a21oi_1
X_15432_ _05719_ _05644_ _05735_ VGND VGND VPWR VPWR _05737_ sky130_fd_sc_hd__o21a_1
X_12644_ _02735_ _02736_ VGND VGND VPWR VPWR _02737_ sky130_fd_sc_hd__nor2_1
XFILLER_0_66_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18151_ _03120_ _06021_ _08687_ _08690_ VGND VGND VPWR VPWR _08691_ sky130_fd_sc_hd__o211a_1
XFILLER_0_25_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15363_ _02999_ _03153_ _05661_ VGND VGND VPWR VPWR _05662_ sky130_fd_sc_hd__nand3_1
X_12575_ _02655_ _02666_ _02667_ VGND VGND VPWR VPWR _02668_ sky130_fd_sc_hd__a21o_1
XFILLER_0_25_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17102_ _07546_ _07547_ VGND VGND VPWR VPWR _07549_ sky130_fd_sc_hd__nand2_1
X_14314_ _00112_ _09350_ _01005_ _08409_ VGND VGND VPWR VPWR _04518_ sky130_fd_sc_hd__and4_1
XFILLER_0_80_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11526_ _01610_ _01617_ _01618_ VGND VGND VPWR VPWR _01619_ sky130_fd_sc_hd__nor3_4
XFILLER_0_108_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18082_ _08563_ _08564_ VGND VGND VPWR VPWR _08616_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15294_ _05585_ _05586_ VGND VGND VPWR VPWR _05587_ sky130_fd_sc_hd__nand2_1
XFILLER_0_151_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17033_ _04247_ _06727_ VGND VGND VPWR VPWR _07474_ sky130_fd_sc_hd__nand2_1
X_14245_ _04434_ _04435_ _04441_ VGND VGND VPWR VPWR _04442_ sky130_fd_sc_hd__nand3_1
X_11457_ _01548_ _01549_ VGND VGND VPWR VPWR _01550_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_7_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10408_ _00499_ _00500_ VGND VGND VPWR VPWR _00501_ sky130_fd_sc_hd__nor2_1
X_14176_ _04360_ _04366_ VGND VGND VPWR VPWR _04367_ sky130_fd_sc_hd__xnor2_1
X_11388_ _01479_ _01480_ VGND VGND VPWR VPWR _01481_ sky130_fd_sc_hd__nor2_2
XFILLER_0_110_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10339_ _03651_ _03662_ _04460_ _04657_ VGND VGND VPWR VPWR _00432_ sky130_fd_sc_hd__nand4_2
X_13127_ _00611_ _00616_ _00610_ VGND VGND VPWR VPWR _03223_ sky130_fd_sc_hd__a21bo_1
XTAP_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18984_ clknet_4_3_0_clk _09380_ VGND VGND VPWR VPWR salida\[37\] sky130_fd_sc_hd__dfxtp_1
XTAP_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13058_ _03025_ _03149_ VGND VGND VPWR VPWR _03150_ sky130_fd_sc_hd__and2_1
X_17935_ _08454_ _08455_ VGND VGND VPWR VPWR _08456_ sky130_fd_sc_hd__or2_1
XFILLER_0_84_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12009_ _02092_ _02097_ VGND VGND VPWR VPWR _02102_ sky130_fd_sc_hd__or2b_1
X_17866_ _08304_ _08305_ _08307_ VGND VGND VPWR VPWR _08381_ sky130_fd_sc_hd__a21o_1
XFILLER_0_17_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16817_ _07235_ _07236_ VGND VGND VPWR VPWR _07238_ sky130_fd_sc_hd__nor2_1
X_17797_ _08304_ _08305_ VGND VGND VPWR VPWR _08306_ sky130_fd_sc_hd__xor2_1
X_16748_ _07162_ _02831_ _04238_ VGND VGND VPWR VPWR _07163_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_88_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16679_ _07087_ VGND VGND VPWR VPWR _07088_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18418_ _06408_ _08428_ _03016_ VGND VGND VPWR VPWR _08980_ sky130_fd_sc_hd__or3b_1
XFILLER_0_33_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18349_ _08904_ _08852_ _08851_ VGND VGND VPWR VPWR _08905_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_127_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput60 i_wb_data[3] VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__buf_2
XFILLER_0_114_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09984_ _07799_ _09256_ VGND VGND VPWR VPWR _09263_ sky130_fd_sc_hd__and2_4
XFILLER_0_0_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwb_buttons_leds_158 VGND VGND VPWR VPWR wb_buttons_leds_158/HI led_enb[7] sky130_fd_sc_hd__conb_1
XFILLER_0_67_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10690_ _04722_ _00780_ _00782_ VGND VGND VPWR VPWR _00783_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_54_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12360_ _02375_ _02443_ _02445_ VGND VGND VPWR VPWR _02453_ sky130_fd_sc_hd__or3_1
XFILLER_0_7_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11311_ _01401_ _01403_ VGND VGND VPWR VPWR _01404_ sky130_fd_sc_hd__xor2_1
XFILLER_0_133_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12291_ _02279_ _02280_ _02281_ _02231_ VGND VGND VPWR VPWR _02384_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_121_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14030_ _04195_ _04206_ VGND VGND VPWR VPWR _04207_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_133_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11242_ _01312_ _01332_ _01333_ _01334_ VGND VGND VPWR VPWR _01335_ sky130_fd_sc_hd__and4_1
XFILLER_0_30_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11173_ _01263_ _01265_ VGND VGND VPWR VPWR _01266_ sky130_fd_sc_hd__xor2_4
XFILLER_0_38_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10124_ _04242_ VGND VGND VPWR VPWR _00217_ sky130_fd_sc_hd__clkbuf_4
X_15981_ _03013_ _03073_ VGND VGND VPWR VPWR _06328_ sky130_fd_sc_hd__nand2_2
XFILLER_0_100_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17720_ _08218_ _08220_ _08221_ VGND VGND VPWR VPWR _08222_ sky130_fd_sc_hd__or3_1
X_10055_ cla_inst.in2\[27\] VGND VGND VPWR VPWR _00148_ sky130_fd_sc_hd__clkbuf_4
X_14932_ _05191_ _05054_ _05051_ VGND VGND VPWR VPWR _05193_ sky130_fd_sc_hd__o21ai_1
X_17651_ _08124_ _08128_ _08146_ _06463_ _03111_ VGND VGND VPWR VPWR _08147_ sky130_fd_sc_hd__a32o_1
X_14863_ _04977_ _04980_ _04978_ VGND VGND VPWR VPWR _05117_ sky130_fd_sc_hd__o21ba_1
X_16602_ _03921_ _06998_ _07003_ _06484_ VGND VGND VPWR VPWR _07005_ sky130_fd_sc_hd__o211a_1
X_13814_ _05279_ _05355_ cla_inst.in1\[29\] cla_inst.in1\[28\] VGND VGND VPWR VPWR
+ _03971_ sky130_fd_sc_hd__and4_1
X_17582_ _07109_ net146 VGND VGND VPWR VPWR _08072_ sky130_fd_sc_hd__nand2_1
X_14794_ _01505_ _05758_ VGND VGND VPWR VPWR _05042_ sky130_fd_sc_hd__nand2_1
X_16533_ _06923_ _06925_ _06929_ _06720_ VGND VGND VPWR VPWR _06930_ sky130_fd_sc_hd__and4b_1
X_13745_ _03725_ _03726_ _03724_ VGND VGND VPWR VPWR _03896_ sky130_fd_sc_hd__o21ba_2
X_10957_ _01039_ _01048_ _01049_ VGND VGND VPWR VPWR _01050_ sky130_fd_sc_hd__nor3_1
XFILLER_0_85_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16464_ _06348_ _06545_ _06854_ _03166_ VGND VGND VPWR VPWR _06855_ sky130_fd_sc_hd__a22o_1
X_13676_ _03818_ _00563_ cla_inst.in2\[28\] _03819_ VGND VGND VPWR VPWR _03820_ sky130_fd_sc_hd__and4b_1
X_10888_ _05213_ _04460_ VGND VGND VPWR VPWR _00981_ sky130_fd_sc_hd__nand2_1
X_18203_ _08741_ _08745_ _08747_ _03195_ VGND VGND VPWR VPWR _08748_ sky130_fd_sc_hd__a31o_1
X_15415_ _05651_ _05670_ VGND VGND VPWR VPWR _05718_ sky130_fd_sc_hd__or2_1
XFILLER_0_26_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12627_ _07799_ _00181_ VGND VGND VPWR VPWR _02720_ sky130_fd_sc_hd__and2_2
XFILLER_0_54_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16395_ _02780_ _06673_ _01248_ VGND VGND VPWR VPWR _06780_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_26_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18134_ _01997_ _08593_ _01995_ VGND VGND VPWR VPWR _08673_ sky130_fd_sc_hd__o21a_1
X_15346_ _05545_ _05642_ VGND VGND VPWR VPWR _05643_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_14_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12558_ _02648_ _02649_ _02650_ VGND VGND VPWR VPWR _02651_ sky130_fd_sc_hd__and3_1
XFILLER_0_26_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_124_742 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_172 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18065_ _04887_ _06394_ _06393_ VGND VGND VPWR VPWR _08598_ sky130_fd_sc_hd__a21o_1
X_11509_ _01593_ _01600_ _01585_ _01586_ VGND VGND VPWR VPWR _01602_ sky130_fd_sc_hd__o211ai_4
X_15277_ _05470_ _05465_ VGND VGND VPWR VPWR _05568_ sky130_fd_sc_hd__and2b_1
XFILLER_0_41_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12489_ _02574_ _02580_ _02581_ VGND VGND VPWR VPWR _02582_ sky130_fd_sc_hd__nor3_1
Xhold107 _00030_ VGND VGND VPWR VPWR net270 sky130_fd_sc_hd__dlygate4sd3_1
Xhold118 net98 VGND VGND VPWR VPWR net281 sky130_fd_sc_hd__dlygate4sd3_1
X_17016_ _02839_ _07454_ VGND VGND VPWR VPWR _07455_ sky130_fd_sc_hd__nor2_1
Xhold129 _00019_ VGND VGND VPWR VPWR net292 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14228_ _04387_ VGND VGND VPWR VPWR _04423_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14159_ _01745_ _01695_ _04346_ VGND VGND VPWR VPWR _04348_ sky130_fd_sc_hd__a21o_1
XTAP_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18967_ clknet_4_4_0_clk _09398_ VGND VGND VPWR VPWR salida\[20\] sky130_fd_sc_hd__dfxtp_1
XTAP_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17918_ _06420_ _08437_ VGND VGND VPWR VPWR _08438_ sky130_fd_sc_hd__nand2_1
XFILLER_0_119_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18898_ clknet_4_12_0_clk _00052_ VGND VGND VPWR VPWR cla_inst.in1\[16\] sky130_fd_sc_hd__dfxtp_2
X_17849_ _08356_ _08361_ VGND VGND VPWR VPWR _08362_ sky130_fd_sc_hd__xor2_1
XFILLER_0_89_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_712 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_119_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_134_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09967_ _09080_ _09131_ VGND VGND VPWR VPWR _09137_ sky130_fd_sc_hd__xor2_2
X_09898_ _08365_ _08376_ _08387_ VGND VGND VPWR VPWR _08398_ sky130_fd_sc_hd__nand3_1
XTAP_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11860_ _01950_ _01952_ VGND VGND VPWR VPWR _01953_ sky130_fd_sc_hd__or2_1
XFILLER_0_95_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10811_ _00900_ _00902_ _00903_ VGND VGND VPWR VPWR _00904_ sky130_fd_sc_hd__nor3_1
X_11791_ _01841_ _01881_ _01882_ _01883_ VGND VGND VPWR VPWR _01884_ sky130_fd_sc_hd__nand4_2
XFILLER_0_39_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13530_ _03653_ _03659_ VGND VGND VPWR VPWR _03660_ sky130_fd_sc_hd__xor2_2
XFILLER_0_94_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10742_ _00832_ _05704_ _00833_ _00834_ VGND VGND VPWR VPWR _00835_ sky130_fd_sc_hd__and4_1
XFILLER_0_94_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_149_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10673_ _03673_ _00764_ _00765_ VGND VGND VPWR VPWR _00766_ sky130_fd_sc_hd__a21bo_1
X_13461_ _03573_ _03583_ _02976_ VGND VGND VPWR VPWR _03584_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15200_ _01505_ _09059_ VGND VGND VPWR VPWR _05484_ sky130_fd_sc_hd__nand2_1
X_12412_ _00120_ VGND VGND VPWR VPWR _02505_ sky130_fd_sc_hd__buf_4
X_16180_ _06545_ VGND VGND VPWR VPWR _06546_ sky130_fd_sc_hd__buf_4
X_13392_ _03490_ _03507_ _03508_ VGND VGND VPWR VPWR _03510_ sky130_fd_sc_hd__nand3b_4
XFILLER_0_23_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15131_ _04947_ net117 VGND VGND VPWR VPWR _05409_ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12343_ _07788_ _00120_ _04067_ _00166_ VGND VGND VPWR VPWR _02436_ sky130_fd_sc_hd__and4_2
XFILLER_0_106_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_121_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15062_ _07504_ _05845_ _05878_ _00679_ VGND VGND VPWR VPWR _05334_ sky130_fd_sc_hd__a22o_1
X_12274_ _02356_ _02365_ _02366_ VGND VGND VPWR VPWR _02367_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_50_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14013_ _04186_ _04188_ VGND VGND VPWR VPWR _04189_ sky130_fd_sc_hd__nor2_2
X_11225_ _00846_ _01317_ _00861_ VGND VGND VPWR VPWR _01318_ sky130_fd_sc_hd__a21oi_2
X_11156_ cla_inst.in2\[20\] _01248_ VGND VGND VPWR VPWR _01249_ sky130_fd_sc_hd__nand2_2
X_18821_ _03011_ net58 _09250_ VGND VGND VPWR VPWR _09325_ sky130_fd_sc_hd__mux2_1
X_10107_ _00170_ _00194_ _00198_ _00199_ VGND VGND VPWR VPWR _00200_ sky130_fd_sc_hd__and4_1
X_18752_ _09245_ _09270_ VGND VGND VPWR VPWR _09272_ sky130_fd_sc_hd__and2_1
X_11087_ _01039_ _01049_ _01048_ VGND VGND VPWR VPWR _01180_ sky130_fd_sc_hd__o21ai_2
X_15964_ _06308_ _06311_ VGND VGND VPWR VPWR _06312_ sky130_fd_sc_hd__xnor2_1
X_17703_ _08079_ _08081_ VGND VGND VPWR VPWR _08204_ sky130_fd_sc_hd__and2_1
X_14915_ _05047_ _05048_ _05046_ VGND VGND VPWR VPWR _05174_ sky130_fd_sc_hd__o21ai_1
X_10038_ _00130_ VGND VGND VPWR VPWR _00131_ sky130_fd_sc_hd__clkbuf_8
X_18683_ _01862_ _09190_ _09191_ VGND VGND VPWR VPWR _09220_ sky130_fd_sc_hd__a21oi_1
X_15895_ _06237_ _06208_ VGND VGND VPWR VPWR _06238_ sky130_fd_sc_hd__nand2_1
X_17634_ _02988_ _06510_ _03111_ VGND VGND VPWR VPWR _08129_ sky130_fd_sc_hd__a21bo_1
X_14846_ _03117_ _05097_ VGND VGND VPWR VPWR _05098_ sky130_fd_sc_hd__and2_1
XFILLER_0_59_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17565_ _07935_ _07937_ _07934_ _06800_ VGND VGND VPWR VPWR _08053_ sky130_fd_sc_hd__a2bb2o_1
X_14777_ _05022_ VGND VGND VPWR VPWR _05023_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_743 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11989_ _05017_ _00131_ VGND VGND VPWR VPWR _02082_ sky130_fd_sc_hd__nand2_1
XFILLER_0_105_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16516_ _06908_ _06909_ _06910_ VGND VGND VPWR VPWR _06911_ sky130_fd_sc_hd__o21a_1
XFILLER_0_14_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13728_ _03856_ _03875_ _03876_ VGND VGND VPWR VPWR _03877_ sky130_fd_sc_hd__or3_2
XFILLER_0_18_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17496_ _06579_ _07124_ _07511_ _07861_ VGND VGND VPWR VPWR _07978_ sky130_fd_sc_hd__or4_4
XFILLER_0_58_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16447_ _06589_ VGND VGND VPWR VPWR _06836_ sky130_fd_sc_hd__buf_4
XFILLER_0_129_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13659_ _03797_ _03798_ _03799_ VGND VGND VPWR VPWR _03801_ sky130_fd_sc_hd__a21o_1
XFILLER_0_144_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16378_ _03313_ _06760_ VGND VGND VPWR VPWR _06761_ sky130_fd_sc_hd__nor2_1
XFILLER_0_109_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_121_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_312 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18117_ _08652_ _08653_ VGND VGND VPWR VPWR _08654_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15329_ _03534_ _03556_ _03536_ VGND VGND VPWR VPWR _05624_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_594 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18048_ _08486_ _08492_ VGND VGND VPWR VPWR _08579_ sky130_fd_sc_hd__nand2_1
XFILLER_0_69_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_255 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09821_ _07548_ VGND VGND VPWR VPWR _07559_ sky130_fd_sc_hd__clkbuf_8
X_09752_ _06667_ _06798_ VGND VGND VPWR VPWR _06808_ sky130_fd_sc_hd__xnor2_1
X_09683_ _05617_ VGND VGND VPWR VPWR _06062_ sky130_fd_sc_hd__buf_4
XTAP_2109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_107_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_134_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11010_ _01097_ _01101_ _01102_ VGND VGND VPWR VPWR _01103_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_130_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12961_ _03024_ _03053_ VGND VGND VPWR VPWR _03054_ sky130_fd_sc_hd__nand2_1
X_14700_ _04832_ _04938_ VGND VGND VPWR VPWR _04939_ sky130_fd_sc_hd__and2b_1
X_11912_ ApproximateM_inst.lob_16.lob2.genblk1\[11\].genblk1.mux.sel _00180_ VGND
+ VGND VPWR VPWR _02005_ sky130_fd_sc_hd__nand2_1
X_15680_ _05956_ _06004_ _06005_ VGND VGND VPWR VPWR _06006_ sky130_fd_sc_hd__nor3_1
XTAP_2610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12892_ _02984_ VGND VGND VPWR VPWR _02985_ sky130_fd_sc_hd__buf_4
XTAP_2621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14631_ _04860_ _04861_ _04723_ _04834_ VGND VGND VPWR VPWR _04863_ sky130_fd_sc_hd__a211oi_4
XTAP_2643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11843_ _01933_ _01934_ _01935_ VGND VGND VPWR VPWR _01936_ sky130_fd_sc_hd__a21o_1
XTAP_2654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17350_ _07256_ _07804_ _07805_ _07818_ VGND VGND VPWR VPWR _07819_ sky130_fd_sc_hd__a31o_1
XTAP_2687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14562_ _04780_ _04787_ VGND VGND VPWR VPWR _04789_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_51_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11774_ _00846_ _01866_ _01674_ VGND VGND VPWR VPWR _01867_ sky130_fd_sc_hd__a21oi_4
XTAP_1964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16301_ _06672_ _06674_ _06675_ VGND VGND VPWR VPWR _06677_ sky130_fd_sc_hd__nand3_1
XTAP_1986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13513_ _03624_ _03639_ _03641_ VGND VGND VPWR VPWR _03642_ sky130_fd_sc_hd__and3_2
X_10725_ _00810_ _00816_ _00801_ _00802_ VGND VGND VPWR VPWR _00818_ sky130_fd_sc_hd__o211ai_2
XTAP_1997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17281_ _06814_ VGND VGND VPWR VPWR _07743_ sky130_fd_sc_hd__clkbuf_4
X_14493_ _04709_ _04710_ _04705_ _04706_ VGND VGND VPWR VPWR _04713_ sky130_fd_sc_hd__a211o_1
XFILLER_0_126_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_153_634 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16232_ _06543_ _06429_ _06601_ _06546_ _06333_ VGND VGND VPWR VPWR _06603_ sky130_fd_sc_hd__a32o_1
XFILLER_0_125_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13444_ _02982_ _03141_ VGND VGND VPWR VPWR _03566_ sky130_fd_sc_hd__or2_1
X_10656_ _00578_ _00580_ VGND VGND VPWR VPWR _00749_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16163_ ApproximateM_inst.lob_16.lob1.genblk2.mux_final.sel ApproximateM_inst.lob_16.lob1.genblk1\[14\].genblk1.mux.sel
+ ApproximateM_inst.lob_16.lob1.genblk1\[13\].genblk1.mux.sel VGND VGND VPWR VPWR
+ _06528_ sky130_fd_sc_hd__or3_4
X_13375_ _03318_ _03330_ VGND VGND VPWR VPWR _03491_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10587_ _00678_ _00147_ _00132_ _00679_ VGND VGND VPWR VPWR _00680_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_140_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15114_ _05387_ _05389_ _05347_ VGND VGND VPWR VPWR _05391_ sky130_fd_sc_hd__o21a_1
X_12326_ _07221_ _07243_ _04242_ _00176_ VGND VGND VPWR VPWR _02419_ sky130_fd_sc_hd__and4_1
X_16094_ _06246_ _06452_ VGND VGND VPWR VPWR _06453_ sky130_fd_sc_hd__nand2_1
XFILLER_0_23_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_121_564 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15045_ _02988_ _03455_ _09311_ _02984_ VGND VGND VPWR VPWR _05315_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_50_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12257_ _02346_ _02349_ VGND VGND VPWR VPWR _02350_ sky130_fd_sc_hd__and2b_1
XFILLER_0_121_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11208_ _05878_ _00839_ _00838_ VGND VGND VPWR VPWR _01301_ sky130_fd_sc_hd__a21bo_1
X_12188_ _02203_ _02229_ _02228_ VGND VGND VPWR VPWR _02281_ sky130_fd_sc_hd__o21a_1
X_18804_ _09298_ _09312_ VGND VGND VPWR VPWR _09313_ sky130_fd_sc_hd__and2_1
X_11139_ _01143_ _01230_ _01229_ _01196_ VGND VGND VPWR VPWR _01232_ sky130_fd_sc_hd__a211oi_2
X_16996_ _07300_ _07327_ _07298_ VGND VGND VPWR VPWR _07433_ sky130_fd_sc_hd__o21a_1
X_18735_ _09258_ VGND VGND VPWR VPWR _00070_ sky130_fd_sc_hd__clkbuf_1
X_15947_ _03537_ _06293_ _03123_ VGND VGND VPWR VPWR _06294_ sky130_fd_sc_hd__a21o_1
X_18666_ _02099_ _09190_ _09191_ VGND VGND VPWR VPWR _09208_ sky130_fd_sc_hd__a21oi_1
X_15878_ _06193_ _06175_ _06218_ VGND VGND VPWR VPWR _06220_ sky130_fd_sc_hd__or3_1
X_17617_ _08108_ _08109_ VGND VGND VPWR VPWR _08110_ sky130_fd_sc_hd__nor2_1
X_14829_ _05077_ _05079_ VGND VGND VPWR VPWR _05080_ sky130_fd_sc_hd__nand2_1
XFILLER_0_116_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18597_ salida\[18\] _09141_ _09142_ salida\[50\] _09146_ VGND VGND VPWR VPWR _09155_
+ sky130_fd_sc_hd__a221o_1
X_17548_ _06378_ _06546_ _08034_ _03693_ VGND VGND VPWR VPWR _08035_ sky130_fd_sc_hd__a22o_1
XFILLER_0_74_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17479_ _07957_ _07958_ VGND VGND VPWR VPWR _07959_ sky130_fd_sc_hd__or2b_1
XFILLER_0_46_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_132_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_520 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09804_ cla_inst.in1\[27\] VGND VGND VPWR VPWR _07374_ sky130_fd_sc_hd__clkbuf_4
X_09735_ _05355_ _06613_ net231 _05399_ VGND VGND VPWR VPWR _06624_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_805 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09666_ _05388_ VGND VGND VPWR VPWR _05878_ sky130_fd_sc_hd__buf_4
XFILLER_0_96_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09597_ _04526_ _04602_ _04406_ VGND VGND VPWR VPWR _05126_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_38_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10510_ _00450_ _00463_ _00464_ VGND VGND VPWR VPWR _00603_ sky130_fd_sc_hd__nor3_1
XFILLER_0_108_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11490_ _01582_ _01538_ _01534_ VGND VGND VPWR VPWR _01583_ sky130_fd_sc_hd__a21o_1
XFILLER_0_107_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10441_ _00489_ _00490_ net184 net340 VGND VGND VPWR VPWR _00534_ sky130_fd_sc_hd__a211o_2
XFILLER_0_135_689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_116_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10372_ _00450_ _00463_ _00464_ VGND VGND VPWR VPWR _00465_ sky130_fd_sc_hd__or3_4
X_13160_ _03242_ _03256_ _03257_ VGND VGND VPWR VPWR _03258_ sky130_fd_sc_hd__and3_1
XFILLER_0_103_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12111_ _05235_ _00147_ _02179_ _02180_ VGND VGND VPWR VPWR _02204_ sky130_fd_sc_hd__a22oi_2
X_13091_ _03047_ _03182_ VGND VGND VPWR VPWR _03183_ sky130_fd_sc_hd__or2_1
XFILLER_0_103_586 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_130_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12042_ _02107_ _02134_ _02049_ VGND VGND VPWR VPWR _02135_ sky130_fd_sc_hd__o21ai_2
X_16850_ _06422_ _06459_ VGND VGND VPWR VPWR _07274_ sky130_fd_sc_hd__or2_2
X_15801_ _06135_ _06136_ VGND VGND VPWR VPWR _06137_ sky130_fd_sc_hd__nor2_1
X_16781_ _07196_ _07197_ VGND VGND VPWR VPWR _07198_ sky130_fd_sc_hd__xnor2_1
X_13993_ _04146_ _04147_ _04164_ VGND VGND VPWR VPWR _04167_ sky130_fd_sc_hd__or3_1
X_18520_ _03120_ _06325_ _09088_ VGND VGND VPWR VPWR _09089_ sky130_fd_sc_hd__o21ai_1
X_15732_ _06000_ _06002_ VGND VGND VPWR VPWR _06063_ sky130_fd_sc_hd__nand2_1
X_12944_ _02728_ _02965_ _03292_ _03217_ VGND VGND VPWR VPWR _03037_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_87_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18451_ _08969_ _08978_ _09013_ VGND VGND VPWR VPWR _09015_ sky130_fd_sc_hd__o21ai_1
X_15663_ _05985_ _05987_ VGND VGND VPWR VPWR _05988_ sky130_fd_sc_hd__nor2_1
XTAP_2440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_130 _04132_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12875_ _02967_ VGND VGND VPWR VPWR _02968_ sky130_fd_sc_hd__clkbuf_4
XANTENNA_141 _07091_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17402_ _07858_ _07874_ VGND VGND VPWR VPWR _07876_ sky130_fd_sc_hd__xnor2_1
XANTENNA_152 _08762_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14614_ _03859_ _03793_ _07755_ cla_inst.in1\[28\] VGND VGND VPWR VPWR _04845_ sky130_fd_sc_hd__and4_4
XTAP_2473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18382_ _05896_ _06407_ _06421_ _08940_ VGND VGND VPWR VPWR _08942_ sky130_fd_sc_hd__o211ai_1
XANTENNA_163 _08934_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11826_ _01917_ _01918_ VGND VGND VPWR VPWR _01919_ sky130_fd_sc_hd__nand2_1
XTAP_2484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15594_ _05894_ _05825_ _05911_ VGND VGND VPWR VPWR _05913_ sky130_fd_sc_hd__nor3_1
XTAP_1750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_174 _02646_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17333_ _02200_ _06510_ _02045_ VGND VGND VPWR VPWR _07801_ sky130_fd_sc_hd__a21o_1
X_14545_ _04768_ _04769_ VGND VGND VPWR VPWR _04770_ sky130_fd_sc_hd__and2_1
XTAP_1783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11757_ _05584_ _03388_ ApproximateM_inst.lob_16.lob1.genblk1\[9\].genblk1.mux.sel
+ _06008_ VGND VGND VPWR VPWR _01850_ sky130_fd_sc_hd__a22o_1
XTAP_1794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_612 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10708_ _06138_ _00799_ _00800_ VGND VGND VPWR VPWR _00801_ sky130_fd_sc_hd__nand3_2
X_17264_ _07042_ _07106_ VGND VGND VPWR VPWR _07725_ sky130_fd_sc_hd__nor2_1
X_14476_ _04691_ _04694_ VGND VGND VPWR VPWR _04695_ sky130_fd_sc_hd__nor2_1
XFILLER_0_43_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11688_ _01771_ _01779_ _01780_ VGND VGND VPWR VPWR _01781_ sky130_fd_sc_hd__nor3_4
XFILLER_0_70_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_45 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19003_ clknet_4_5_0_clk _09370_ VGND VGND VPWR VPWR salida\[56\] sky130_fd_sc_hd__dfxtp_1
X_16215_ _06561_ _06572_ _06581_ _06563_ VGND VGND VPWR VPWR _06584_ sky130_fd_sc_hd__o22a_1
X_13427_ _03544_ _03546_ _03547_ VGND VGND VPWR VPWR _03548_ sky130_fd_sc_hd__mux2_1
X_10639_ _00724_ _00731_ VGND VGND VPWR VPWR _00732_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_24_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17195_ _07649_ VGND VGND VPWR VPWR _07650_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_12_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16146_ _03239_ op_code\[3\] op_code\[2\] _03217_ VGND VGND VPWR VPWR _06509_ sky130_fd_sc_hd__and4bb_2
XFILLER_0_23_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13358_ _03267_ _03290_ VGND VGND VPWR VPWR _03472_ sky130_fd_sc_hd__and2_1
XFILLER_0_11_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12309_ _00645_ _05235_ _07570_ _07602_ VGND VGND VPWR VPWR _02402_ sky130_fd_sc_hd__and4_2
X_16077_ _06433_ VGND VGND VPWR VPWR _06434_ sky130_fd_sc_hd__inv_2
X_13289_ _03728_ _00459_ _03216_ _03215_ _05845_ VGND VGND VPWR VPWR _03396_ sky130_fd_sc_hd__a32o_1
X_15028_ _05207_ _05176_ _05295_ VGND VGND VPWR VPWR _05297_ sky130_fd_sc_hd__and3_1
XFILLER_0_20_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput3 i_wb_addr[10] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16979_ _06579_ _07313_ VGND VGND VPWR VPWR _07414_ sky130_fd_sc_hd__or2_1
X_09520_ _04198_ _04209_ _04274_ VGND VGND VPWR VPWR _04285_ sky130_fd_sc_hd__a21o_1
X_18718_ _09244_ VGND VGND VPWR VPWR _00065_ sky130_fd_sc_hd__clkbuf_1
X_09451_ _03520_ VGND VGND VPWR VPWR _03531_ sky130_fd_sc_hd__buf_8
X_18649_ _09176_ _09194_ VGND VGND VPWR VPWR _09195_ sky130_fd_sc_hd__and2_1
XFILLER_0_78_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_882 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_117_623 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_278 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_144_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_602 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_131_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09718_ _06395_ _06428_ VGND VGND VPWR VPWR _06439_ sky130_fd_sc_hd__xnor2_2
X_10990_ _01081_ cla_inst.in1\[20\] net233 _01082_ VGND VGND VPWR VPWR _01083_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09649_ cla_inst.in1\[23\] VGND VGND VPWR VPWR _05693_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_97_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12660_ _02724_ VGND VGND VPWR VPWR _02753_ sky130_fd_sc_hd__inv_2
XTAP_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11611_ _01669_ _01681_ _01702_ _01703_ VGND VGND VPWR VPWR _01704_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_93_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12591_ _02674_ _02682_ _02681_ VGND VGND VPWR VPWR _02684_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_108_612 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14330_ _04491_ _04378_ _04533_ _04534_ VGND VGND VPWR VPWR _04535_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_53_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11542_ _01573_ _01581_ VGND VGND VPWR VPWR _01635_ sky130_fd_sc_hd__nand2_1
XFILLER_0_92_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14261_ _04457_ _04458_ VGND VGND VPWR VPWR _04459_ sky130_fd_sc_hd__nor2_2
X_11473_ _05224_ _04143_ VGND VGND VPWR VPWR _01566_ sky130_fd_sc_hd__and2_1
XFILLER_0_122_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16000_ _02972_ _01264_ VGND VGND VPWR VPWR _06349_ sky130_fd_sc_hd__nand2_1
X_13212_ _03310_ _03312_ VGND VGND VPWR VPWR _03314_ sky130_fd_sc_hd__xor2_2
XFILLER_0_61_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10424_ _00515_ _00516_ VGND VGND VPWR VPWR _00517_ sky130_fd_sc_hd__nor2_4
XFILLER_0_123_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14192_ _04334_ _04382_ _04383_ VGND VGND VPWR VPWR _04385_ sky130_fd_sc_hd__nand3_4
XFILLER_0_33_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13143_ _03237_ _03238_ _00620_ net136 VGND VGND VPWR VPWR _03241_ sky130_fd_sc_hd__a211o_1
X_10355_ _00438_ _00446_ _00445_ VGND VGND VPWR VPWR _00448_ sky130_fd_sc_hd__a21o_1
XTAP_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10286_ _09339_ VGND VGND VPWR VPWR _00379_ sky130_fd_sc_hd__inv_2
X_13074_ _01264_ VGND VGND VPWR VPWR _03166_ sky130_fd_sc_hd__clkbuf_4
X_17951_ _07394_ _07604_ _07649_ _07780_ VGND VGND VPWR VPWR _08473_ sky130_fd_sc_hd__and4_1
X_12025_ _02116_ _02117_ VGND VGND VPWR VPWR _02118_ sky130_fd_sc_hd__xnor2_2
X_16902_ _07328_ _07329_ VGND VGND VPWR VPWR _07331_ sky130_fd_sc_hd__xnor2_1
X_17882_ _08397_ VGND VGND VPWR VPWR _08399_ sky130_fd_sc_hd__inv_2
X_16833_ _06508_ VGND VGND VPWR VPWR _07256_ sky130_fd_sc_hd__buf_4
X_16764_ _06424_ _07179_ _07180_ VGND VGND VPWR VPWR _07181_ sky130_fd_sc_hd__or3_1
X_13976_ _03792_ _03995_ VGND VGND VPWR VPWR _04148_ sky130_fd_sc_hd__and2_1
XFILLER_0_88_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15715_ _06036_ _06043_ VGND VGND VPWR VPWR _06044_ sky130_fd_sc_hd__xnor2_1
X_18503_ _09051_ _09057_ _09071_ _06463_ _03155_ VGND VGND VPWR VPWR _09409_ sky130_fd_sc_hd__a32oi_2
X_12927_ _03018_ _03019_ VGND VGND VPWR VPWR _03020_ sky130_fd_sc_hd__or2_1
X_16695_ _06812_ _06575_ _06871_ VGND VGND VPWR VPWR _07105_ sky130_fd_sc_hd__o21ai_4
X_15646_ _05914_ _05926_ VGND VGND VPWR VPWR _05969_ sky130_fd_sc_hd__and2_1
X_18434_ _06559_ _08977_ _08978_ _08997_ VGND VGND VPWR VPWR _08998_ sky130_fd_sc_hd__o31a_1
X_12858_ _02949_ _02950_ VGND VGND VPWR VPWR _02951_ sky130_fd_sc_hd__or2_1
XTAP_2270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11809_ _01900_ _01899_ _01812_ _01811_ VGND VGND VPWR VPWR _01902_ sky130_fd_sc_hd__o211ai_1
X_18365_ _08873_ _08893_ _08921_ VGND VGND VPWR VPWR _08923_ sky130_fd_sc_hd__o21ai_1
X_15577_ _05767_ _05822_ VGND VGND VPWR VPWR _05894_ sky130_fd_sc_hd__and2b_1
XFILLER_0_28_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_852 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12789_ _02871_ _02881_ VGND VGND VPWR VPWR _02882_ sky130_fd_sc_hd__and2_1
XFILLER_0_113_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17316_ _07779_ _07781_ VGND VGND VPWR VPWR _07782_ sky130_fd_sc_hd__xnor2_2
X_14528_ _04743_ _04749_ VGND VGND VPWR VPWR _04751_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_896 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18296_ _04023_ _07516_ _08260_ VGND VGND VPWR VPWR _08848_ sky130_fd_sc_hd__or3_2
XFILLER_0_126_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17247_ _02059_ _06889_ VGND VGND VPWR VPWR _07706_ sky130_fd_sc_hd__nand2_4
X_14459_ _04628_ _04629_ _04674_ _04675_ VGND VGND VPWR VPWR _04676_ sky130_fd_sc_hd__or4bb_4
XFILLER_0_52_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17178_ _06944_ _06957_ _07115_ _07035_ VGND VGND VPWR VPWR _07631_ sky130_fd_sc_hd__or4_1
XFILLER_0_3_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16129_ _08180_ _03144_ VGND VGND VPWR VPWR _06490_ sky130_fd_sc_hd__or2_1
XFILLER_0_12_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_191 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09503_ _04088_ VGND VGND VPWR VPWR _04099_ sky130_fd_sc_hd__buf_6
XFILLER_0_149_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_679 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09434_ cla_inst.in2\[19\] VGND VGND VPWR VPWR _03345_ sky130_fd_sc_hd__buf_6
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_137_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_30 _01225_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_41 _01697_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_52 _03618_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_63 _04414_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_74 _06554_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_85 _08750_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_96 _08880_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10140_ _00144_ _00155_ VGND VGND VPWR VPWR _00233_ sky130_fd_sc_hd__nand2_1
X_10071_ _00163_ VGND VGND VPWR VPWR _00164_ sky130_fd_sc_hd__clkbuf_8
X_13830_ _09172_ _03673_ _00211_ _09166_ VGND VGND VPWR VPWR _03988_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13761_ _03912_ VGND VGND VPWR VPWR _03913_ sky130_fd_sc_hd__buf_4
X_10973_ _00439_ _01064_ _01065_ VGND VGND VPWR VPWR _01066_ sky130_fd_sc_hd__a21bo_1
X_15500_ _05734_ _05733_ VGND VGND VPWR VPWR _05810_ sky130_fd_sc_hd__and2b_1
XFILLER_0_85_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12712_ _00120_ _07559_ VGND VGND VPWR VPWR _02805_ sky130_fd_sc_hd__and2_2
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16480_ _06870_ VGND VGND VPWR VPWR _06871_ sky130_fd_sc_hd__buf_4
XFILLER_0_97_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13692_ _03669_ _03652_ VGND VGND VPWR VPWR _03838_ sky130_fd_sc_hd__and2b_1
XFILLER_0_38_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15431_ _05733_ _05734_ VGND VGND VPWR VPWR _05735_ sky130_fd_sc_hd__xnor2_1
X_12643_ _02689_ _02734_ VGND VGND VPWR VPWR _02736_ sky130_fd_sc_hd__nor2_1
XFILLER_0_93_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18150_ _07089_ _08141_ _08689_ _06721_ VGND VGND VPWR VPWR _08690_ sky130_fd_sc_hd__o211a_1
XFILLER_0_38_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15362_ _05658_ _05659_ VGND VGND VPWR VPWR _05661_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_81_822 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12574_ _02656_ _02665_ VGND VGND VPWR VPWR _02667_ sky130_fd_sc_hd__and2b_1
X_17101_ _07536_ _07538_ _07545_ VGND VGND VPWR VPWR _07547_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_142_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14313_ _03321_ _01005_ _01575_ _03322_ VGND VGND VPWR VPWR _04517_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_124_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11525_ _01607_ _01608_ _01609_ VGND VGND VPWR VPWR _01618_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_123_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18081_ _08502_ _08585_ VGND VGND VPWR VPWR _08614_ sky130_fd_sc_hd__nor2_1
XFILLER_0_151_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15293_ _02999_ _03071_ _05583_ VGND VGND VPWR VPWR _05586_ sky130_fd_sc_hd__a21o_1
X_17032_ _06680_ _07471_ VGND VGND VPWR VPWR _07473_ sky130_fd_sc_hd__nor2_1
XFILLER_0_123_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14244_ _04439_ _04440_ VGND VGND VPWR VPWR _04441_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_151_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11456_ _01527_ _01529_ VGND VGND VPWR VPWR _01549_ sky130_fd_sc_hd__nand2_1
XFILLER_0_150_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10407_ _07047_ _07080_ _09303_ _07722_ VGND VGND VPWR VPWR _00500_ sky130_fd_sc_hd__and4_1
X_14175_ _04364_ _04365_ VGND VGND VPWR VPWR _04366_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_110_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11387_ _01478_ _01475_ _01476_ VGND VGND VPWR VPWR _01480_ sky130_fd_sc_hd__nor3_1
XFILLER_0_0_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13126_ _03213_ _03214_ _03220_ VGND VGND VPWR VPWR _03222_ sky130_fd_sc_hd__a21o_1
X_10338_ _00291_ _00301_ _00302_ VGND VGND VPWR VPWR _00431_ sky130_fd_sc_hd__nor3_2
XTAP_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_191 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18983_ clknet_4_1_0_clk _09379_ VGND VGND VPWR VPWR salida\[36\] sky130_fd_sc_hd__dfxtp_1
XTAP_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13057_ _00339_ VGND VGND VPWR VPWR _03149_ sky130_fd_sc_hd__buf_4
X_17934_ _07751_ _07595_ _08453_ VGND VGND VPWR VPWR _08455_ sky130_fd_sc_hd__and3_1
X_10269_ _07526_ VGND VGND VPWR VPWR _00362_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_84_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12008_ _02034_ _02100_ VGND VGND VPWR VPWR _02101_ sky130_fd_sc_hd__nor2_1
X_17865_ _08378_ _08379_ VGND VGND VPWR VPWR _08380_ sky130_fd_sc_hd__xor2_1
XFILLER_0_84_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16816_ _07235_ _07236_ VGND VGND VPWR VPWR _07237_ sky130_fd_sc_hd__and2_1
X_17796_ _08190_ _08193_ _08189_ VGND VGND VPWR VPWR _08305_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_17_86 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13959_ _03951_ _03959_ VGND VGND VPWR VPWR _04129_ sky130_fd_sc_hd__nand2_1
X_16747_ _02832_ _02801_ VGND VGND VPWR VPWR _07162_ sky130_fd_sc_hd__and2b_1
X_16678_ _06726_ _06729_ _03098_ VGND VGND VPWR VPWR _07087_ sky130_fd_sc_hd__mux2_1
XFILLER_0_146_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18417_ _03016_ _06512_ _06408_ VGND VGND VPWR VPWR _08979_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_119_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15629_ _05796_ _05949_ _05950_ VGND VGND VPWR VPWR _05951_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_57_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18348_ _08847_ VGND VGND VPWR VPWR _08904_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18279_ _04238_ _08820_ _08824_ _08829_ VGND VGND VPWR VPWR _08830_ sky130_fd_sc_hd__o211a_1
XFILLER_0_154_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput50 i_wb_data[23] VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__buf_1
XFILLER_0_130_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput61 i_wb_data[4] VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__buf_2
XFILLER_0_114_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_149_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09983_ cla_inst.in1\[30\] VGND VGND VPWR VPWR _09256_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_110_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_218 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwb_buttons_leds_159 VGND VGND VPWR VPWR wb_buttons_leds_159/HI led_enb[8] sky130_fd_sc_hd__conb_1
XFILLER_0_79_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_885 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_118_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11310_ _01319_ _01323_ _01402_ VGND VGND VPWR VPWR _01403_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_62_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12290_ _02352_ _02380_ _02381_ _02382_ VGND VGND VPWR VPWR _02383_ sky130_fd_sc_hd__nor4_2
XFILLER_0_133_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_132_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_752 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11241_ _01310_ _01311_ net220 _01020_ VGND VGND VPWR VPWR _01334_ sky130_fd_sc_hd__a211o_2
X_11172_ _00163_ _01264_ VGND VGND VPWR VPWR _01265_ sky130_fd_sc_hd__nand2_2
XFILLER_0_101_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10123_ _00184_ _00183_ _00171_ _00177_ VGND VGND VPWR VPWR _00216_ sky130_fd_sc_hd__and4_1
XFILLER_0_100_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15980_ _00908_ _02963_ VGND VGND VPWR VPWR _06327_ sky130_fd_sc_hd__or2_1
XFILLER_0_100_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14931_ _05036_ _05037_ _05049_ VGND VGND VPWR VPWR _05191_ sky130_fd_sc_hd__and3_1
X_10054_ _00146_ VGND VGND VPWR VPWR _00147_ sky130_fd_sc_hd__buf_4
X_14862_ _05113_ _05114_ VGND VGND VPWR VPWR _05116_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_89_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17650_ _08135_ _08138_ _08145_ VGND VGND VPWR VPWR _08146_ sky130_fd_sc_hd__and3_1
X_13813_ _05301_ _07755_ cla_inst.in1\[28\] _05410_ VGND VGND VPWR VPWR _03970_ sky130_fd_sc_hd__a22oi_1
X_16601_ _03921_ _07002_ VGND VGND VPWR VPWR _07003_ sky130_fd_sc_hd__nand2_1
X_17581_ _08068_ _08069_ VGND VGND VPWR VPWR _08070_ sky130_fd_sc_hd__nand2_1
X_14793_ _05038_ _05040_ VGND VGND VPWR VPWR _05041_ sky130_fd_sc_hd__nor2_1
X_16532_ _06344_ _06346_ _06926_ _06927_ _06598_ VGND VGND VPWR VPWR _06929_ sky130_fd_sc_hd__a311o_1
X_13744_ _03893_ _03894_ VGND VGND VPWR VPWR _03895_ sky130_fd_sc_hd__nor2_2
XFILLER_0_58_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10956_ _01022_ _01023_ _01038_ VGND VGND VPWR VPWR _01049_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_57_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16463_ _02972_ _06592_ _06551_ VGND VGND VPWR VPWR _06854_ sky130_fd_sc_hd__a21o_1
X_13675_ cla_inst.in2\[29\] _03432_ _00205_ cla_inst.in2\[30\] VGND VGND VPWR VPWR
+ _03819_ sky130_fd_sc_hd__a22o_1
X_10887_ net195 _00955_ _00978_ _00979_ VGND VGND VPWR VPWR _00980_ sky130_fd_sc_hd__o211a_1
X_15414_ _05646_ _05650_ VGND VGND VPWR VPWR _05717_ sky130_fd_sc_hd__nand2_1
X_18202_ _08018_ _08415_ _08743_ VGND VGND VPWR VPWR _08747_ sky130_fd_sc_hd__or3_4
XFILLER_0_72_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12626_ _02716_ _02718_ VGND VGND VPWR VPWR _02719_ sky130_fd_sc_hd__xnor2_2
X_16394_ _06582_ _06665_ _06774_ VGND VGND VPWR VPWR _06779_ sky130_fd_sc_hd__or3b_4
X_18133_ _08669_ _08671_ VGND VGND VPWR VPWR _08672_ sky130_fd_sc_hd__nand2_1
X_15345_ _05631_ _05641_ VGND VGND VPWR VPWR _05642_ sky130_fd_sc_hd__xor2_1
XFILLER_0_53_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12557_ _02608_ _02647_ VGND VGND VPWR VPWR _02650_ sky130_fd_sc_hd__or2_1
XFILLER_0_13_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18064_ _04887_ _06393_ _06394_ VGND VGND VPWR VPWR _08597_ sky130_fd_sc_hd__nand3_1
X_11508_ _01585_ _01586_ _01593_ _01600_ VGND VGND VPWR VPWR _01601_ sky130_fd_sc_hd__a211o_1
XFILLER_0_124_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15276_ _05452_ _05566_ VGND VGND VPWR VPWR _05567_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_112_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12488_ _02521_ _02579_ _02570_ _02578_ VGND VGND VPWR VPWR _02581_ sky130_fd_sc_hd__o211a_1
Xhold108 net113 VGND VGND VPWR VPWR net271 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17015_ _02837_ _02838_ VGND VGND VPWR VPWR _07454_ sky130_fd_sc_hd__nor2_1
X_14227_ _04421_ _04353_ VGND VGND VPWR VPWR _04422_ sky130_fd_sc_hd__nand2_1
Xhold119 _00027_ VGND VGND VPWR VPWR net282 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11439_ _03717_ _00197_ _01510_ _01531_ VGND VGND VPWR VPWR _01532_ sky130_fd_sc_hd__a31o_1
X_14158_ _02999_ _01695_ _04346_ VGND VGND VPWR VPWR _04347_ sky130_fd_sc_hd__nand3_1
XFILLER_0_21_284 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13109_ _00747_ _00748_ _00749_ VGND VGND VPWR VPWR _03203_ sky130_fd_sc_hd__nor3_2
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14089_ _02986_ _05975_ _04269_ _04270_ VGND VGND VPWR VPWR _04271_ sky130_fd_sc_hd__nand4_4
XTAP_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18966_ clknet_4_5_0_clk _09396_ VGND VGND VPWR VPWR salida\[19\] sky130_fd_sc_hd__dfxtp_1
XTAP_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17917_ _04337_ _06390_ _06389_ VGND VGND VPWR VPWR _08437_ sky130_fd_sc_hd__a21o_1
X_18897_ clknet_4_11_0_clk _00051_ VGND VGND VPWR VPWR ApproximateM_inst.lob_16.lob1.genblk2.mux_final.sel
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17848_ _08358_ _08359_ _08360_ VGND VGND VPWR VPWR _08361_ sky130_fd_sc_hd__or3_1
X_17779_ _08280_ _08285_ VGND VGND VPWR VPWR _08286_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_89_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_119_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_170 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_674 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_114_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09966_ _09091_ _09123_ VGND VGND VPWR VPWR _09131_ sky130_fd_sc_hd__xnor2_2
X_09897_ _06213_ _06224_ _06202_ VGND VGND VPWR VPWR _08387_ sky130_fd_sc_hd__a21bo_1
XTAP_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_903 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10810_ _00430_ _00899_ _00893_ _00898_ VGND VGND VPWR VPWR _00903_ sky130_fd_sc_hd__o211a_1
X_11790_ _01540_ _01880_ _01879_ VGND VGND VPWR VPWR _01883_ sky130_fd_sc_hd__a21o_1
XFILLER_0_94_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10741_ _07973_ cla_inst.in1\[22\] _08746_ _07984_ VGND VGND VPWR VPWR _00834_ sky130_fd_sc_hd__a22o_1
XFILLER_0_95_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_276 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13460_ _03577_ _03582_ _03079_ VGND VGND VPWR VPWR _03583_ sky130_fd_sc_hd__mux2_1
X_10672_ _03782_ _03399_ _03476_ _03848_ VGND VGND VPWR VPWR _00765_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12411_ _02436_ _02502_ VGND VGND VPWR VPWR _02504_ sky130_fd_sc_hd__or2_1
X_13391_ _03491_ _03492_ _03506_ VGND VGND VPWR VPWR _03508_ sky130_fd_sc_hd__nand3_2
XFILLER_0_152_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15130_ _05199_ _05077_ _05198_ _05302_ VGND VGND VPWR VPWR _05408_ sky130_fd_sc_hd__nor4_1
X_12342_ _02433_ _02434_ VGND VGND VPWR VPWR _02435_ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15061_ _03008_ _07515_ _05856_ _05878_ VGND VGND VPWR VPWR _05332_ sky130_fd_sc_hd__and4_1
XFILLER_0_105_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12273_ _02361_ _02364_ VGND VGND VPWR VPWR _02366_ sky130_fd_sc_hd__and2b_1
X_14012_ _04174_ _04016_ _04185_ VGND VGND VPWR VPWR _04188_ sky130_fd_sc_hd__and3_1
X_11224_ _00318_ VGND VGND VPWR VPWR _01317_ sky130_fd_sc_hd__buf_4
X_18820_ _09324_ VGND VGND VPWR VPWR _00097_ sky130_fd_sc_hd__buf_1
X_11155_ _00134_ VGND VGND VPWR VPWR _01248_ sky130_fd_sc_hd__clkbuf_8
X_10106_ _00183_ _00181_ _00197_ _00173_ VGND VGND VPWR VPWR _00199_ sky130_fd_sc_hd__a22o_1
X_18751_ _02533_ net65 _09251_ VGND VGND VPWR VPWR _09270_ sky130_fd_sc_hd__mux2_1
X_11086_ _01039_ _01048_ _01049_ VGND VGND VPWR VPWR _01179_ sky130_fd_sc_hd__or3_4
X_15963_ _06282_ _06310_ VGND VGND VPWR VPWR _06311_ sky130_fd_sc_hd__or2_1
X_17702_ _08185_ _08201_ VGND VGND VPWR VPWR _08203_ sky130_fd_sc_hd__xor2_1
X_14914_ _05171_ _05172_ VGND VGND VPWR VPWR _05173_ sky130_fd_sc_hd__nand2_1
X_10037_ _00129_ VGND VGND VPWR VPWR _00130_ sky130_fd_sc_hd__buf_6
X_18682_ net41 _09189_ _09218_ VGND VGND VPWR VPWR _00051_ sky130_fd_sc_hd__o21a_1
X_15894_ _06156_ _06204_ VGND VGND VPWR VPWR _06237_ sky130_fd_sc_hd__or2_1
X_17633_ _02848_ _08125_ _08127_ VGND VGND VPWR VPWR _08128_ sky130_fd_sc_hd__a21o_2
X_14845_ _04077_ _04083_ _02978_ VGND VGND VPWR VPWR _05097_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14776_ _09352_ _00460_ _05020_ _05021_ VGND VGND VPWR VPWR _05022_ sky130_fd_sc_hd__and4_1
X_17564_ _08050_ _08051_ VGND VGND VPWR VPWR _08052_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_85_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11988_ _01990_ _02000_ _02080_ VGND VGND VPWR VPWR _02081_ sky130_fd_sc_hd__and3_1
XFILLER_0_147_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13727_ _03857_ _03858_ _03874_ VGND VGND VPWR VPWR _03876_ sky130_fd_sc_hd__and3_1
XFILLER_0_58_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16515_ _06839_ _06840_ _06838_ VGND VGND VPWR VPWR _06910_ sky130_fd_sc_hd__a21oi_2
X_10939_ _03454_ _01031_ VGND VGND VPWR VPWR _01032_ sky130_fd_sc_hd__and2_1
X_17495_ _07124_ _07511_ _07861_ _06581_ VGND VGND VPWR VPWR _07977_ sky130_fd_sc_hd__o22a_1
XFILLER_0_14_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13658_ _03797_ _03798_ _03799_ VGND VGND VPWR VPWR _03800_ sky130_fd_sc_hd__nand3_2
XFILLER_0_45_129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16446_ _06649_ _06834_ VGND VGND VPWR VPWR _06835_ sky130_fd_sc_hd__nand2_1
XFILLER_0_144_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12609_ _02650_ net203 VGND VGND VPWR VPWR _02702_ sky130_fd_sc_hd__xnor2_1
XPHY_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16377_ _06529_ _06565_ _06759_ _06520_ VGND VGND VPWR VPWR _06760_ sky130_fd_sc_hd__o22a_1
XFILLER_0_121_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13589_ _03722_ _03723_ _03469_ _03516_ VGND VGND VPWR VPWR _03725_ sky130_fd_sc_hd__o211a_1
XFILLER_0_81_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15328_ _03538_ _03121_ VGND VGND VPWR VPWR _05623_ sky130_fd_sc_hd__nor2_2
XFILLER_0_124_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18116_ _08650_ _08651_ VGND VGND VPWR VPWR _08653_ sky130_fd_sc_hd__or2_1
XFILLER_0_41_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_152_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15259_ _05536_ _05547_ VGND VGND VPWR VPWR _05548_ sky130_fd_sc_hd__xor2_1
X_18047_ _08576_ _08577_ VGND VGND VPWR VPWR _08578_ sky130_fd_sc_hd__or2_1
XFILLER_0_112_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09820_ ApproximateM_inst.lob_16.lob1.genblk1\[1\].genblk1.mux.sel VGND VGND VPWR
+ VPWR _07548_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_39_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09751_ _06743_ _06787_ VGND VGND VPWR VPWR _06798_ sky130_fd_sc_hd__nor2_1
X_18949_ clknet_4_5_0_clk _09408_ VGND VGND VPWR VPWR salida\[2\] sky130_fd_sc_hd__dfxtp_2
X_09682_ _05649_ VGND VGND VPWR VPWR _06051_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_146_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_120 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_310 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_146_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_611 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_278 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_130_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09949_ _06646_ _06656_ VGND VGND VPWR VPWR _08951_ sky130_fd_sc_hd__and2_1
X_12960_ _03027_ _03052_ _01224_ VGND VGND VPWR VPWR _03053_ sky130_fd_sc_hd__a21o_1
X_11911_ _04548_ _00197_ _02003_ VGND VGND VPWR VPWR _02004_ sky130_fd_sc_hd__and3_1
X_12891_ _03629_ VGND VGND VPWR VPWR _02984_ sky130_fd_sc_hd__buf_4
XTAP_2600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14630_ _04723_ _04834_ _04860_ _04861_ VGND VGND VPWR VPWR _04862_ sky130_fd_sc_hd__o211a_4
XTAP_2633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11842_ _01837_ _01838_ VGND VGND VPWR VPWR _01935_ sky130_fd_sc_hd__xnor2_1
XTAP_2644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14561_ _04781_ _04786_ VGND VGND VPWR VPWR _04787_ sky130_fd_sc_hd__xnor2_1
XTAP_1943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11773_ _06482_ VGND VGND VPWR VPWR _01866_ sky130_fd_sc_hd__clkbuf_8
XTAP_1954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13512_ _03637_ _03638_ _03630_ VGND VGND VPWR VPWR _03641_ sky130_fd_sc_hd__a21o_1
X_16300_ _06672_ _06674_ _06675_ VGND VGND VPWR VPWR _06676_ sky130_fd_sc_hd__a21o_1
XTAP_1976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10724_ _00801_ _00802_ _00810_ _00816_ VGND VGND VPWR VPWR _00817_ sky130_fd_sc_hd__a211o_1
XFILLER_0_83_736 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17280_ _06561_ _07124_ _07314_ _07741_ VGND VGND VPWR VPWR _07742_ sky130_fd_sc_hd__or4_4
X_14492_ _04705_ _04706_ _04709_ _04710_ VGND VGND VPWR VPWR _04712_ sky130_fd_sc_hd__o211ai_4
XTAP_1998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16231_ _01746_ _03029_ VGND VGND VPWR VPWR _06601_ sky130_fd_sc_hd__or2_1
X_13443_ _03538_ _03564_ VGND VGND VPWR VPWR _03565_ sky130_fd_sc_hd__nand2_1
XFILLER_0_126_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10655_ _00745_ _00746_ _00537_ net124 VGND VGND VPWR VPWR _00748_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_153_646 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_540 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16162_ _06522_ _06525_ _01113_ VGND VGND VPWR VPWR _06527_ sky130_fd_sc_hd__a21oi_4
X_13374_ _03488_ _03489_ VGND VGND VPWR VPWR _03490_ sky130_fd_sc_hd__xor2_2
XFILLER_0_51_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10586_ _09166_ VGND VGND VPWR VPWR _00679_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_140_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15113_ _05347_ _05387_ _05389_ VGND VGND VPWR VPWR _05390_ sky130_fd_sc_hd__nor3_2
X_12325_ _02356_ _02365_ VGND VGND VPWR VPWR _02418_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_134_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16093_ _03155_ _06451_ VGND VGND VPWR VPWR _06452_ sky130_fd_sc_hd__and2_1
X_15044_ _02987_ _00495_ _05214_ VGND VGND VPWR VPWR _05314_ sky130_fd_sc_hd__and3_1
X_12256_ _02190_ _02348_ VGND VGND VPWR VPWR _02349_ sky130_fd_sc_hd__and2_1
XFILLER_0_121_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11207_ _06711_ _00460_ VGND VGND VPWR VPWR _01300_ sky130_fd_sc_hd__nand2_1
XFILLER_0_76_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12187_ _02277_ _02278_ _02254_ _02264_ VGND VGND VPWR VPWR _02280_ sky130_fd_sc_hd__o211a_1
X_18803_ _02994_ net51 _09301_ VGND VGND VPWR VPWR _09312_ sky130_fd_sc_hd__mux2_1
X_11138_ _01196_ _01229_ _01230_ _01143_ VGND VGND VPWR VPWR _01231_ sky130_fd_sc_hd__o211a_1
X_16995_ _07430_ _07431_ VGND VGND VPWR VPWR _07432_ sky130_fd_sc_hd__or2_1
X_18734_ _09245_ _09257_ VGND VGND VPWR VPWR _09258_ sky130_fd_sc_hd__and2_1
X_11069_ _01159_ _01160_ _01161_ VGND VGND VPWR VPWR _01162_ sky130_fd_sc_hd__o21a_1
X_15946_ _03917_ _03908_ _02979_ VGND VGND VPWR VPWR _06293_ sky130_fd_sc_hd__mux2_1
X_18665_ _09207_ VGND VGND VPWR VPWR _00044_ sky130_fd_sc_hd__buf_1
X_15877_ _06193_ _06175_ _06218_ VGND VGND VPWR VPWR _06219_ sky130_fd_sc_hd__o21ai_1
X_17616_ _08106_ _08107_ VGND VGND VPWR VPWR _08109_ sky130_fd_sc_hd__and2_1
X_14828_ _05078_ _04953_ VGND VGND VPWR VPWR _05079_ sky130_fd_sc_hd__and2_1
X_18596_ net275 _09140_ _09154_ _09144_ VGND VGND VPWR VPWR _00021_ sky130_fd_sc_hd__o211a_1
XFILLER_0_148_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17547_ _02989_ _06920_ _06921_ VGND VGND VPWR VPWR _08034_ sky130_fd_sc_hd__a21o_1
X_14759_ _00678_ _08452_ _01005_ _00679_ VGND VGND VPWR VPWR _05003_ sky130_fd_sc_hd__a22o_1
XFILLER_0_74_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17478_ _06957_ _07035_ _07195_ _07608_ VGND VGND VPWR VPWR _07958_ sky130_fd_sc_hd__or4_1
XFILLER_0_128_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_116_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_698 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16429_ _06815_ VGND VGND VPWR VPWR _06816_ sky130_fd_sc_hd__buf_2
XFILLER_0_116_326 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_128_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_112_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09803_ _07352_ VGND VGND VPWR VPWR _07363_ sky130_fd_sc_hd__buf_4
XFILLER_0_66_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09734_ cla_inst.in1\[20\] VGND VGND VPWR VPWR _06613_ sky130_fd_sc_hd__buf_6
X_09665_ _05834_ _05856_ _05475_ _05519_ VGND VGND VPWR VPWR _05867_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09596_ _05006_ _05104_ VGND VGND VPWR VPWR _05115_ sky130_fd_sc_hd__xnor2_2
XTAP_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_135_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10440_ _00349_ _00531_ _00529_ _00530_ VGND VGND VPWR VPWR _00533_ sky130_fd_sc_hd__a211o_1
XFILLER_0_122_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10371_ _00447_ _00448_ _00449_ VGND VGND VPWR VPWR _00464_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_131_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12110_ _02198_ _02199_ _02202_ VGND VGND VPWR VPWR _02203_ sky130_fd_sc_hd__and3_1
X_13090_ _02370_ _03181_ _03022_ VGND VGND VPWR VPWR _03182_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_103_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12041_ _02122_ _02132_ _02107_ _02133_ VGND VGND VPWR VPWR _02134_ sky130_fd_sc_hd__a211oi_2
X_15800_ _06065_ _06068_ _06133_ VGND VGND VPWR VPWR _06136_ sky130_fd_sc_hd__nor3_1
X_13992_ _04146_ _04147_ _04164_ VGND VGND VPWR VPWR _04166_ sky130_fd_sc_hd__o21ai_1
X_16780_ _06572_ _07106_ VGND VGND VPWR VPWR _07197_ sky130_fd_sc_hd__nor2_1
XFILLER_0_99_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15731_ _06034_ _06060_ VGND VGND VPWR VPWR _06061_ sky130_fd_sc_hd__xor2_1
X_12943_ _08865_ VGND VGND VPWR VPWR _03036_ sky130_fd_sc_hd__clkbuf_4
X_18450_ _08969_ _08978_ _09013_ VGND VGND VPWR VPWR _09014_ sky130_fd_sc_hd__or3_1
X_15662_ _05903_ _05905_ _05984_ VGND VGND VPWR VPWR _05987_ sky130_fd_sc_hd__nor3_1
XANTENNA_120 _02188_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12874_ _02965_ _02966_ VGND VGND VPWR VPWR _02967_ sky130_fd_sc_hd__or2_1
XTAP_2430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_131 _04132_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17401_ _07866_ _07873_ VGND VGND VPWR VPWR _07874_ sky130_fd_sc_hd__xnor2_1
XANTENNA_142 _08180_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14613_ _03793_ _09303_ _00498_ _03859_ VGND VGND VPWR VPWR _04844_ sky130_fd_sc_hd__a22oi_1
X_11825_ _01877_ _01878_ VGND VGND VPWR VPWR _01918_ sky130_fd_sc_hd__xor2_1
XANTENNA_153 _08762_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15593_ _05894_ _05825_ _05911_ VGND VGND VPWR VPWR _05912_ sky130_fd_sc_hd__o21a_1
X_18381_ _06330_ _06405_ _06404_ VGND VGND VPWR VPWR _08940_ sky130_fd_sc_hd__a21o_1
XANTENNA_164 _08934_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_175 _02646_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14544_ _01745_ _01139_ _04767_ VGND VGND VPWR VPWR _04769_ sky130_fd_sc_hd__a21o_1
XTAP_1773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17332_ _07797_ _03930_ _07798_ VGND VGND VPWR VPWR _07800_ sky130_fd_sc_hd__and3_2
X_11756_ _06008_ ApproximateM_inst.lob_16.lob2.genblk1\[6\].genblk1.mux.sel _03388_
+ ApproximateM_inst.lob_16.lob1.genblk1\[9\].genblk1.mux.sel VGND VGND VPWR VPWR _01849_
+ sky130_fd_sc_hd__and4_1
XTAP_1784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_624 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10707_ _05943_ _05954_ _06127_ VGND VGND VPWR VPWR _00800_ sky130_fd_sc_hd__a21o_1
XFILLER_0_153_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14475_ _04410_ _04692_ _04693_ _04551_ VGND VGND VPWR VPWR _04694_ sky130_fd_sc_hd__o2bb2a_1
X_17263_ _07018_ _07721_ _07723_ VGND VGND VPWR VPWR _07724_ sky130_fd_sc_hd__o21a_1
X_11687_ net198 _01770_ _01721_ _01739_ VGND VGND VPWR VPWR _01780_ sky130_fd_sc_hd__o211a_1
XFILLER_0_126_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_114_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19002_ clknet_4_7_0_clk _09369_ VGND VGND VPWR VPWR salida\[55\] sky130_fd_sc_hd__dfxtp_1
X_16214_ _06582_ VGND VGND VPWR VPWR _06583_ sky130_fd_sc_hd__inv_2
X_13426_ _03081_ VGND VGND VPWR VPWR _03547_ sky130_fd_sc_hd__clkbuf_4
X_10638_ _00725_ _00730_ VGND VGND VPWR VPWR _00731_ sky130_fd_sc_hd__xor2_1
XFILLER_0_3_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17194_ _00399_ _07311_ VGND VGND VPWR VPWR _07649_ sky130_fd_sc_hd__and2_2
XFILLER_0_141_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16145_ _06507_ VGND VGND VPWR VPWR _06508_ sky130_fd_sc_hd__buf_4
X_13357_ _03289_ _03268_ VGND VGND VPWR VPWR _03471_ sky130_fd_sc_hd__and2b_1
X_10569_ _00659_ _00660_ _00601_ _00602_ VGND VGND VPWR VPWR _00662_ sky130_fd_sc_hd__a211oi_2
X_12308_ _08615_ _01357_ VGND VGND VPWR VPWR _02401_ sky130_fd_sc_hd__nand2_1
X_16076_ _03169_ _06432_ VGND VGND VPWR VPWR _06433_ sky130_fd_sc_hd__and2_1
X_13288_ _03230_ _03231_ VGND VGND VPWR VPWR _03395_ sky130_fd_sc_hd__nand2_1
X_15027_ _05207_ _05176_ _05295_ VGND VGND VPWR VPWR _05296_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_20_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12239_ _07591_ _02205_ VGND VGND VPWR VPWR _02332_ sky130_fd_sc_hd__nand2_1
X_16978_ _07411_ _07412_ VGND VGND VPWR VPWR _07413_ sky130_fd_sc_hd__or2b_1
Xinput4 i_wb_addr[11] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18717_ _09209_ _09243_ VGND VGND VPWR VPWR _09244_ sky130_fd_sc_hd__and2_1
X_15929_ _06195_ _06199_ VGND VGND VPWR VPWR _06274_ sky130_fd_sc_hd__and2b_1
XFILLER_0_78_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09450_ cla_inst.in2\[19\] VGND VGND VPWR VPWR _03520_ sky130_fd_sc_hd__buf_6
X_18648_ net60 _03083_ _09193_ VGND VGND VPWR VPWR _09194_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18579_ salida\[10\] _09141_ _09142_ salida\[42\] _09128_ VGND VGND VPWR VPWR _09143_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_148_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_635 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_144_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_112_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09717_ _06406_ _06417_ VGND VGND VPWR VPWR _06428_ sky130_fd_sc_hd__and2b_1
XFILLER_0_69_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09648_ _05671_ VGND VGND VPWR VPWR _05682_ sky130_fd_sc_hd__buf_4
XTAP_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09579_ _04810_ _04821_ _04831_ VGND VGND VPWR VPWR _04930_ sky130_fd_sc_hd__a21o_1
XTAP_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11610_ _01701_ _01700_ _01602_ _01585_ VGND VGND VPWR VPWR _01703_ sky130_fd_sc_hd__o211a_1
XFILLER_0_139_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12590_ _02674_ _02681_ _02682_ VGND VGND VPWR VPWR _02683_ sky130_fd_sc_hd__and3_1
XFILLER_0_136_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11541_ _01630_ _01632_ _01631_ VGND VGND VPWR VPWR _01634_ sky130_fd_sc_hd__a21o_1
XFILLER_0_147_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_108_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14260_ _04445_ _04446_ _04456_ VGND VGND VPWR VPWR _04458_ sky130_fd_sc_hd__nor3_4
XFILLER_0_123_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11472_ _05453_ _05464_ _04154_ _00563_ VGND VGND VPWR VPWR _01565_ sky130_fd_sc_hd__nand4_2
XFILLER_0_107_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13211_ _00164_ _03311_ VGND VGND VPWR VPWR _03312_ sky130_fd_sc_hd__nand2_1
XFILLER_0_122_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10423_ _00509_ VGND VGND VPWR VPWR _00516_ sky130_fd_sc_hd__inv_4
XFILLER_0_33_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14191_ _04380_ _04381_ _04208_ _04212_ VGND VGND VPWR VPWR _04383_ sky130_fd_sc_hd__o211ai_4
X_13142_ _00620_ net136 _03237_ _03238_ VGND VGND VPWR VPWR _03240_ sky130_fd_sc_hd__o211ai_2
X_10354_ _00438_ _00445_ _00446_ VGND VGND VPWR VPWR _00447_ sky130_fd_sc_hd__nand3_1
XFILLER_0_131_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13073_ _03139_ _03148_ _03160_ _03163_ _03164_ _03081_ VGND VGND VPWR VPWR _03165_
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_130_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17950_ _07608_ _07410_ _07511_ _07195_ VGND VGND VPWR VPWR _08472_ sky130_fd_sc_hd__o22a_1
X_10285_ _09346_ _00274_ net338 _00377_ VGND VGND VPWR VPWR _00378_ sky130_fd_sc_hd__a211oi_4
X_12024_ _02030_ _02029_ VGND VGND VPWR VPWR _02117_ sky130_fd_sc_hd__and2b_1
X_16901_ _07205_ _07227_ _07203_ VGND VGND VPWR VPWR _07329_ sky130_fd_sc_hd__a21o_1
X_17881_ _08381_ _08396_ VGND VGND VPWR VPWR _08397_ sky130_fd_sc_hd__xnor2_1
X_16832_ _07250_ _07252_ _07253_ VGND VGND VPWR VPWR _07255_ sky130_fd_sc_hd__o21a_1
XFILLER_0_88_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16763_ _03094_ _06435_ VGND VGND VPWR VPWR _07180_ sky130_fd_sc_hd__nor2_1
X_13975_ _04144_ _04145_ _03963_ _03982_ VGND VGND VPWR VPWR _04147_ sky130_fd_sc_hd__o211a_1
XFILLER_0_87_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18502_ _06414_ _07084_ _09058_ _09062_ _09069_ VGND VGND VPWR VPWR _09071_ sky130_fd_sc_hd__o311a_1
X_15714_ _06041_ _06042_ VGND VGND VPWR VPWR _06043_ sky130_fd_sc_hd__or2_1
XFILLER_0_87_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12926_ _00806_ _06591_ VGND VGND VPWR VPWR _03019_ sky130_fd_sc_hd__or2_1
X_16694_ _02347_ _06871_ VGND VGND VPWR VPWR _07104_ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18433_ _06836_ _08983_ _08987_ _08996_ VGND VGND VPWR VPWR _08997_ sky130_fd_sc_hd__o211a_1
X_15645_ _05966_ _05967_ VGND VGND VPWR VPWR _05968_ sky130_fd_sc_hd__and2_1
XTAP_2260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12857_ _02948_ _02941_ _02933_ VGND VGND VPWR VPWR _02950_ sky130_fd_sc_hd__nor3_1
XTAP_2271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11808_ _01811_ _01812_ _01899_ _01900_ VGND VGND VPWR VPWR _01901_ sky130_fd_sc_hd__a211o_1
X_18364_ _08873_ _08893_ _08921_ VGND VGND VPWR VPWR _08922_ sky130_fd_sc_hd__or3_1
X_15576_ _05830_ _05843_ VGND VGND VPWR VPWR _05893_ sky130_fd_sc_hd__and2_1
XTAP_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12788_ _02879_ _02880_ VGND VGND VPWR VPWR _02881_ sky130_fd_sc_hd__and2b_2
XFILLER_0_17_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17315_ _06750_ _07780_ VGND VGND VPWR VPWR _07781_ sky130_fd_sc_hd__nand2_1
X_14527_ _04743_ _04749_ VGND VGND VPWR VPWR _04750_ sky130_fd_sc_hd__or2_1
XFILLER_0_16_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11739_ _01829_ _01830_ _01831_ VGND VGND VPWR VPWR _01832_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_126_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18295_ _08845_ _08846_ VGND VGND VPWR VPWR _08847_ sky130_fd_sc_hd__xor2_1
XFILLER_0_138_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17246_ _07590_ _07600_ VGND VGND VPWR VPWR _07705_ sky130_fd_sc_hd__nand2_1
XFILLER_0_154_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14458_ _04672_ _04673_ _04529_ _04531_ VGND VGND VPWR VPWR _04675_ sky130_fd_sc_hd__a211o_1
XFILLER_0_4_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_141_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13409_ _03525_ _03526_ _03349_ _03365_ VGND VGND VPWR VPWR _03528_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_141_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14389_ _04596_ _04597_ _04445_ net335 VGND VGND VPWR VPWR _04599_ sky130_fd_sc_hd__a211o_1
XFILLER_0_4_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17177_ _06875_ VGND VGND VPWR VPWR _07630_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_51_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16128_ _00861_ _03140_ VGND VGND VPWR VPWR _06489_ sky130_fd_sc_hd__or2_1
XFILLER_0_122_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110_833 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_122_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16059_ _06328_ _06412_ _06413_ _06248_ VGND VGND VPWR VPWR _06414_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_20_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09502_ _04078_ VGND VGND VPWR VPWR _04088_ sky130_fd_sc_hd__buf_6
XFILLER_0_154_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09433_ _03324_ _03206_ _03228_ _03292_ VGND VGND VPWR VPWR _00000_ sky130_fd_sc_hd__a22o_1
XFILLER_0_149_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_568 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_20 _01115_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_31 _01225_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_42 _02188_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_53 _03618_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_105_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_64 _04420_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_75 _06693_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_86 _08762_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_97 _08880_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_844 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_112_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10070_ cla_inst.in2\[20\] VGND VGND VPWR VPWR _00163_ sky130_fd_sc_hd__buf_4
XFILLER_0_69_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13760_ _02978_ VGND VGND VPWR VPWR _03912_ sky130_fd_sc_hd__buf_4
X_10972_ _05584_ cla_inst.in1\[16\] ApproximateM_inst.lob_16.lob1.genblk2.mux_final.sel
+ _05562_ VGND VGND VPWR VPWR _01065_ sky130_fd_sc_hd__a22o_1
XFILLER_0_58_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12711_ _02755_ _02785_ VGND VGND VPWR VPWR _02804_ sky130_fd_sc_hd__nor2_1
X_13691_ _03697_ _03698_ _03712_ VGND VGND VPWR VPWR _03836_ sky130_fd_sc_hd__a21o_1
XFILLER_0_84_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15430_ _05631_ _05641_ _05639_ VGND VGND VPWR VPWR _05734_ sky130_fd_sc_hd__a21oi_1
X_12642_ _02689_ _02734_ VGND VGND VPWR VPWR _02735_ sky130_fd_sc_hd__and2_1
X_15361_ _05577_ _05580_ _05578_ VGND VGND VPWR VPWR _05659_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_65_363 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_108_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12573_ _02656_ _02665_ VGND VGND VPWR VPWR _02666_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_26_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17100_ _07536_ _07538_ _07545_ VGND VGND VPWR VPWR _07546_ sky130_fd_sc_hd__or3_1
X_14312_ _04320_ _04322_ VGND VGND VPWR VPWR _04516_ sky130_fd_sc_hd__nor2_1
X_11524_ _01615_ _01616_ VGND VGND VPWR VPWR _01617_ sky130_fd_sc_hd__xnor2_2
X_15292_ _03000_ _03071_ _05583_ VGND VGND VPWR VPWR _05585_ sky130_fd_sc_hd__nand3_1
X_18080_ _08592_ _08596_ _08613_ _06721_ _01136_ VGND VGND VPWR VPWR _09400_ sky130_fd_sc_hd__o32a_2
XFILLER_0_123_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14243_ _02059_ _08224_ VGND VGND VPWR VPWR _04440_ sky130_fd_sc_hd__nand2_1
X_17031_ _06364_ _06545_ _07470_ _00593_ VGND VGND VPWR VPWR _07471_ sky130_fd_sc_hd__a22o_1
X_11455_ _01546_ _01547_ VGND VGND VPWR VPWR _01548_ sky130_fd_sc_hd__and2b_1
XFILLER_0_104_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10406_ _07080_ _09303_ _00498_ _07058_ VGND VGND VPWR VPWR _00499_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_21_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_68_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14174_ _09352_ _01962_ VGND VGND VPWR VPWR _04365_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11386_ _01475_ _01476_ _01478_ VGND VGND VPWR VPWR _01479_ sky130_fd_sc_hd__o21a_1
XFILLER_0_104_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13125_ _03213_ _03214_ _03220_ VGND VGND VPWR VPWR _03221_ sky130_fd_sc_hd__nand3_2
XFILLER_0_0_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10337_ _00428_ _00270_ _00427_ _00429_ VGND VGND VPWR VPWR _00430_ sky130_fd_sc_hd__a211oi_4
X_18982_ clknet_4_0_0_clk _09377_ VGND VGND VPWR VPWR salida\[35\] sky130_fd_sc_hd__dfxtp_1
XTAP_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13056_ _03147_ VGND VGND VPWR VPWR _03148_ sky130_fd_sc_hd__inv_2
X_17933_ _07751_ _07596_ _08453_ VGND VGND VPWR VPWR _08454_ sky130_fd_sc_hd__a21oi_1
X_10268_ _00357_ _00359_ _00360_ VGND VGND VPWR VPWR _00361_ sky130_fd_sc_hd__a21bo_1
X_12007_ _06765_ _02099_ _02032_ _02033_ VGND VGND VPWR VPWR _02100_ sky130_fd_sc_hd__o22a_1
X_17864_ _08277_ _08290_ _08275_ VGND VGND VPWR VPWR _08379_ sky130_fd_sc_hd__a21o_1
X_10199_ _08420_ _08463_ _08431_ VGND VGND VPWR VPWR _00292_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_108_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16815_ _06665_ _07130_ VGND VGND VPWR VPWR _07236_ sky130_fd_sc_hd__nor2_1
X_17795_ _08302_ _08303_ VGND VGND VPWR VPWR _08304_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_17_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16746_ _07158_ _07159_ _03195_ VGND VGND VPWR VPWR _07161_ sky130_fd_sc_hd__a21o_1
XFILLER_0_17_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13958_ _03952_ _03958_ VGND VGND VPWR VPWR _04128_ sky130_fd_sc_hd__or2_1
X_12909_ _02990_ _02995_ _03001_ VGND VGND VPWR VPWR _03002_ sky130_fd_sc_hd__or3_2
X_16677_ _03062_ _06724_ VGND VGND VPWR VPWR _07086_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13889_ _04050_ _04051_ _03834_ net321 VGND VGND VPWR VPWR _04053_ sky130_fd_sc_hd__a211oi_1
X_18416_ _08971_ _08976_ VGND VGND VPWR VPWR _08978_ sky130_fd_sc_hd__nor2_4
X_15628_ _05876_ _05873_ _05874_ VGND VGND VPWR VPWR _05950_ sky130_fd_sc_hd__o21ai_1
XTAP_2090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18347_ _08901_ _08902_ VGND VGND VPWR VPWR _08903_ sky130_fd_sc_hd__and2_1
X_15559_ _05873_ _05874_ VGND VGND VPWR VPWR _05875_ sky130_fd_sc_hd__or2b_1
XFILLER_0_127_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_126_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18278_ _03036_ _06148_ _06426_ _08825_ _08828_ VGND VGND VPWR VPWR _08829_ sky130_fd_sc_hd__o221a_1
XFILLER_0_127_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput40 i_wb_data[14] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__buf_2
X_17229_ _04247_ _06914_ VGND VGND VPWR VPWR _07687_ sky130_fd_sc_hd__nor2_1
XFILLER_0_142_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput51 i_wb_data[24] VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_12_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput62 i_wb_data[5] VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__buf_2
XFILLER_0_71_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_619 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_141_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09982_ _07755_ VGND VGND VPWR VPWR _09248_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_40_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_466 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_137_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_694 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_251 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_700 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11240_ _01330_ _01331_ _01313_ _01314_ VGND VGND VPWR VPWR _01333_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_15_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11171_ _00193_ VGND VGND VPWR VPWR _01264_ sky130_fd_sc_hd__buf_4
XFILLER_0_31_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10122_ _00203_ _00214_ VGND VGND VPWR VPWR _00215_ sky130_fd_sc_hd__nand2_1
XFILLER_0_100_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14930_ _05188_ _05189_ VGND VGND VPWR VPWR _05190_ sky130_fd_sc_hd__nand2_1
X_10053_ _00145_ VGND VGND VPWR VPWR _00146_ sky130_fd_sc_hd__buf_4
X_14861_ _04975_ _04982_ VGND VGND VPWR VPWR _05114_ sky130_fd_sc_hd__nand2_2
X_16600_ _06999_ _07001_ _03080_ VGND VGND VPWR VPWR _07002_ sky130_fd_sc_hd__mux2_1
X_13812_ _03790_ _03455_ VGND VGND VPWR VPWR _03969_ sky130_fd_sc_hd__nand2_1
X_17580_ _07130_ _07126_ _07195_ _07608_ VGND VGND VPWR VPWR _08069_ sky130_fd_sc_hd__or4_1
X_14792_ _00190_ _00192_ _05986_ _01223_ VGND VGND VPWR VPWR _05040_ sky130_fd_sc_hd__and4_1
X_16531_ _06344_ _06346_ _06926_ VGND VGND VPWR VPWR _06927_ sky130_fd_sc_hd__a21oi_1
X_13743_ net119 _03889_ _03891_ VGND VGND VPWR VPWR _03894_ sky130_fd_sc_hd__o21a_1
X_10955_ _01044_ _01047_ VGND VGND VPWR VPWR _01048_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_97_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16462_ _03166_ _06431_ VGND VGND VPWR VPWR _06853_ sky130_fd_sc_hd__nor2_1
XFILLER_0_128_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13674_ cla_inst.in2\[30\] cla_inst.in2\[29\] _03432_ _00205_ VGND VGND VPWR VPWR
+ _03818_ sky130_fd_sc_hd__and4_1
XFILLER_0_39_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10886_ _00967_ _00977_ _00976_ VGND VGND VPWR VPWR _00979_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_128_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18201_ _08588_ _08742_ _08743_ _08417_ _08744_ VGND VGND VPWR VPWR _08745_ sky130_fd_sc_hd__o221a_1
X_15413_ _05691_ _05690_ VGND VGND VPWR VPWR _05716_ sky130_fd_sc_hd__or2b_1
XFILLER_0_66_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12625_ _02681_ _02717_ VGND VGND VPWR VPWR _02718_ sky130_fd_sc_hd__or2_2
XFILLER_0_39_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16393_ _06583_ _06750_ _06775_ _06777_ VGND VGND VPWR VPWR _06778_ sky130_fd_sc_hd__a22o_1
XFILLER_0_81_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18132_ _08614_ _08590_ _08668_ _06516_ VGND VGND VPWR VPWR _08671_ sky130_fd_sc_hd__o31a_1
X_15344_ _05639_ _05640_ VGND VGND VPWR VPWR _05641_ sky130_fd_sc_hd__nor2_1
X_12556_ _07788_ _00878_ _02607_ VGND VGND VPWR VPWR _02649_ sky130_fd_sc_hd__a21o_1
XFILLER_0_54_878 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11507_ _01594_ _01599_ VGND VGND VPWR VPWR _01600_ sky130_fd_sc_hd__and2_1
X_18063_ _01997_ _08593_ _08595_ VGND VGND VPWR VPWR _08596_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_108_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15275_ _05556_ _05565_ VGND VGND VPWR VPWR _05566_ sky130_fd_sc_hd__xor2_1
X_12487_ _02570_ _02578_ _02521_ _02579_ VGND VGND VPWR VPWR _02580_ sky130_fd_sc_hd__a211oi_2
Xhold109 _00012_ VGND VGND VPWR VPWR net272 sky130_fd_sc_hd__dlygate4sd3_1
X_17014_ _03195_ _07451_ _07452_ VGND VGND VPWR VPWR _07453_ sky130_fd_sc_hd__or3b_2
X_14226_ _00592_ _04336_ VGND VGND VPWR VPWR _04421_ sky130_fd_sc_hd__and2_1
X_11438_ _04078_ _01151_ _01031_ _09179_ VGND VGND VPWR VPWR _01531_ sky130_fd_sc_hd__and4_1
XFILLER_0_22_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14157_ _04344_ _04345_ VGND VGND VPWR VPWR _04346_ sky130_fd_sc_hd__xnor2_1
X_11369_ _01460_ _01461_ VGND VGND VPWR VPWR _01462_ sky130_fd_sc_hd__or2_1
XTAP_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13108_ _03201_ VGND VGND VPWR VPWR _03202_ sky130_fd_sc_hd__buf_6
X_14088_ _03651_ _03662_ _00308_ _08757_ VGND VGND VPWR VPWR _04270_ sky130_fd_sc_hd__nand4_4
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18965_ clknet_4_7_0_clk _09395_ VGND VGND VPWR VPWR salida\[18\] sky130_fd_sc_hd__dfxtp_1
XTAP_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17916_ _06425_ _06444_ _08435_ VGND VGND VPWR VPWR _08436_ sky130_fd_sc_hd__or3_1
X_13039_ _00494_ _03130_ VGND VGND VPWR VPWR _03131_ sky130_fd_sc_hd__or2_1
X_18896_ clknet_4_11_0_clk _00050_ VGND VGND VPWR VPWR ApproximateM_inst.lob_16.lob1.genblk1\[14\].genblk1.mux.sel
+ sky130_fd_sc_hd__dfxtp_4
X_17847_ _07143_ _07706_ _08260_ _06961_ VGND VGND VPWR VPWR _08360_ sky130_fd_sc_hd__o22a_1
X_17778_ _08283_ _08284_ VGND VGND VPWR VPWR _08285_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_14_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_52 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16729_ _07140_ _07141_ VGND VGND VPWR VPWR _07142_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_44_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_151_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_279 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_686 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_114_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_142_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09965_ _09101_ _09112_ VGND VGND VPWR VPWR _09123_ sky130_fd_sc_hd__and2b_1
X_09896_ _08333_ _08354_ _08344_ VGND VGND VPWR VPWR _08376_ sky130_fd_sc_hd__a21o_1
XTAP_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10740_ _07036_ _07069_ cla_inst.in1\[22\] _08746_ VGND VGND VPWR VPWR _00833_ sky130_fd_sc_hd__nand4_1
XFILLER_0_138_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10671_ _03848_ _03782_ _03399_ VGND VGND VPWR VPWR _00764_ sky130_fd_sc_hd__and3_1
XFILLER_0_138_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12410_ _02436_ _02502_ VGND VGND VPWR VPWR _02503_ sky130_fd_sc_hd__nand2_1
XFILLER_0_153_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13390_ _03491_ _03492_ _03506_ VGND VGND VPWR VPWR _03507_ sky130_fd_sc_hd__a21o_2
XFILLER_0_105_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12341_ _02418_ _02432_ VGND VGND VPWR VPWR _02434_ sky130_fd_sc_hd__nand2_1
XFILLER_0_145_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15060_ _03006_ _01866_ VGND VGND VPWR VPWR _05331_ sky130_fd_sc_hd__nand2_1
XFILLER_0_50_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12272_ _02361_ _02364_ VGND VGND VPWR VPWR _02365_ sky130_fd_sc_hd__xnor2_1
X_14011_ _04174_ _04016_ _04185_ VGND VGND VPWR VPWR _04186_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_105_298 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11223_ _00862_ _01107_ VGND VGND VPWR VPWR _01316_ sky130_fd_sc_hd__and2_1
X_11154_ _01240_ _01246_ VGND VGND VPWR VPWR _01247_ sky130_fd_sc_hd__xnor2_4
X_10105_ _00195_ _00175_ _00181_ _00197_ VGND VGND VPWR VPWR _00198_ sky130_fd_sc_hd__nand4_1
X_18750_ _09269_ VGND VGND VPWR VPWR _00075_ sky130_fd_sc_hd__buf_1
X_11085_ _01166_ _01176_ _01177_ VGND VGND VPWR VPWR _01178_ sky130_fd_sc_hd__nor3_1
X_15962_ _06258_ _06284_ VGND VGND VPWR VPWR _06310_ sky130_fd_sc_hd__nor2_1
X_17701_ _08187_ _08200_ VGND VGND VPWR VPWR _08201_ sky130_fd_sc_hd__xnor2_1
X_14913_ _02999_ _03055_ _05169_ VGND VGND VPWR VPWR _05172_ sky130_fd_sc_hd__a21o_1
X_10036_ ApproximateM_inst.lob_16.lob1.genblk1\[3\].genblk1.mux.sel VGND VGND VPWR
+ VPWR _00129_ sky130_fd_sc_hd__buf_6
X_18681_ _02044_ _09190_ _09191_ VGND VGND VPWR VPWR _09218_ sky130_fd_sc_hd__a21oi_1
X_15893_ _06171_ _06214_ _06216_ VGND VGND VPWR VPWR _06236_ sky130_fd_sc_hd__a21oi_1
X_17632_ _02848_ _08125_ _03201_ VGND VGND VPWR VPWR _08127_ sky130_fd_sc_hd__o21ai_1
X_14844_ _02974_ _05095_ VGND VGND VPWR VPWR _05096_ sky130_fd_sc_hd__nor2_1
XFILLER_0_98_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17563_ _06766_ _07706_ VGND VGND VPWR VPWR _08051_ sky130_fd_sc_hd__nor2_1
X_14775_ _03322_ _03321_ _05486_ _05878_ VGND VGND VPWR VPWR _05021_ sky130_fd_sc_hd__nand4_1
XFILLER_0_98_594 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11987_ _02053_ _02078_ _02079_ VGND VGND VPWR VPWR _02080_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_14_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16514_ _08865_ _06509_ _00223_ VGND VGND VPWR VPWR _06909_ sky130_fd_sc_hd__a21boi_1
X_13726_ _03857_ _03858_ _03874_ VGND VGND VPWR VPWR _03875_ sky130_fd_sc_hd__a21oi_1
X_10938_ ApproximateM_inst.lob_16.lob1.genblk1\[2\].genblk1.mux.sel VGND VGND VPWR
+ VPWR _01031_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_105_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17494_ _07841_ _07848_ VGND VGND VPWR VPWR _07976_ sky130_fd_sc_hd__and2b_1
XFILLER_0_73_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16445_ _06775_ _06779_ _06832_ VGND VGND VPWR VPWR _06834_ sky130_fd_sc_hd__a21o_1
X_13657_ _03632_ _03634_ _03633_ VGND VGND VPWR VPWR _03799_ sky130_fd_sc_hd__a21bo_1
X_10869_ _03465_ _00171_ _00771_ _00773_ VGND VGND VPWR VPWR _00962_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_143_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12608_ _02662_ _02695_ _02700_ VGND VGND VPWR VPWR _02701_ sky130_fd_sc_hd__or3b_4
XPHY_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16376_ _04384_ _03281_ VGND VGND VPWR VPWR _06759_ sky130_fd_sc_hd__and2_1
XPHY_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13588_ _03469_ _03516_ _03722_ _03723_ VGND VGND VPWR VPWR _03724_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_27_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18115_ _08650_ _08651_ VGND VGND VPWR VPWR _08652_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15327_ _05619_ _05620_ _05622_ VGND VGND VPWR VPWR _09363_ sky130_fd_sc_hd__a21bo_1
X_12539_ _02592_ _02631_ VGND VGND VPWR VPWR _02632_ sky130_fd_sc_hd__or2_1
XFILLER_0_152_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18046_ _08482_ _08531_ _08575_ VGND VGND VPWR VPWR _08577_ sky130_fd_sc_hd__and3_1
X_15258_ _05545_ _05546_ VGND VGND VPWR VPWR _05547_ sky130_fd_sc_hd__and2_1
XFILLER_0_112_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14209_ _03742_ _04402_ VGND VGND VPWR VPWR _04403_ sky130_fd_sc_hd__nand2_1
XFILLER_0_112_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15189_ _05463_ _05471_ VGND VGND VPWR VPWR _05472_ sky130_fd_sc_hd__xor2_1
XFILLER_0_111_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09750_ _06754_ _06700_ _06765_ _06776_ VGND VGND VPWR VPWR _06787_ sky130_fd_sc_hd__o2bb2a_1
X_18948_ clknet_4_5_0_clk _09397_ VGND VGND VPWR VPWR salida\[1\] sky130_fd_sc_hd__dfxtp_2
X_09681_ _06029_ VGND VGND VPWR VPWR _06040_ sky130_fd_sc_hd__buf_4
X_18879_ clknet_4_15_0_clk net247 VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_119_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_130_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09948_ _08692_ _08702_ _08919_ VGND VGND VPWR VPWR _08941_ sky130_fd_sc_hd__nand3_2
X_09879_ _07700_ _08158_ _08180_ VGND VGND VPWR VPWR _08191_ sky130_fd_sc_hd__and3_1
X_11910_ _02001_ _02002_ VGND VGND VPWR VPWR _02003_ sky130_fd_sc_hd__nor2_1
XFILLER_0_99_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12890_ _02982_ VGND VGND VPWR VPWR _02983_ sky130_fd_sc_hd__clkbuf_4
XTAP_2601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11841_ _01908_ _01912_ VGND VGND VPWR VPWR _01934_ sky130_fd_sc_hd__or2b_1
XTAP_2634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14560_ _04784_ _04785_ VGND VGND VPWR VPWR _04786_ sky130_fd_sc_hd__xnor2_1
X_11772_ _01675_ _01864_ VGND VGND VPWR VPWR _01865_ sky130_fd_sc_hd__and2_1
XTAP_2678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13511_ _03630_ _03637_ _03638_ VGND VGND VPWR VPWR _03639_ sky130_fd_sc_hd__nand3_1
X_10723_ _00811_ _00815_ VGND VGND VPWR VPWR _00816_ sky130_fd_sc_hd__and2_1
XTAP_1977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14491_ _01521_ _07156_ _04707_ _04708_ VGND VGND VPWR VPWR _04710_ sky130_fd_sc_hd__a22o_1
XFILLER_0_82_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_748 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16230_ _01746_ _06595_ _06596_ _06599_ VGND VGND VPWR VPWR _06600_ sky130_fd_sc_hd__o2bb2a_1
X_10654_ _00537_ _00600_ _00745_ _00746_ VGND VGND VPWR VPWR _00747_ sky130_fd_sc_hd__o211a_2
X_13442_ _02979_ _03562_ VGND VGND VPWR VPWR _03564_ sky130_fd_sc_hd__nor2_1
XFILLER_0_153_658 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13373_ _01873_ _03107_ VGND VGND VPWR VPWR _03489_ sky130_fd_sc_hd__nand2_1
X_16161_ _06051_ _05682_ _07047_ _06524_ VGND VGND VPWR VPWR _06525_ sky130_fd_sc_hd__or4_4
XFILLER_0_91_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10585_ _09172_ VGND VGND VPWR VPWR _00678_ sky130_fd_sc_hd__buf_2
XFILLER_0_50_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15112_ _05260_ _05283_ _05386_ VGND VGND VPWR VPWR _05389_ sky130_fd_sc_hd__and3_1
XFILLER_0_2_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12324_ _02414_ _02415_ VGND VGND VPWR VPWR _02417_ sky130_fd_sc_hd__xor2_1
XFILLER_0_51_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16092_ _03073_ _06408_ _06449_ VGND VGND VPWR VPWR _06451_ sky130_fd_sc_hd__and3_1
XFILLER_0_32_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15043_ _05210_ _05218_ VGND VGND VPWR VPWR _05313_ sky130_fd_sc_hd__or2b_1
XFILLER_0_50_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12255_ _08615_ _01746_ _01357_ _02347_ VGND VGND VPWR VPWR _02348_ sky130_fd_sc_hd__a22o_1
X_11206_ _01297_ _01298_ VGND VGND VPWR VPWR _01299_ sky130_fd_sc_hd__xor2_1
XFILLER_0_121_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12186_ _02254_ _02264_ _02277_ _02278_ VGND VGND VPWR VPWR _02279_ sky130_fd_sc_hd__a211oi_2
X_11137_ _01138_ _01140_ _01141_ _01135_ _01134_ VGND VGND VPWR VPWR _01230_ sky130_fd_sc_hd__a32o_1
X_18802_ _09310_ VGND VGND VPWR VPWR _00091_ sky130_fd_sc_hd__clkbuf_1
X_16994_ _07427_ _07429_ _07407_ VGND VGND VPWR VPWR _07431_ sky130_fd_sc_hd__a21oi_1
X_18733_ _03077_ net57 _09251_ VGND VGND VPWR VPWR _09257_ sky130_fd_sc_hd__mux2_1
X_11068_ _03509_ _00871_ _07581_ _03345_ VGND VGND VPWR VPWR _01161_ sky130_fd_sc_hd__a22o_1
X_15945_ _03911_ _03926_ _03912_ VGND VGND VPWR VPWR _06292_ sky130_fd_sc_hd__mux2_1
X_10019_ _00109_ VGND VGND VPWR VPWR _00112_ sky130_fd_sc_hd__clkbuf_4
X_18664_ _09176_ _09206_ VGND VGND VPWR VPWR _09207_ sky130_fd_sc_hd__and2_1
XFILLER_0_116_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15876_ _06216_ _06217_ VGND VGND VPWR VPWR _06218_ sky130_fd_sc_hd__nor2_1
X_17615_ _08106_ _08107_ VGND VGND VPWR VPWR _08108_ sky130_fd_sc_hd__nor2_1
XFILLER_0_149_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14827_ _04942_ _04945_ VGND VGND VPWR VPWR _05078_ sky130_fd_sc_hd__or2_1
XFILLER_0_116_56 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18595_ salida\[17\] _09141_ _09142_ salida\[49\] _09146_ VGND VGND VPWR VPWR _09154_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_86_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17546_ _03693_ _06441_ _08032_ VGND VGND VPWR VPWR _08033_ sky130_fd_sc_hd__o21a_1
X_14758_ _00679_ _00678_ _04591_ _01005_ VGND VGND VPWR VPWR _05002_ sky130_fd_sc_hd__and4_1
XFILLER_0_128_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13709_ _03854_ _03855_ VGND VGND VPWR VPWR _03856_ sky130_fd_sc_hd__or2_1
XFILLER_0_58_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17477_ _07130_ _07195_ _07608_ _07042_ VGND VGND VPWR VPWR _07957_ sky130_fd_sc_hd__o22a_1
X_14689_ _04924_ _04925_ _04794_ _04796_ VGND VGND VPWR VPWR _04927_ sky130_fd_sc_hd__a211o_1
XFILLER_0_46_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_129_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16428_ _06811_ _06814_ _00181_ VGND VGND VPWR VPWR _06815_ sky130_fd_sc_hd__or3b_1
XFILLER_0_117_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_143_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16359_ _00881_ _03094_ _00167_ _03101_ _06477_ _03161_ VGND VGND VPWR VPWR _06740_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_14_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18029_ _08556_ _08557_ VGND VGND VPWR VPWR _08558_ sky130_fd_sc_hd__and2_1
X_09802_ ApproximateM_inst.lob_16.lob2.genblk1\[2\].genblk1.mux.sel VGND VGND VPWR
+ VPWR _07352_ sky130_fd_sc_hd__buf_4
X_09733_ _05399_ _06591_ cla_inst.in1\[20\] net233 VGND VGND VPWR VPWR _06602_ sky130_fd_sc_hd__and4_1
X_09664_ _05845_ VGND VGND VPWR VPWR _05856_ sky130_fd_sc_hd__buf_4
X_09595_ _05061_ _05093_ VGND VGND VPWR VPWR _05104_ sky130_fd_sc_hd__xnor2_2
XTAP_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_135_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_134_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_150_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10370_ _00458_ _00462_ VGND VGND VPWR VPWR _00463_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_143_680 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12040_ _02050_ _02106_ _02105_ _02090_ VGND VGND VPWR VPWR _02133_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_130_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13991_ _04148_ _04163_ VGND VGND VPWR VPWR _04164_ sky130_fd_sc_hd__xnor2_1
X_15730_ _06058_ _06059_ VGND VGND VPWR VPWR _06060_ sky130_fd_sc_hd__nand2_1
X_12942_ _02979_ _03034_ VGND VGND VPWR VPWR _03035_ sky130_fd_sc_hd__or2_4
XFILLER_0_99_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15661_ _05903_ _05905_ _05984_ VGND VGND VPWR VPWR _05985_ sky130_fd_sc_hd__o21a_1
XTAP_2420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_110 net42 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12873_ _03239_ _03217_ VGND VGND VPWR VPWR _02966_ sky130_fd_sc_hd__or2_1
XTAP_2431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_121 _02476_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_132 _04191_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17400_ _07871_ _07872_ VGND VGND VPWR VPWR _07873_ sky130_fd_sc_hd__xnor2_1
X_14612_ _04839_ _04840_ _04835_ _04836_ VGND VGND VPWR VPWR _04843_ sky130_fd_sc_hd__a211o_1
XANTENNA_143 _08180_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11824_ _01913_ _01916_ VGND VGND VPWR VPWR _01917_ sky130_fd_sc_hd__and2b_1
X_18380_ _03120_ _06229_ _08938_ VGND VGND VPWR VPWR _08939_ sky130_fd_sc_hd__o21a_1
XTAP_2464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15592_ _05908_ _05909_ VGND VGND VPWR VPWR _05911_ sky130_fd_sc_hd__xnor2_1
XTAP_1730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_154 _08762_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_165 _09380_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_176 _02646_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17331_ _02589_ _02844_ VGND VGND VPWR VPWR _07798_ sky130_fd_sc_hd__nand2_1
XTAP_2497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14543_ _01745_ _01139_ _04767_ VGND VGND VPWR VPWR _04768_ sky130_fd_sc_hd__nand3_2
XFILLER_0_68_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11755_ _07363_ _01575_ _01846_ _01847_ VGND VGND VPWR VPWR _01848_ sky130_fd_sc_hd__a31o_2
XTAP_1774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_247 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10706_ _00798_ _00791_ _00784_ VGND VGND VPWR VPWR _00799_ sky130_fd_sc_hd__a21o_1
XFILLER_0_71_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17262_ _06969_ _07394_ _07396_ _06891_ VGND VGND VPWR VPWR _07723_ sky130_fd_sc_hd__a22o_1
X_14474_ _04399_ _04400_ _04549_ VGND VGND VPWR VPWR _04693_ sky130_fd_sc_hd__o21a_1
XFILLER_0_126_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11686_ _01748_ _01778_ VGND VGND VPWR VPWR _01779_ sky130_fd_sc_hd__xor2_1
XFILLER_0_125_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19001_ clknet_4_7_0_clk _09368_ VGND VGND VPWR VPWR salida\[54\] sky130_fd_sc_hd__dfxtp_1
X_16213_ _06561_ _06563_ _06572_ _06581_ VGND VGND VPWR VPWR _06582_ sky130_fd_sc_hd__or4_2
XFILLER_0_126_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13425_ _03164_ _03545_ VGND VGND VPWR VPWR _03546_ sky130_fd_sc_hd__nor2_1
XFILLER_0_36_483 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10637_ _00728_ _00729_ VGND VGND VPWR VPWR _00730_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_11_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17193_ _07645_ _07647_ VGND VGND VPWR VPWR _07648_ sky130_fd_sc_hd__or2b_1
XFILLER_0_23_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16144_ _03239_ _06418_ VGND VGND VPWR VPWR _06507_ sky130_fd_sc_hd__nor2_1
X_10568_ _00601_ _00602_ _00659_ _00660_ VGND VGND VPWR VPWR _00661_ sky130_fd_sc_hd__o211a_2
X_13356_ _03467_ _03468_ net131 _03373_ VGND VGND VPWR VPWR _03470_ sky130_fd_sc_hd__a211o_1
XFILLER_0_24_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12307_ _02395_ _02399_ VGND VGND VPWR VPWR _02400_ sky130_fd_sc_hd__or2_1
X_16075_ _03086_ _01264_ _06431_ VGND VGND VPWR VPWR _06432_ sky130_fd_sc_hd__and3_1
X_13287_ _03390_ _03391_ _03392_ VGND VGND VPWR VPWR _03394_ sky130_fd_sc_hd__a21oi_1
X_10499_ _00591_ VGND VGND VPWR VPWR _00592_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_121_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15026_ _05292_ _05294_ VGND VGND VPWR VPWR _05295_ sky130_fd_sc_hd__xor2_2
X_12238_ _08724_ _00132_ _02206_ _02207_ VGND VGND VPWR VPWR _02331_ sky130_fd_sc_hd__a22oi_2
X_12169_ _00846_ _00557_ _02257_ VGND VGND VPWR VPWR _02262_ sky130_fd_sc_hd__a21oi_2
X_16977_ net237 _06951_ _07035_ _07410_ VGND VGND VPWR VPWR _07412_ sky130_fd_sc_hd__or4_1
Xinput5 i_wb_addr[12] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_127_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18716_ net56 _03073_ _09182_ VGND VGND VPWR VPWR _09243_ sky130_fd_sc_hd__mux2_1
X_15928_ _06237_ _06208_ _06240_ VGND VGND VPWR VPWR _06273_ sky130_fd_sc_hd__a21o_1
X_18647_ _09182_ VGND VGND VPWR VPWR _09193_ sky130_fd_sc_hd__clkbuf_4
X_15859_ _03007_ _03149_ _06198_ VGND VGND VPWR VPWR _06199_ sky130_fd_sc_hd__and3_1
X_18578_ _09117_ VGND VGND VPWR VPWR _09142_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_93_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17529_ _07931_ _07932_ _08013_ VGND VGND VPWR VPWR _08014_ sky130_fd_sc_hd__o21ba_2
XFILLER_0_74_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_117_647 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_144_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_472 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_280 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_144_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09716_ _04362_ _05028_ _04569_ _04635_ VGND VGND VPWR VPWR _06417_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09647_ ApproximateM_inst.lob_16.lob2.genblk1\[5\].genblk1.mux.sel VGND VGND VPWR
+ VPWR _05671_ sky130_fd_sc_hd__buf_4
XTAP_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09578_ _04853_ _04908_ VGND VGND VPWR VPWR _04919_ sky130_fd_sc_hd__xnor2_2
XTAP_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11540_ _01630_ _01631_ _01632_ VGND VGND VPWR VPWR _01633_ sky130_fd_sc_hd__nand3_2
XFILLER_0_25_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_147_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_386 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_108_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11471_ _01525_ _01540_ _01562_ _01563_ VGND VGND VPWR VPWR _01564_ sky130_fd_sc_hd__a211o_2
XFILLER_0_151_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_751 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13210_ _02124_ VGND VGND VPWR VPWR _03311_ sky130_fd_sc_hd__buf_4
X_10422_ _00514_ VGND VGND VPWR VPWR _00515_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_150_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14190_ _04208_ _04212_ _04380_ _04381_ VGND VGND VPWR VPWR _04382_ sky130_fd_sc_hd__a211o_2
XFILLER_0_60_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10353_ _00435_ _00436_ _00437_ VGND VGND VPWR VPWR _00446_ sky130_fd_sc_hd__a21o_1
X_13141_ _03224_ _03225_ _03236_ VGND VGND VPWR VPWR _03238_ sky130_fd_sc_hd__or3_1
XFILLER_0_103_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13072_ _03062_ VGND VGND VPWR VPWR _03164_ sky130_fd_sc_hd__clkbuf_4
X_10284_ _00372_ _00373_ _00376_ _00336_ VGND VGND VPWR VPWR _00377_ sky130_fd_sc_hd__o2bb2a_1
X_12023_ _00832_ _03815_ VGND VGND VPWR VPWR _02116_ sky130_fd_sc_hd__nand2_1
X_16900_ _07300_ _07327_ VGND VGND VPWR VPWR _07328_ sky130_fd_sc_hd__xnor2_1
X_17880_ _08394_ _08395_ VGND VGND VPWR VPWR _08396_ sky130_fd_sc_hd__nor2_1
X_16831_ _07250_ _07252_ _06559_ VGND VGND VPWR VPWR _07253_ sky130_fd_sc_hd__a21oi_1
X_16762_ _03094_ _06435_ VGND VGND VPWR VPWR _07179_ sky130_fd_sc_hd__and2_1
X_13974_ _03963_ _03982_ _04144_ _04145_ VGND VGND VPWR VPWR _04146_ sky130_fd_sc_hd__a211oi_2
X_18501_ _06426_ _06452_ _09063_ _09068_ VGND VGND VPWR VPWR _09069_ sky130_fd_sc_hd__o31a_1
X_15713_ _01359_ _04125_ _06038_ _06039_ VGND VGND VPWR VPWR _06042_ sky130_fd_sc_hd__a22oi_1
X_12925_ ApproximateM_inst.lob_16.lob2.genblk1\[8\].genblk1.mux.sel _06008_ VGND VGND
+ VPWR VPWR _03018_ sky130_fd_sc_hd__or2_1
X_16693_ _07019_ _07046_ VGND VGND VPWR VPWR _07103_ sky130_fd_sc_hd__nor2_1
XFILLER_0_87_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18432_ _06410_ _07084_ _08988_ _08990_ _08994_ VGND VGND VPWR VPWR _08996_ sky130_fd_sc_hd__o311a_1
X_15644_ _05958_ _05965_ VGND VGND VPWR VPWR _05967_ sky130_fd_sc_hd__nand2_1
XTAP_2250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12856_ _02941_ _02933_ _02948_ VGND VGND VPWR VPWR _02949_ sky130_fd_sc_hd__o21a_1
XFILLER_0_69_873 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11807_ _01897_ VGND VGND VPWR VPWR _01900_ sky130_fd_sc_hd__inv_2
XTAP_2294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18363_ _08917_ _08920_ VGND VGND VPWR VPWR _08921_ sky130_fd_sc_hd__xnor2_1
X_15575_ _05890_ _05891_ VGND VGND VPWR VPWR _05892_ sky130_fd_sc_hd__and2_1
XTAP_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12787_ _02863_ _02872_ _02878_ VGND VGND VPWR VPWR _02880_ sky130_fd_sc_hd__a21o_1
XFILLER_0_22_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17314_ _02259_ _06814_ VGND VGND VPWR VPWR _07780_ sky130_fd_sc_hd__nor2_4
XFILLER_0_139_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14526_ _04747_ _04748_ VGND VGND VPWR VPWR _04749_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_56_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11738_ _05279_ _05355_ _03607_ _00217_ VGND VGND VPWR VPWR _01831_ sky130_fd_sc_hd__nand4_2
XFILLER_0_113_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18294_ _03107_ _07390_ VGND VGND VPWR VPWR _08846_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17245_ _07603_ _07615_ VGND VGND VPWR VPWR _07704_ sky130_fd_sc_hd__nor2_1
X_14457_ _04529_ _04531_ _04672_ _04673_ VGND VGND VPWR VPWR _04674_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_114_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11669_ _01217_ _01219_ _01227_ VGND VGND VPWR VPWR _01762_ sky130_fd_sc_hd__o21a_1
XFILLER_0_154_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13408_ _03349_ _03365_ _03525_ _03526_ VGND VGND VPWR VPWR _03527_ sky130_fd_sc_hd__a211o_1
XFILLER_0_113_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17176_ _07627_ _07628_ VGND VGND VPWR VPWR _07629_ sky130_fd_sc_hd__or2_1
X_14388_ _04445_ net335 _04596_ _04597_ VGND VGND VPWR VPWR _04598_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_40_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16127_ _03152_ _06485_ _06486_ _06487_ VGND VGND VPWR VPWR _06488_ sky130_fd_sc_hd__a211o_1
XFILLER_0_24_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13339_ _03279_ _03285_ VGND VGND VPWR VPWR _03451_ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16058_ _03011_ _03155_ VGND VGND VPWR VPWR _06413_ sky130_fd_sc_hd__nor2_1
XFILLER_0_110_845 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15009_ _05263_ _05171_ _05275_ VGND VGND VPWR VPWR _05276_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_44_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09501_ cla_inst.in2\[16\] VGND VGND VPWR VPWR _04078_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_514 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09432_ _03313_ VGND VGND VPWR VPWR _03324_ sky130_fd_sc_hd__buf_4
XFILLER_0_2_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_10 _00516_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_21 _01115_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_32 _01266_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_43 _02200_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_54 _03618_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_65 _04537_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_76 _06799_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_87 _08820_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_98 _08880_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_856 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10971_ _05562_ _05584_ ApproximateM_inst.lob_16.lob1.genblk2.mux_final.sel VGND
+ VGND VPWR VPWR _01064_ sky130_fd_sc_hd__and3_1
X_12710_ _02794_ _02802_ VGND VGND VPWR VPWR _02803_ sky130_fd_sc_hd__or2_1
XFILLER_0_69_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13690_ _03832_ _03833_ _03649_ _03751_ VGND VGND VPWR VPWR _03835_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_57_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12641_ _02691_ _02711_ _02726_ VGND VGND VPWR VPWR _02734_ sky130_fd_sc_hd__and3_1
XFILLER_0_84_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15360_ _05656_ _05657_ VGND VGND VPWR VPWR _05658_ sky130_fd_sc_hd__xnor2_1
X_12572_ _02658_ _02663_ _02664_ VGND VGND VPWR VPWR _02665_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_38_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14311_ _01356_ _01962_ _04364_ _04363_ VGND VGND VPWR VPWR _04514_ sky130_fd_sc_hd__a31o_1
XFILLER_0_92_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11523_ _01541_ _01543_ VGND VGND VPWR VPWR _01616_ sky130_fd_sc_hd__nand2_1
XFILLER_0_81_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15291_ _05581_ _05582_ VGND VGND VPWR VPWR _05583_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_108_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17030_ _08615_ _06592_ _06551_ VGND VGND VPWR VPWR _07470_ sky130_fd_sc_hd__a21o_1
X_14242_ _04436_ _04437_ VGND VGND VPWR VPWR _04439_ sky130_fd_sc_hd__nor2_1
XFILLER_0_135_285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11454_ _01543_ _01545_ _01544_ VGND VGND VPWR VPWR _01547_ sky130_fd_sc_hd__a21o_1
XFILLER_0_22_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10405_ cla_inst.in1\[28\] VGND VGND VPWR VPWR _00498_ sky130_fd_sc_hd__buf_2
XFILLER_0_123_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14173_ _04361_ _04363_ VGND VGND VPWR VPWR _04364_ sky130_fd_sc_hd__nor2_1
X_11385_ _01477_ _00879_ VGND VGND VPWR VPWR _01478_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_21_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13124_ _03218_ _03219_ VGND VGND VPWR VPWR _03220_ sky130_fd_sc_hd__xor2_2
X_10336_ _00424_ _00426_ _09348_ _00273_ VGND VGND VPWR VPWR _00429_ sky130_fd_sc_hd__o211a_1
X_18981_ clknet_4_1_0_clk _09366_ VGND VGND VPWR VPWR salida\[34\] sky130_fd_sc_hd__dfxtp_1
XTAP_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_9_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_9_0_clk sky130_fd_sc_hd__clkbuf_8
XTAP_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10267_ _07504_ _00127_ _07559_ _00358_ VGND VGND VPWR VPWR _00360_ sky130_fd_sc_hd__a22o_1
X_13055_ _03141_ _03146_ _03049_ VGND VGND VPWR VPWR _03147_ sky130_fd_sc_hd__mux2_1
X_17932_ _07218_ _07486_ VGND VGND VPWR VPWR _08453_ sky130_fd_sc_hd__nor2_1
X_12006_ _00563_ VGND VGND VPWR VPWR _02099_ sky130_fd_sc_hd__inv_4
X_17863_ _08366_ _08377_ VGND VGND VPWR VPWR _08378_ sky130_fd_sc_hd__xor2_1
X_10198_ _00288_ _00289_ _00290_ VGND VGND VPWR VPWR _00291_ sky130_fd_sc_hd__and3_2
XFILLER_0_17_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16814_ _07233_ _07234_ VGND VGND VPWR VPWR _07235_ sky130_fd_sc_hd__xor2_1
X_17794_ _07630_ _07741_ VGND VGND VPWR VPWR _08303_ sky130_fd_sc_hd__nor2_1
X_16745_ _07158_ _07159_ VGND VGND VPWR VPWR _07160_ sky130_fd_sc_hd__nor2_1
X_13957_ _03974_ _03975_ _04126_ VGND VGND VPWR VPWR _04127_ sky130_fd_sc_hd__a21o_1
X_12908_ _02997_ _02998_ _03000_ _00591_ VGND VGND VPWR VPWR _03001_ sky130_fd_sc_hd__or4_1
X_16676_ _06343_ _06342_ _06997_ _07084_ VGND VGND VPWR VPWR _07085_ sky130_fd_sc_hd__a31o_1
X_13888_ _03834_ net321 _04050_ _04051_ VGND VGND VPWR VPWR _04052_ sky130_fd_sc_hd__o211a_1
XFILLER_0_124_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15627_ _05948_ _05875_ VGND VGND VPWR VPWR _05949_ sky130_fd_sc_hd__nor2_1
X_18415_ _08971_ _08976_ VGND VGND VPWR VPWR _08977_ sky130_fd_sc_hd__and2_1
XFILLER_0_33_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12839_ _02930_ _02931_ VGND VGND VPWR VPWR _02932_ sky130_fd_sc_hd__xnor2_2
XTAP_2080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_651 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18346_ _04537_ _07743_ _08900_ VGND VGND VPWR VPWR _08902_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_139_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15558_ _05870_ _05871_ _05872_ VGND VGND VPWR VPWR _05874_ sky130_fd_sc_hd__o21ai_1
XTAP_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14509_ _04576_ _04577_ _04729_ VGND VGND VPWR VPWR _04730_ sky130_fd_sc_hd__o21ai_4
X_18277_ _07269_ _08141_ _08827_ _06721_ VGND VGND VPWR VPWR _08828_ sky130_fd_sc_hd__o211a_1
XFILLER_0_115_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_154_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15489_ _02973_ _03564_ VGND VGND VPWR VPWR _05799_ sky130_fd_sc_hd__nand2_1
XFILLER_0_127_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17228_ _06639_ _06627_ _02981_ VGND VGND VPWR VPWR _07686_ sky130_fd_sc_hd__mux2_1
Xinput30 i_wb_addr[6] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__clkbuf_1
Xinput41 i_wb_data[15] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__buf_2
XFILLER_0_4_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput52 i_wb_data[25] VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__buf_1
XFILLER_0_71_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput63 i_wb_data[6] VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__buf_2
XFILLER_0_52_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_678 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17159_ _06764_ _07018_ _07194_ _07608_ VGND VGND VPWR VPWR _07610_ sky130_fd_sc_hd__or4_1
XFILLER_0_40_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09981_ _09226_ _09232_ VGND VGND VPWR VPWR _09240_ sky130_fd_sc_hd__or2_2
XFILLER_0_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_478 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_364 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_712 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_879 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11170_ _01261_ _01262_ VGND VGND VPWR VPWR _01263_ sky130_fd_sc_hd__nor2_2
XFILLER_0_113_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10121_ _00213_ VGND VGND VPWR VPWR _00214_ sky130_fd_sc_hd__buf_4
XFILLER_0_100_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10052_ ApproximateM_inst.lob_16.lob1.genblk1\[4\].genblk1.mux.sel VGND VGND VPWR
+ VPWR _00145_ sky130_fd_sc_hd__clkbuf_4
X_14860_ _05109_ _05112_ VGND VGND VPWR VPWR _05113_ sky130_fd_sc_hd__xnor2_1
X_13811_ _03774_ net171 _03966_ VGND VGND VPWR VPWR _03967_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_98_732 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14791_ _02996_ _01139_ _01223_ _02993_ VGND VGND VPWR VPWR _05038_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_97_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16530_ _06338_ _06348_ _06349_ VGND VGND VPWR VPWR _06926_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_97_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13742_ net119 _03889_ _03891_ VGND VGND VPWR VPWR _03893_ sky130_fd_sc_hd__nor3_1
XFILLER_0_98_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10954_ _06460_ _04067_ _01045_ _01046_ VGND VGND VPWR VPWR _01047_ sky130_fd_sc_hd__a31o_1
XFILLER_0_97_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16461_ _03166_ _03083_ _06430_ VGND VGND VPWR VPWR _06851_ sky130_fd_sc_hd__and3_1
X_13673_ cla_inst.in2\[31\] _00172_ VGND VGND VPWR VPWR _03817_ sky130_fd_sc_hd__nand2_1
X_10885_ _00967_ _00976_ _00977_ VGND VGND VPWR VPWR _00978_ sky130_fd_sc_hd__or3_1
XFILLER_0_66_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18200_ _08582_ _08614_ _08667_ VGND VGND VPWR VPWR _08744_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_39_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15412_ _03548_ _05623_ _05625_ _03125_ _05714_ VGND VGND VPWR VPWR _09364_ sky130_fd_sc_hd__a221o_1
XFILLER_0_128_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12624_ _02675_ _02680_ _02679_ VGND VGND VPWR VPWR _02717_ sky130_fd_sc_hd__a21oi_1
X_16392_ _06659_ _06668_ _06774_ VGND VGND VPWR VPWR _06777_ sky130_fd_sc_hd__a21o_1
XFILLER_0_109_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18131_ _08614_ _08590_ _08668_ VGND VGND VPWR VPWR _08669_ sky130_fd_sc_hd__o21ai_1
X_15343_ _05636_ _05637_ _05632_ VGND VGND VPWR VPWR _05640_ sky130_fd_sc_hd__a21oi_1
X_12555_ _02608_ _02647_ VGND VGND VPWR VPWR _02648_ sky130_fd_sc_hd__nand2_1
XFILLER_0_81_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11506_ _01595_ _01598_ VGND VGND VPWR VPWR _01599_ sky130_fd_sc_hd__xor2_2
X_18062_ _01997_ _08593_ _03930_ VGND VGND VPWR VPWR _08595_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_123_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15274_ _05563_ _05564_ VGND VGND VPWR VPWR _05565_ sky130_fd_sc_hd__nor2_1
X_12486_ _02515_ _02520_ _02519_ VGND VGND VPWR VPWR _02579_ sky130_fd_sc_hd__o21a_1
XFILLER_0_123_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17013_ _07345_ _07349_ _07449_ VGND VGND VPWR VPWR _07452_ sky130_fd_sc_hd__or3_1
X_14225_ _04390_ _04391_ _04392_ VGND VGND VPWR VPWR _04420_ sky130_fd_sc_hd__or3_4
X_11437_ ApproximateM_inst.lob_16.lob2.genblk1\[11\].genblk1.mux.sel _03618_ _01527_
+ _01528_ VGND VGND VPWR VPWR _01530_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14156_ _04175_ _04179_ _04177_ VGND VGND VPWR VPWR _04345_ sky130_fd_sc_hd__o21ba_1
X_11368_ _01458_ _01459_ _01455_ _01456_ VGND VGND VPWR VPWR _01461_ sky130_fd_sc_hd__o211a_1
XTAP_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13107_ _03200_ VGND VGND VPWR VPWR _03201_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_0_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10319_ _00401_ _00402_ _00411_ VGND VGND VPWR VPWR _00412_ sky130_fd_sc_hd__o21a_1
X_14087_ _03662_ _05704_ _08757_ _03629_ VGND VGND VPWR VPWR _04269_ sky130_fd_sc_hd__a22o_1
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18964_ clknet_4_7_0_clk _09394_ VGND VGND VPWR VPWR salida\[17\] sky130_fd_sc_hd__dfxtp_1
XTAP_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11299_ _01382_ _01389_ _01390_ _01391_ VGND VGND VPWR VPWR _01392_ sky130_fd_sc_hd__nand4_4
XTAP_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17915_ _03041_ _06443_ _04336_ VGND VGND VPWR VPWR _08435_ sky130_fd_sc_hd__a21oi_1
X_13038_ _03127_ _03129_ _03048_ VGND VGND VPWR VPWR _03130_ sky130_fd_sc_hd__mux2_1
X_18895_ clknet_4_11_0_clk _00049_ VGND VGND VPWR VPWR ApproximateM_inst.lob_16.lob1.genblk1\[13\].genblk1.mux.sel
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_28_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17846_ _07143_ _08262_ VGND VGND VPWR VPWR _08359_ sky130_fd_sc_hd__and2_1
XFILLER_0_89_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14989_ _05248_ _05253_ VGND VGND VPWR VPWR _05254_ sky130_fd_sc_hd__xnor2_1
X_17777_ _07109_ _07649_ VGND VGND VPWR VPWR _08284_ sky130_fd_sc_hd__nand2_1
XFILLER_0_135_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16728_ _07040_ _07043_ _07037_ VGND VGND VPWR VPWR _07141_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_44_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16659_ _07063_ _07065_ VGND VGND VPWR VPWR _07066_ sky130_fd_sc_hd__and2b_1
XFILLER_0_76_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_146_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18329_ _06403_ _06546_ _08883_ _03143_ VGND VGND VPWR VPWR _08884_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_115_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_562 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09964_ _07080_ _07374_ _07406_ _07047_ VGND VGND VPWR VPWR _09112_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09895_ _08333_ _08344_ _08354_ VGND VGND VPWR VPWR _08365_ sky130_fd_sc_hd__nand3_1
XTAP_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_149_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10670_ _04296_ _04285_ _04187_ VGND VGND VPWR VPWR _00763_ sky130_fd_sc_hd__a21o_1
XFILLER_0_63_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_643 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12340_ _02418_ _02432_ VGND VGND VPWR VPWR _02433_ sky130_fd_sc_hd__or2_1
XFILLER_0_106_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12271_ _02362_ _02363_ VGND VGND VPWR VPWR _02364_ sky130_fd_sc_hd__xnor2_1
X_14010_ _04183_ _04184_ VGND VGND VPWR VPWR _04185_ sky130_fd_sc_hd__nand2_1
X_11222_ _00862_ _01107_ VGND VGND VPWR VPWR _01315_ sky130_fd_sc_hd__nor2_1
XFILLER_0_31_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11153_ _01243_ _01245_ VGND VGND VPWR VPWR _01246_ sky130_fd_sc_hd__nor2_2
X_10104_ _00196_ VGND VGND VPWR VPWR _00197_ sky130_fd_sc_hd__buf_4
X_11084_ _01149_ _01150_ _01165_ VGND VGND VPWR VPWR _01177_ sky130_fd_sc_hd__a21oi_2
X_15961_ _06306_ _06307_ VGND VGND VPWR VPWR _06308_ sky130_fd_sc_hd__and2_1
X_17700_ _08198_ _08199_ VGND VGND VPWR VPWR _08200_ sky130_fd_sc_hd__nor2_1
X_14912_ _02999_ _03055_ _05169_ VGND VGND VPWR VPWR _05171_ sky130_fd_sc_hd__nand3_1
X_10035_ _00125_ _00127_ _09188_ _00109_ VGND VGND VPWR VPWR _00128_ sky130_fd_sc_hd__a22o_1
X_18680_ net40 _09189_ _09217_ VGND VGND VPWR VPWR _00050_ sky130_fd_sc_hd__o21a_1
X_15892_ _06190_ _06225_ _06231_ _06184_ _06233_ VGND VGND VPWR VPWR _06235_ sky130_fd_sc_hd__o221a_1
X_14843_ _03912_ _04082_ _05094_ VGND VGND VPWR VPWR _05095_ sky130_fd_sc_hd__o21ai_1
X_17631_ _02846_ _02847_ _02465_ VGND VGND VPWR VPWR _08125_ sky130_fd_sc_hd__a21bo_1
X_17562_ _08045_ _08046_ _08048_ VGND VGND VPWR VPWR _08050_ sky130_fd_sc_hd__a21o_1
X_14774_ _09350_ _05486_ _05878_ _00112_ VGND VGND VPWR VPWR _05020_ sky130_fd_sc_hd__a22o_1
X_11986_ _02073_ _02077_ _01984_ _02054_ VGND VGND VPWR VPWR _02079_ sky130_fd_sc_hd__o211a_1
X_16513_ _03086_ _06509_ _08865_ VGND VGND VPWR VPWR _06908_ sky130_fd_sc_hd__and3b_1
X_13725_ _03861_ _03873_ VGND VGND VPWR VPWR _03874_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_85_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10937_ _00936_ _00935_ _00934_ VGND VGND VPWR VPWR _01030_ sky130_fd_sc_hd__a21o_1
XFILLER_0_86_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17493_ _07843_ _07847_ VGND VGND VPWR VPWR _07975_ sky130_fd_sc_hd__and2b_1
XFILLER_0_128_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16444_ _06775_ _06779_ _06832_ VGND VGND VPWR VPWR _06833_ sky130_fd_sc_hd__and3_1
X_13656_ _08713_ _09303_ _03795_ _03796_ VGND VGND VPWR VPWR _03798_ sky130_fd_sc_hd__nand4_2
XFILLER_0_38_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10868_ _00958_ _00960_ VGND VGND VPWR VPWR _00961_ sky130_fd_sc_hd__or2_1
XFILLER_0_26_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12607_ _02693_ _02696_ _02699_ VGND VGND VPWR VPWR _02700_ sky130_fd_sc_hd__nor3b_2
XPHY_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16375_ _06531_ _06533_ VGND VGND VPWR VPWR _06758_ sky130_fd_sc_hd__nor2_1
XFILLER_0_109_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13587_ _03674_ _03675_ _03720_ _03721_ VGND VGND VPWR VPWR _03723_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_53_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10799_ _00270_ _00271_ _00272_ _09348_ VGND VGND VPWR VPWR _00892_ sky130_fd_sc_hd__a22o_1
XPHY_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18114_ _08548_ _08562_ _08546_ VGND VGND VPWR VPWR _08651_ sky130_fd_sc_hd__a21o_1
X_15326_ _03165_ _05307_ _05621_ _03039_ VGND VGND VPWR VPWR _05622_ sky130_fd_sc_hd__o22a_1
X_12538_ _02628_ _02630_ VGND VGND VPWR VPWR _02631_ sky130_fd_sc_hd__and2_1
XFILLER_0_121_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_124_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18045_ _08482_ _08531_ _08575_ VGND VGND VPWR VPWR _08576_ sky130_fd_sc_hd__a21oi_1
X_15257_ _05537_ _05544_ VGND VGND VPWR VPWR _05546_ sky130_fd_sc_hd__nand2_1
X_12469_ _02561_ VGND VGND VPWR VPWR _02562_ sky130_fd_sc_hd__inv_2
XFILLER_0_124_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14208_ _03741_ _03902_ _04068_ _04236_ VGND VGND VPWR VPWR _04402_ sky130_fd_sc_hd__nor4_2
XFILLER_0_111_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15188_ _05465_ _05470_ VGND VGND VPWR VPWR _05471_ sky130_fd_sc_hd__xnor2_1
X_14139_ _04322_ _04324_ _04319_ VGND VGND VPWR VPWR _04326_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_10_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_120_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18947_ clknet_4_3_0_clk _09386_ VGND VGND VPWR VPWR salida\[0\] sky130_fd_sc_hd__dfxtp_2
X_09680_ _06019_ VGND VGND VPWR VPWR _06029_ sky130_fd_sc_hd__clkbuf_4
X_18878_ clknet_4_15_0_clk net248 VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__dfxtp_1
X_17829_ _06734_ _08243_ _08340_ _06461_ VGND VGND VPWR VPWR _08341_ sky130_fd_sc_hd__a211o_1
XFILLER_0_49_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09947_ _08692_ _08702_ _08919_ VGND VGND VPWR VPWR _08930_ sky130_fd_sc_hd__a21o_2
XTAP_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09878_ _07799_ _08169_ VGND VGND VPWR VPWR _08180_ sky130_fd_sc_hd__and2_2
XFILLER_0_99_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11840_ _01905_ _01907_ VGND VGND VPWR VPWR _01933_ sky130_fd_sc_hd__or2_1
XTAP_2624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_724 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11771_ _01106_ _01862_ _01863_ VGND VGND VPWR VPWR _01864_ sky130_fd_sc_hd__or3b_4
XTAP_1934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13510_ _03635_ _03636_ _03631_ _03419_ VGND VGND VPWR VPWR _03638_ sky130_fd_sc_hd__a211o_1
XTAP_1956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10722_ _08082_ _00814_ VGND VGND VPWR VPWR _00815_ sky130_fd_sc_hd__nor2_1
XTAP_1967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14490_ _02986_ _07156_ _04707_ _04708_ VGND VGND VPWR VPWR _04709_ sky130_fd_sc_hd__nand4_2
XTAP_1978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13441_ _03560_ _03561_ _03098_ VGND VGND VPWR VPWR _03562_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10653_ _00696_ _00697_ _00743_ _00744_ VGND VGND VPWR VPWR _00746_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_137_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_120 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_125_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16160_ _03003_ _03004_ _03018_ _06523_ VGND VGND VPWR VPWR _06524_ sky130_fd_sc_hd__or4_4
XFILLER_0_51_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13372_ _03484_ _03486_ VGND VGND VPWR VPWR _03488_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_63_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10584_ _00663_ _00664_ _00675_ VGND VGND VPWR VPWR _00677_ sky130_fd_sc_hd__and3_1
XFILLER_0_24_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15111_ _05260_ _05283_ _05386_ VGND VGND VPWR VPWR _05387_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_140_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12323_ _02414_ _02415_ VGND VGND VPWR VPWR _02416_ sky130_fd_sc_hd__or2_1
X_16091_ _03068_ _06448_ VGND VGND VPWR VPWR _06449_ sky130_fd_sc_hd__and2_1
XFILLER_0_133_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15042_ _05216_ _05217_ VGND VGND VPWR VPWR _05312_ sky130_fd_sc_hd__nand2_1
X_12254_ _02188_ VGND VGND VPWR VPWR _02347_ sky130_fd_sc_hd__buf_4
XFILLER_0_32_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11205_ _08713_ _08452_ _01002_ _01001_ VGND VGND VPWR VPWR _01298_ sky130_fd_sc_hd__a31o_1
XFILLER_0_76_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12185_ _02275_ _02276_ _02224_ VGND VGND VPWR VPWR _02278_ sky130_fd_sc_hd__a21oi_1
X_18801_ _09298_ _09309_ VGND VGND VPWR VPWR _09310_ sky130_fd_sc_hd__and2_1
X_11136_ _01187_ _01192_ _01196_ _01197_ VGND VGND VPWR VPWR _01229_ sky130_fd_sc_hd__a211oi_2
X_16993_ _07407_ _07427_ _07429_ VGND VGND VPWR VPWR _07430_ sky130_fd_sc_hd__and3_1
X_18732_ _09255_ VGND VGND VPWR VPWR _00069_ sky130_fd_sc_hd__clkbuf_1
X_11067_ _03345_ net242 _01031_ _07581_ VGND VGND VPWR VPWR _01160_ sky130_fd_sc_hd__and4_1
X_15944_ _02976_ _04241_ _03918_ _03036_ VGND VGND VPWR VPWR _06291_ sky130_fd_sc_hd__a31o_1
X_10018_ _00110_ VGND VGND VPWR VPWR _00111_ sky130_fd_sc_hd__inv_2
X_15875_ _06203_ _06215_ VGND VGND VPWR VPWR _06217_ sky130_fd_sc_hd__nor2_1
X_18663_ net65 _03094_ _09193_ VGND VGND VPWR VPWR _09206_ sky130_fd_sc_hd__mux2_1
X_17614_ _06750_ _07859_ VGND VGND VPWR VPWR _08107_ sky130_fd_sc_hd__nand2_1
XFILLER_0_59_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14826_ _05074_ _05076_ VGND VGND VPWR VPWR _05077_ sky130_fd_sc_hd__nand2_2
X_18594_ net289 _09140_ _09153_ _09144_ VGND VGND VPWR VPWR _00020_ sky130_fd_sc_hd__o211a_1
XFILLER_0_86_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_77 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14757_ _03006_ _02124_ VGND VGND VPWR VPWR _05001_ sky130_fd_sc_hd__nand2_1
X_17545_ _03693_ _06441_ _06426_ VGND VGND VPWR VPWR _08032_ sky130_fd_sc_hd__a21oi_1
X_11969_ _01913_ _01916_ VGND VGND VPWR VPWR _02062_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_129_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13708_ _00163_ _01866_ _03853_ VGND VGND VPWR VPWR _03855_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_46_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17476_ _06891_ _07390_ _07836_ _07834_ VGND VGND VPWR VPWR _07956_ sky130_fd_sc_hd__a31o_1
X_14688_ _04794_ _04796_ _04924_ _04925_ VGND VGND VPWR VPWR _04926_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_58_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_128_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13639_ _04690_ _07406_ _03776_ _03777_ VGND VGND VPWR VPWR _03779_ sky130_fd_sc_hd__o2bb2a_1
X_16427_ _06813_ VGND VGND VPWR VPWR _06814_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_128_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16358_ _06736_ _06738_ _03098_ VGND VGND VPWR VPWR _06739_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15309_ _05499_ _05602_ VGND VGND VPWR VPWR _05603_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_81_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_143_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16289_ _06660_ _06663_ _00494_ VGND VGND VPWR VPWR _06664_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_125_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18028_ _08455_ _08549_ _08555_ VGND VGND VPWR VPWR _08557_ sky130_fd_sc_hd__or3_1
XFILLER_0_100_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09801_ _05627_ _05725_ VGND VGND VPWR VPWR _07341_ sky130_fd_sc_hd__or2_1
X_09732_ ApproximateM_inst.lob_16.lob2.genblk1\[9\].genblk1.mux.sel VGND VGND VPWR
+ VPWR _06591_ sky130_fd_sc_hd__buf_4
X_09663_ _05322_ VGND VGND VPWR VPWR _05845_ sky130_fd_sc_hd__clkbuf_8
X_09594_ _05072_ _05083_ VGND VGND VPWR VPWR _05093_ sky130_fd_sc_hd__and2b_1
XTAP_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_687 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_143_692 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_131_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13990_ _04161_ _04162_ VGND VGND VPWR VPWR _04163_ sky130_fd_sc_hd__and2_1
XFILLER_0_99_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12941_ _02981_ _03033_ VGND VGND VPWR VPWR _03034_ sky130_fd_sc_hd__or2_1
XFILLER_0_87_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15660_ _05890_ _05983_ VGND VGND VPWR VPWR _05984_ sky130_fd_sc_hd__xnor2_1
X_12872_ op_code\[2\] op_code\[3\] VGND VGND VPWR VPWR _02965_ sky130_fd_sc_hd__nand2b_2
XTAP_2410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_100 _09374_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_111 net43 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14611_ _04835_ _04836_ _04839_ _04840_ VGND VGND VPWR VPWR _04841_ sky130_fd_sc_hd__o211ai_2
XANTENNA_122 _02646_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_133 _04191_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11823_ _01815_ _01915_ VGND VGND VPWR VPWR _01916_ sky130_fd_sc_hd__nor2_1
XFILLER_0_96_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15591_ _05811_ _05821_ _05819_ VGND VGND VPWR VPWR _05909_ sky130_fd_sc_hd__a21oi_1
XANTENNA_144 _08615_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_155 _08762_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_166 net172 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17330_ _02589_ _02844_ VGND VGND VPWR VPWR _07797_ sky130_fd_sc_hd__or2_1
XTAP_2487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14542_ _04764_ _04765_ VGND VGND VPWR VPWR _04767_ sky130_fd_sc_hd__xor2_1
XTAP_1753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_177 _02646_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11754_ _01082_ _01081_ ApproximateM_inst.lob_16.lob1.genblk1\[13\].genblk1.mux.sel
+ ApproximateM_inst.lob_16.lob1.genblk1\[12\].genblk1.mux.sel VGND VGND VPWR VPWR
+ _01847_ sky130_fd_sc_hd__and4_1
XTAP_1764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10705_ _04722_ _00780_ _00782_ VGND VGND VPWR VPWR _00798_ sky130_fd_sc_hd__a21o_1
XTAP_1797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17261_ _06880_ _07194_ _07290_ VGND VGND VPWR VPWR _07721_ sky130_fd_sc_hd__or3_2
X_14473_ _04551_ _04401_ net215 VGND VGND VPWR VPWR _04692_ sky130_fd_sc_hd__and3b_1
XFILLER_0_55_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11685_ _01776_ _01777_ VGND VGND VPWR VPWR _01778_ sky130_fd_sc_hd__nor2_1
X_16212_ _06579_ VGND VGND VPWR VPWR _06581_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_125_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19000_ clknet_4_4_0_clk _09367_ VGND VGND VPWR VPWR salida\[53\] sky130_fd_sc_hd__dfxtp_1
X_13424_ _03065_ _03075_ _02983_ VGND VGND VPWR VPWR _03545_ sky130_fd_sc_hd__mux2_1
X_10636_ _00106_ _00212_ VGND VGND VPWR VPWR _00729_ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17192_ _07643_ _07644_ VGND VGND VPWR VPWR _07647_ sky130_fd_sc_hd__nand2_1
XFILLER_0_51_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_478 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16143_ _02976_ _06505_ VGND VGND VPWR VPWR _06506_ sky130_fd_sc_hd__nand2_1
XFILLER_0_141_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13355_ net131 _03373_ _03467_ _03468_ VGND VGND VPWR VPWR _03469_ sky130_fd_sc_hd__o211ai_4
X_10567_ _00634_ _00635_ _00657_ _00658_ VGND VGND VPWR VPWR _00660_ sky130_fd_sc_hd__nand4_4
XFILLER_0_107_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12306_ _02392_ _02394_ _02393_ VGND VGND VPWR VPWR _02399_ sky130_fd_sc_hd__o21a_1
X_16074_ _01248_ _06430_ VGND VGND VPWR VPWR _06431_ sky130_fd_sc_hd__and2_1
X_13286_ _03390_ _03391_ _03392_ VGND VGND VPWR VPWR _03393_ sky130_fd_sc_hd__and3_2
X_10498_ _00164_ VGND VGND VPWR VPWR _00591_ sky130_fd_sc_hd__buf_4
X_15025_ _05059_ _05186_ _05293_ VGND VGND VPWR VPWR _05294_ sky130_fd_sc_hd__a21o_1
X_12237_ _02326_ _02329_ VGND VGND VPWR VPWR _02330_ sky130_fd_sc_hd__or2_1
X_12168_ _02258_ _02260_ VGND VGND VPWR VPWR _02261_ sky130_fd_sc_hd__and2_1
X_11119_ _05573_ _05595_ _04395_ _03739_ VGND VGND VPWR VPWR _01212_ sky130_fd_sc_hd__and4_1
X_12099_ _02191_ _02085_ VGND VGND VPWR VPWR _02192_ sky130_fd_sc_hd__xnor2_1
X_16976_ _06951_ _07035_ _07410_ net237 VGND VGND VPWR VPWR _07411_ sky130_fd_sc_hd__o22a_1
X_18715_ _09242_ VGND VGND VPWR VPWR _00064_ sky130_fd_sc_hd__clkbuf_1
Xinput6 i_wb_addr[13] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_1
X_15927_ _06270_ _06271_ VGND VGND VPWR VPWR _06272_ sky130_fd_sc_hd__nand2_1
X_18646_ net57 _09189_ _09192_ VGND VGND VPWR VPWR _00038_ sky130_fd_sc_hd__o21a_1
X_15858_ _06196_ _06197_ VGND VGND VPWR VPWR _06198_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_59_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14809_ _04920_ _04922_ VGND VGND VPWR VPWR _05058_ sky130_fd_sc_hd__nand2_1
XFILLER_0_143_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18577_ _09113_ VGND VGND VPWR VPWR _09141_ sky130_fd_sc_hd__clkbuf_4
X_15789_ _06097_ _06123_ VGND VGND VPWR VPWR _06124_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17528_ _08011_ _08012_ VGND VGND VPWR VPWR _08013_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_86_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17459_ _06657_ _07708_ VGND VGND VPWR VPWR _07937_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_602 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_117_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_104_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09715_ _04340_ _04362_ _05028_ cla_inst.in1\[16\] VGND VGND VPWR VPWR _06406_ sky130_fd_sc_hd__and4_1
X_09646_ _05649_ _05606_ _05617_ _05573_ VGND VGND VPWR VPWR _05660_ sky130_fd_sc_hd__a22o_1
XTAP_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09577_ _04875_ _04897_ VGND VGND VPWR VPWR _04908_ sky130_fd_sc_hd__nor2_1
XTAP_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_811 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_154_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_147_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_579 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11470_ _01550_ _01561_ VGND VGND VPWR VPWR _01563_ sky130_fd_sc_hd__and2_1
XFILLER_0_92_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10421_ ApproximateM_inst.lob_16.lob2.mux.sel VGND VGND VPWR VPWR _00514_ sky130_fd_sc_hd__clkinv_4
XFILLER_0_61_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_448 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13140_ _03224_ _03225_ _03236_ VGND VGND VPWR VPWR _03237_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_61_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10352_ _00442_ _00444_ VGND VGND VPWR VPWR _00445_ sky130_fd_sc_hd__xor2_1
XFILLER_0_20_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13071_ _03161_ _03162_ VGND VGND VPWR VPWR _03163_ sky130_fd_sc_hd__nand2_1
X_10283_ _00333_ _00335_ _08681_ _09005_ VGND VGND VPWR VPWR _00376_ sky130_fd_sc_hd__o211a_1
X_12022_ _02112_ _02114_ VGND VGND VPWR VPWR _02115_ sky130_fd_sc_hd__nor2_1
X_16830_ _07158_ _07159_ _07251_ VGND VGND VPWR VPWR _07252_ sky130_fd_sc_hd__a21oi_2
X_13973_ _04123_ _04124_ _04142_ VGND VGND VPWR VPWR _04145_ sky130_fd_sc_hd__nor3_4
XFILLER_0_73_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16761_ _06355_ _06790_ _07176_ _03094_ VGND VGND VPWR VPWR _07177_ sky130_fd_sc_hd__a22o_1
X_18500_ _03916_ _06999_ _08141_ _09066_ _09067_ VGND VGND VPWR VPWR _09068_ sky130_fd_sc_hd__o311a_1
X_15712_ _01359_ _04125_ _06038_ _06039_ VGND VGND VPWR VPWR _06041_ sky130_fd_sc_hd__and4_1
X_12924_ _03007_ _03011_ _03013_ _03016_ VGND VGND VPWR VPWR _03017_ sky130_fd_sc_hd__or4_2
X_16692_ _07072_ _07075_ _07101_ _06723_ _02214_ VGND VGND VPWR VPWR _09415_ sky130_fd_sc_hd__o32a_2
XFILLER_0_69_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18431_ _03119_ _06266_ _07579_ _08141_ _08993_ VGND VGND VPWR VPWR _08994_ sky130_fd_sc_hd__o221a_1
X_15643_ _05958_ _05965_ VGND VGND VPWR VPWR _05966_ sky130_fd_sc_hd__or2_1
X_12855_ _02942_ _02947_ VGND VGND VPWR VPWR _02948_ sky130_fd_sc_hd__xnor2_1
XTAP_2240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11806_ _01876_ _01897_ _01898_ VGND VGND VPWR VPWR _01899_ sky130_fd_sc_hd__and3_1
X_15574_ _05882_ _05889_ VGND VGND VPWR VPWR _05891_ sky130_fd_sc_hd__nand2_1
XTAP_2284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18362_ _08868_ _08918_ VGND VGND VPWR VPWR _08920_ sky130_fd_sc_hd__nor2_1
XTAP_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12786_ _02863_ _02872_ _02878_ VGND VGND VPWR VPWR _02879_ sky130_fd_sc_hd__and3_1
XTAP_2295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14525_ _07537_ _01962_ VGND VGND VPWR VPWR _04748_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17313_ _07776_ _07778_ VGND VGND VPWR VPWR _07779_ sky130_fd_sc_hd__and2b_1
XTAP_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11737_ _06591_ _03607_ _00774_ _00806_ VGND VGND VPWR VPWR _01830_ sky130_fd_sc_hd__a22o_1
XFILLER_0_44_708 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18293_ _04668_ _04679_ _07743_ VGND VGND VPWR VPWR _08845_ sky130_fd_sc_hd__nor3_1
X_14456_ _04670_ _04671_ _04484_ VGND VGND VPWR VPWR _04673_ sky130_fd_sc_hd__o21ai_1
X_17244_ _07589_ _07601_ VGND VGND VPWR VPWR _07703_ sky130_fd_sc_hd__nor2_1
XFILLER_0_4_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11668_ _01201_ _01759_ _01757_ _01758_ VGND VGND VPWR VPWR _01761_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_142_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13407_ _03523_ _03524_ _03367_ _03369_ VGND VGND VPWR VPWR _03526_ sky130_fd_sc_hd__o211a_1
XFILLER_0_98_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10619_ _00700_ _00701_ _00711_ VGND VGND VPWR VPWR _00712_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_107_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17175_ _07622_ _07625_ _07626_ VGND VGND VPWR VPWR _07628_ sky130_fd_sc_hd__a21oi_1
X_14387_ _04584_ _04585_ _04595_ VGND VGND VPWR VPWR _04597_ sky130_fd_sc_hd__or3_4
XFILLER_0_4_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11599_ _05246_ VGND VGND VPWR VPWR _01692_ sky130_fd_sc_hd__inv_6
XFILLER_0_3_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16126_ _02728_ _03002_ _03021_ VGND VGND VPWR VPWR _06487_ sky130_fd_sc_hd__or3_2
X_13338_ _03280_ _03284_ VGND VGND VPWR VPWR _03450_ sky130_fd_sc_hd__nand2_1
X_16057_ _06024_ _06410_ _06411_ _06328_ VGND VGND VPWR VPWR _06412_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_11_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13269_ _00620_ net136 _03237_ _03238_ VGND VGND VPWR VPWR _03374_ sky130_fd_sc_hd__o211a_2
XFILLER_0_121_172 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15008_ _05273_ _05274_ VGND VGND VPWR VPWR _05275_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_37_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16959_ _07388_ _07391_ VGND VGND VPWR VPWR _07392_ sky130_fd_sc_hd__nand2_1
X_09500_ _04056_ VGND VGND VPWR VPWR _04067_ sky130_fd_sc_hd__buf_6
XFILLER_0_79_638 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09431_ sel_op\[0\] VGND VGND VPWR VPWR _03313_ sky130_fd_sc_hd__clkbuf_4
X_18629_ salida\[31\] _09113_ _09117_ salida\[63\] _09127_ VGND VGND VPWR VPWR _09177_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_149_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_11 _00644_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_22 _01115_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_33 _01266_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_44 _02533_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_55 _03760_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_66 _04649_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_77 _07123_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_88 _08820_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_99 _08934_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_868 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10970_ _05671_ _05039_ VGND VGND VPWR VPWR _01063_ sky130_fd_sc_hd__nand2_1
X_09629_ _05453_ _05464_ _05388_ _05050_ VGND VGND VPWR VPWR _05475_ sky130_fd_sc_hd__nand4_2
X_12640_ _02700_ _02731_ _02732_ VGND VGND VPWR VPWR _02733_ sky130_fd_sc_hd__or3_4
XFILLER_0_65_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12571_ _02622_ _02659_ _02662_ VGND VGND VPWR VPWR _02664_ sky130_fd_sc_hd__or3b_1
XFILLER_0_108_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14310_ _04359_ _04367_ VGND VGND VPWR VPWR _04513_ sky130_fd_sc_hd__and2_1
XFILLER_0_135_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11522_ _01613_ _01614_ VGND VGND VPWR VPWR _01615_ sky130_fd_sc_hd__and2b_1
X_15290_ _05481_ _05484_ _05482_ VGND VGND VPWR VPWR _05582_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_124_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14241_ _03859_ _04132_ _07015_ _07112_ VGND VGND VPWR VPWR _04437_ sky130_fd_sc_hd__and4_1
X_11453_ _01543_ _01544_ _01545_ VGND VGND VPWR VPWR _01546_ sky130_fd_sc_hd__and3_1
XFILLER_0_135_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10404_ _05736_ _07025_ _00317_ _00319_ _00318_ VGND VGND VPWR VPWR _00497_ sky130_fd_sc_hd__a32o_1
X_14172_ _00148_ _00149_ _08409_ _03750_ VGND VGND VPWR VPWR _04363_ sky130_fd_sc_hd__and4_1
X_11384_ _00204_ _00878_ VGND VGND VPWR VPWR _01477_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13123_ _04001_ _05257_ VGND VGND VPWR VPWR _03219_ sky130_fd_sc_hd__nand2_1
X_10335_ _00268_ VGND VGND VPWR VPWR _00428_ sky130_fd_sc_hd__inv_2
X_18980_ clknet_4_0_0_clk _09355_ VGND VGND VPWR VPWR salida\[33\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_103_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13054_ _03145_ VGND VGND VPWR VPWR _03146_ sky130_fd_sc_hd__inv_2
X_17931_ _08358_ _08359_ _08360_ _08356_ VGND VGND VPWR VPWR _08451_ sky130_fd_sc_hd__nor4b_1
X_10266_ _00358_ _07504_ _00127_ VGND VGND VPWR VPWR _00359_ sky130_fd_sc_hd__and3_1
X_12005_ _02092_ _02097_ VGND VGND VPWR VPWR _02098_ sky130_fd_sc_hd__xnor2_1
X_17862_ _08367_ _08375_ VGND VGND VPWR VPWR _08377_ sky130_fd_sc_hd__xnor2_1
X_10197_ _08474_ _08485_ _08398_ VGND VGND VPWR VPWR _00290_ sky130_fd_sc_hd__a21bo_1
X_16813_ _07127_ _07131_ _07128_ VGND VGND VPWR VPWR _07234_ sky130_fd_sc_hd__o21ai_2
X_17793_ _08299_ _08301_ VGND VGND VPWR VPWR _08302_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16744_ _07067_ _07070_ _07066_ VGND VGND VPWR VPWR _07159_ sky130_fd_sc_hd__a21o_1
X_13956_ _03790_ _04125_ _03976_ VGND VGND VPWR VPWR _04126_ sky130_fd_sc_hd__and3_1
XFILLER_0_88_424 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12907_ _02999_ VGND VGND VPWR VPWR _03000_ sky130_fd_sc_hd__clkbuf_4
X_13887_ _04004_ _04005_ _04048_ _04049_ VGND VGND VPWR VPWR _04051_ sky130_fd_sc_hd__o22ai_2
X_16675_ _06598_ VGND VGND VPWR VPWR _07084_ sky130_fd_sc_hd__buf_4
XFILLER_0_69_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18414_ _08749_ _08810_ _08972_ _08975_ VGND VGND VPWR VPWR _08976_ sky130_fd_sc_hd__o31a_1
X_12838_ _02909_ _02911_ VGND VGND VPWR VPWR _02931_ sky130_fd_sc_hd__or2b_2
X_15626_ _05786_ _05788_ VGND VGND VPWR VPWR _05948_ sky130_fd_sc_hd__xnor2_1
XTAP_2070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18345_ _04537_ _07743_ _08900_ VGND VGND VPWR VPWR _08901_ sky130_fd_sc_hd__or3_1
X_15557_ _05870_ _05871_ _05872_ VGND VGND VPWR VPWR _05873_ sky130_fd_sc_hd__nor3_1
XTAP_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_663 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12769_ _01802_ _01804_ VGND VGND VPWR VPWR _02862_ sky130_fd_sc_hd__nand2_1
XTAP_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_123_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14508_ _04727_ _04728_ VGND VGND VPWR VPWR _04729_ sky130_fd_sc_hd__xor2_2
XFILLER_0_44_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15488_ _05789_ _05796_ VGND VGND VPWR VPWR _05798_ sky130_fd_sc_hd__nand2_1
X_18276_ _06401_ _06546_ _08826_ _03056_ VGND VGND VPWR VPWR _08827_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_127_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_126_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_142_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_154_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_56 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput20 i_wb_addr[26] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__clkbuf_1
X_17227_ _06508_ _07683_ _07684_ VGND VGND VPWR VPWR _07685_ sky130_fd_sc_hd__and3_1
Xinput31 i_wb_addr[7] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__clkbuf_1
X_14439_ _04475_ _04477_ VGND VGND VPWR VPWR _04654_ sky130_fd_sc_hd__nor2_1
XFILLER_0_141_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput42 i_wb_data[16] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_142_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput53 i_wb_data[26] VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__buf_1
Xinput64 i_wb_data[7] VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__buf_2
XFILLER_0_24_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17158_ _07018_ _07195_ _07608_ _06766_ VGND VGND VPWR VPWR _07609_ sky130_fd_sc_hd__o22a_1
XFILLER_0_12_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16109_ _03089_ _02125_ _03179_ VGND VGND VPWR VPWR _06468_ sky130_fd_sc_hd__or3_1
X_09980_ _07537_ _09219_ _09197_ _09205_ VGND VGND VPWR VPWR _09232_ sky130_fd_sc_hd__o2bb2a_1
X_17089_ _07531_ _07532_ _07507_ VGND VGND VPWR VPWR _07534_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_654 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_595 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_643 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10120_ _00212_ VGND VGND VPWR VPWR _00213_ sky130_fd_sc_hd__buf_4
X_10051_ _00126_ _00133_ VGND VGND VPWR VPWR _00144_ sky130_fd_sc_hd__or2_1
XFILLER_0_100_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13810_ _03775_ _03780_ VGND VGND VPWR VPWR _03966_ sky130_fd_sc_hd__and2_1
X_14790_ _02999_ _01112_ _04893_ VGND VGND VPWR VPWR _05037_ sky130_fd_sc_hd__nand3_1
XFILLER_0_98_744 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13741_ _03718_ _03890_ VGND VGND VPWR VPWR _03891_ sky130_fd_sc_hd__nor2_1
X_10953_ _04493_ _04416_ _00949_ _03421_ VGND VGND VPWR VPWR _01046_ sky130_fd_sc_hd__and4_1
XFILLER_0_39_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_799 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13672_ _03625_ _03628_ _03626_ VGND VGND VPWR VPWR _03816_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_97_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16460_ _02974_ _06847_ _06849_ _06645_ VGND VGND VPWR VPWR _06850_ sky130_fd_sc_hd__a211o_1
X_10884_ _00966_ _00918_ net191 VGND VGND VPWR VPWR _00977_ sky130_fd_sc_hd__nor3_1
X_15411_ _05711_ _05712_ _05713_ VGND VGND VPWR VPWR _05714_ sky130_fd_sc_hd__o21a_1
X_12623_ _02713_ _02715_ VGND VGND VPWR VPWR _02716_ sky130_fd_sc_hd__nand2_1
X_16391_ _06669_ _06774_ VGND VGND VPWR VPWR _06775_ sky130_fd_sc_hd__or2b_1
XFILLER_0_39_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15342_ _05632_ _05636_ _05637_ VGND VGND VPWR VPWR _05639_ sky130_fd_sc_hd__and3_1
X_18130_ _08582_ _08667_ VGND VGND VPWR VPWR _08668_ sky130_fd_sc_hd__xnor2_1
X_12554_ ApproximateM_inst.lob_16.lob2.genblk1\[1\].genblk1.mux.sel _00177_ _02646_
+ VGND VGND VPWR VPWR _02647_ sky130_fd_sc_hd__nand3_1
XFILLER_0_65_195 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11505_ _04045_ _01596_ _01597_ VGND VGND VPWR VPWR _01598_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_136_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15273_ _05446_ _05448_ _05561_ VGND VGND VPWR VPWR _05564_ sky130_fd_sc_hd__nor3_1
X_18061_ _02175_ _08423_ _02170_ VGND VGND VPWR VPWR _08593_ sky130_fd_sc_hd__o21a_1
XFILLER_0_108_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12485_ _02576_ _02577_ VGND VGND VPWR VPWR _02578_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_124_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17012_ _07345_ _07349_ _07449_ VGND VGND VPWR VPWR _07451_ sky130_fd_sc_hd__o21a_1
X_14224_ _03539_ _04241_ _04415_ _04418_ VGND VGND VPWR VPWR _04419_ sky130_fd_sc_hd__a31o_1
X_11436_ _04548_ _03618_ _01527_ _01528_ VGND VGND VPWR VPWR _01529_ sky130_fd_sc_hd__nand4_2
XFILLER_0_21_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14155_ _04342_ _04343_ VGND VGND VPWR VPWR _04344_ sky130_fd_sc_hd__xnor2_1
X_11367_ _01455_ _01456_ _01458_ _01459_ VGND VGND VPWR VPWR _01460_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13106_ _02965_ _02966_ VGND VGND VPWR VPWR _03200_ sky130_fd_sc_hd__nor2_1
XTAP_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10318_ _00403_ _00410_ VGND VGND VPWR VPWR _00411_ sky130_fd_sc_hd__xnor2_1
X_14086_ _04100_ _04105_ VGND VGND VPWR VPWR _04268_ sky130_fd_sc_hd__nor2_1
X_18963_ clknet_4_6_0_clk _09393_ VGND VGND VPWR VPWR salida\[16\] sky130_fd_sc_hd__dfxtp_1
XTAP_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11298_ _00794_ _01381_ _01279_ _01380_ VGND VGND VPWR VPWR _01391_ sky130_fd_sc_hd__a211o_1
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17914_ _06847_ _08036_ _03197_ _05800_ VGND VGND VPWR VPWR _08434_ sky130_fd_sc_hd__a2bb2o_1
X_13037_ _03023_ _03128_ VGND VGND VPWR VPWR _03129_ sky130_fd_sc_hd__nand2_1
X_10249_ _07363_ _09248_ VGND VGND VPWR VPWR _00342_ sky130_fd_sc_hd__nand2_1
X_18894_ clknet_4_11_0_clk _00048_ VGND VGND VPWR VPWR ApproximateM_inst.lob_16.lob1.genblk1\[12\].genblk1.mux.sel
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_0_119_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17845_ _08262_ _08357_ VGND VGND VPWR VPWR _08358_ sky130_fd_sc_hd__nor2_1
XFILLER_0_88_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17776_ _08281_ _08282_ VGND VGND VPWR VPWR _08283_ sky130_fd_sc_hd__nand2_1
X_14988_ _05251_ _05252_ VGND VGND VPWR VPWR _05253_ sky130_fd_sc_hd__or2_1
XFILLER_0_88_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16727_ _07021_ _07045_ VGND VGND VPWR VPWR _07140_ sky130_fd_sc_hd__nor2_1
X_13939_ _04092_ _03945_ _04106_ VGND VGND VPWR VPWR _04107_ sky130_fd_sc_hd__o21a_2
XFILLER_0_76_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16658_ _06936_ _06979_ _07064_ VGND VGND VPWR VPWR _07065_ sky130_fd_sc_hd__a21o_1
XFILLER_0_69_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15609_ _05828_ _05893_ _05927_ _05928_ VGND VGND VPWR VPWR _05929_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_151_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16589_ _02728_ _06988_ _06989_ VGND VGND VPWR VPWR _06990_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_60_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18328_ _01417_ _06593_ _06594_ VGND VGND VPWR VPWR _08883_ sky130_fd_sc_hd__a21o_1
XFILLER_0_127_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18259_ _08804_ _08806_ VGND VGND VPWR VPWR _08808_ sky130_fd_sc_hd__or2_1
XFILLER_0_114_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_733 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_114_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09963_ _07232_ _07080_ _07374_ _07406_ VGND VGND VPWR VPWR _09101_ sky130_fd_sc_hd__and4_1
X_09894_ _03377_ _04886_ _03837_ _03356_ VGND VGND VPWR VPWR _08354_ sky130_fd_sc_hd__a22o_1
XTAP_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_758 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_137_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_8_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_8_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_63_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_145_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12270_ _02242_ _02241_ VGND VGND VPWR VPWR _02363_ sky130_fd_sc_hd__and2b_1
XFILLER_0_121_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11221_ _01104_ _01116_ VGND VGND VPWR VPWR _01314_ sky130_fd_sc_hd__or2_1
XFILLER_0_120_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11152_ cla_inst.in2\[21\] _00108_ _01241_ _01244_ VGND VGND VPWR VPWR _01245_ sky130_fd_sc_hd__o2bb2a_1
X_10103_ ApproximateM_inst.lob_16.lob1.genblk1\[3\].genblk1.mux.sel VGND VGND VPWR
+ VPWR _00196_ sky130_fd_sc_hd__buf_6
XFILLER_0_101_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11083_ _01171_ _01175_ VGND VGND VPWR VPWR _01176_ sky130_fd_sc_hd__xor2_2
X_15960_ _06304_ _06305_ VGND VGND VPWR VPWR _06307_ sky130_fd_sc_hd__nand2_1
X_14911_ _05167_ _05168_ VGND VGND VPWR VPWR _05169_ sky130_fd_sc_hd__xnor2_1
X_10034_ _09212_ VGND VGND VPWR VPWR _00127_ sky130_fd_sc_hd__clkbuf_8
X_15891_ _06221_ _06222_ VGND VGND VPWR VPWR _06233_ sky130_fd_sc_hd__nand2_1
X_17630_ _06559_ _08123_ VGND VGND VPWR VPWR _08124_ sky130_fd_sc_hd__or2_1
X_14842_ _03912_ _04075_ VGND VGND VPWR VPWR _05094_ sky130_fd_sc_hd__nand2_1
X_17561_ _06653_ _06756_ _08047_ VGND VGND VPWR VPWR _08048_ sky130_fd_sc_hd__nor3_1
X_14773_ _03014_ _05921_ _04871_ _04870_ VGND VGND VPWR VPWR _05019_ sky130_fd_sc_hd__a31o_1
X_11985_ _01984_ _02054_ _02073_ _02077_ VGND VGND VPWR VPWR _02078_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_85_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16512_ _02828_ _02968_ _06905_ VGND VGND VPWR VPWR _06907_ sky130_fd_sc_hd__or3_1
X_13724_ _03862_ _03872_ VGND VGND VPWR VPWR _03873_ sky130_fd_sc_hd__xor2_1
X_10936_ _00936_ _00934_ _00935_ VGND VGND VPWR VPWR _01029_ sky130_fd_sc_hd__nand3_1
X_17492_ _07971_ _07972_ VGND VGND VPWR VPWR _07974_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16443_ _06828_ _06831_ VGND VGND VPWR VPWR _06832_ sky130_fd_sc_hd__xor2_1
X_13655_ _08724_ _09248_ _03795_ _03796_ VGND VGND VPWR VPWR _03797_ sky130_fd_sc_hd__a22o_1
X_10867_ _03717_ _03410_ _00956_ _00959_ VGND VGND VPWR VPWR _00960_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_85_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12606_ _02697_ _02698_ VGND VGND VPWR VPWR _02699_ sky130_fd_sc_hd__xnor2_1
X_13586_ _03674_ _03675_ _03720_ _03721_ VGND VGND VPWR VPWR _03722_ sky130_fd_sc_hd__and4_1
X_16374_ _06563_ _06756_ VGND VGND VPWR VPWR _06757_ sky130_fd_sc_hd__nor2_1
XPHY_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10798_ _00856_ _00889_ _00890_ VGND VGND VPWR VPWR _00891_ sky130_fd_sc_hd__nor3_2
XPHY_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18113_ _08634_ _08649_ VGND VGND VPWR VPWR _08650_ sky130_fd_sc_hd__xor2_1
X_15325_ _03132_ _03193_ _03536_ VGND VGND VPWR VPWR _05621_ sky130_fd_sc_hd__mux2_1
X_12537_ _02616_ _02629_ VGND VGND VPWR VPWR _02630_ sky130_fd_sc_hd__or2b_1
XFILLER_0_121_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18044_ _08573_ _08574_ VGND VGND VPWR VPWR _08575_ sky130_fd_sc_hd__nand2_1
X_15256_ _05537_ _05544_ VGND VGND VPWR VPWR _05545_ sky130_fd_sc_hd__or2_1
X_12468_ _02502_ _02559_ VGND VGND VPWR VPWR _02561_ sky130_fd_sc_hd__nand2_1
X_14207_ _04399_ _04400_ VGND VGND VPWR VPWR _04401_ sky130_fd_sc_hd__xor2_2
X_11419_ _04984_ _00131_ VGND VGND VPWR VPWR _01512_ sky130_fd_sc_hd__nand2_1
X_15187_ _05468_ _05469_ VGND VGND VPWR VPWR _05470_ sky130_fd_sc_hd__or2_1
X_12399_ ApproximateM_inst.lob_16.lob2.genblk1\[2\].genblk1.mux.sel _00774_ VGND VGND
+ VPWR VPWR _02492_ sky130_fd_sc_hd__and2_1
X_14138_ _04319_ _04322_ _04324_ VGND VGND VPWR VPWR _04325_ sky130_fd_sc_hd__or3_1
XFILLER_0_10_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_120_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18946_ clknet_4_2_0_clk _00100_ VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__dfxtp_2
X_14069_ _02975_ _03547_ _04249_ VGND VGND VPWR VPWR _04250_ sky130_fd_sc_hd__or3_1
XFILLER_0_55_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18877_ clknet_4_15_0_clk net313 VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__dfxtp_1
X_17828_ _06387_ _06545_ _08339_ _03041_ VGND VGND VPWR VPWR _08340_ sky130_fd_sc_hd__a22o_1
X_17759_ _08153_ _08154_ _08152_ VGND VGND VPWR VPWR _08264_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_76_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_30 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_279 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_119_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_cap150 _06804_ VGND VGND VPWR VPWR net150 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_13_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09946_ _08822_ _08908_ VGND VGND VPWR VPWR _08919_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_110_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09877_ cla_inst.in1\[27\] VGND VGND VPWR VPWR _08169_ sky130_fd_sc_hd__buf_4
XTAP_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11770_ _00120_ _06471_ VGND VGND VPWR VPWR _01863_ sky130_fd_sc_hd__and2_4
XTAP_1924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10721_ _00812_ _08071_ _06765_ _00813_ VGND VGND VPWR VPWR _00814_ sky130_fd_sc_hd__o2bb2a_1
XTAP_1957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13440_ _03129_ _03168_ _03048_ VGND VGND VPWR VPWR _03561_ sky130_fd_sc_hd__mux2_1
X_10652_ _00696_ _00697_ _00743_ _00744_ VGND VGND VPWR VPWR _00745_ sky130_fd_sc_hd__or4_4
XFILLER_0_137_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13371_ _03485_ _03305_ VGND VGND VPWR VPWR _03486_ sky130_fd_sc_hd__nand2_1
XFILLER_0_91_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10583_ _00663_ _00664_ _00675_ VGND VGND VPWR VPWR _00676_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_63_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15110_ _05384_ _05385_ VGND VGND VPWR VPWR _05386_ sky130_fd_sc_hd__nand2_1
X_12322_ _02346_ _02349_ VGND VGND VPWR VPWR _02415_ sky130_fd_sc_hd__xor2_1
X_16090_ _03143_ _03056_ _06447_ VGND VGND VPWR VPWR _06448_ sky130_fd_sc_hd__and3_1
XFILLER_0_106_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15041_ _05285_ _05286_ VGND VGND VPWR VPWR _05310_ sky130_fd_sc_hd__nor2_1
XFILLER_0_32_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12253_ _02344_ _02345_ VGND VGND VPWR VPWR _02346_ sky130_fd_sc_hd__or2_1
X_11204_ _01295_ _01296_ VGND VGND VPWR VPWR _01297_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_31_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12184_ _02275_ _02224_ _02276_ VGND VGND VPWR VPWR _02277_ sky130_fd_sc_hd__and3_1
X_18800_ _02997_ net50 _09301_ VGND VGND VPWR VPWR _09309_ sky130_fd_sc_hd__mux2_1
X_11135_ _01217_ _01219_ _01227_ VGND VGND VPWR VPWR _01228_ sky130_fd_sc_hd__or3_1
XFILLER_0_101_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16992_ _07408_ _07323_ _07425_ VGND VGND VPWR VPWR _07429_ sky130_fd_sc_hd__nand3_1
X_18731_ _09245_ _09254_ VGND VGND VPWR VPWR _09255_ sky130_fd_sc_hd__and2_1
X_11066_ _03454_ _07548_ VGND VGND VPWR VPWR _01159_ sky130_fd_sc_hd__and2_1
X_15943_ _06265_ _06269_ _06287_ VGND VGND VPWR VPWR _06290_ sky130_fd_sc_hd__o21ai_1
X_10017_ _00109_ _09349_ _09188_ _07591_ VGND VGND VPWR VPWR _00110_ sky130_fd_sc_hd__and4_1
X_18662_ _09204_ VGND VGND VPWR VPWR _00043_ sky130_fd_sc_hd__clkbuf_1
X_15874_ _06203_ _06215_ VGND VGND VPWR VPWR _06216_ sky130_fd_sc_hd__and2_1
XFILLER_0_99_850 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17613_ _07978_ _08105_ VGND VGND VPWR VPWR _08106_ sky130_fd_sc_hd__xnor2_1
X_14825_ _05075_ VGND VGND VPWR VPWR _05076_ sky130_fd_sc_hd__inv_2
X_18593_ salida\[16\] _09141_ _09142_ salida\[48\] _09146_ VGND VGND VPWR VPWR _09153_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_99_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17544_ _06379_ _06378_ _06377_ VGND VGND VPWR VPWR _08031_ sky130_fd_sc_hd__a21o_1
X_14756_ _04997_ _04998_ _04862_ _04969_ VGND VGND VPWR VPWR _05000_ sky130_fd_sc_hd__a211o_1
XFILLER_0_25_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11968_ _01905_ _02058_ _02060_ VGND VGND VPWR VPWR _02061_ sky130_fd_sc_hd__and3_1
XFILLER_0_47_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13707_ _00163_ _01866_ _03853_ VGND VGND VPWR VPWR _03854_ sky130_fd_sc_hd__and3_1
X_10919_ _01008_ _01011_ VGND VGND VPWR VPWR _01012_ sky130_fd_sc_hd__xor2_1
XFILLER_0_58_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17475_ _07143_ _07721_ _07844_ _07846_ VGND VGND VPWR VPWR _07955_ sky130_fd_sc_hd__o22ai_2
X_14687_ _04922_ _04923_ _04884_ VGND VGND VPWR VPWR _04925_ sky130_fd_sc_hd__a21o_1
X_11899_ _01899_ _01904_ _01991_ VGND VGND VPWR VPWR _01992_ sky130_fd_sc_hd__or3_4
X_16426_ _06812_ net150 VGND VGND VPWR VPWR _06813_ sky130_fd_sc_hd__and2_1
X_13638_ _03776_ _03777_ _04548_ _07406_ VGND VGND VPWR VPWR _03778_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_41_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_690 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16357_ _03089_ _02272_ _03104_ _06626_ _06737_ VGND VGND VPWR VPWR _06738_ sky130_fd_sc_hd__o311a_1
X_13569_ _09350_ _04154_ _00165_ _00112_ VGND VGND VPWR VPWR _03703_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_125_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15308_ _05600_ _05601_ VGND VGND VPWR VPWR _05602_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_41_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16288_ _06661_ _06662_ _03324_ VGND VGND VPWR VPWR _06663_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_140_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18027_ _08455_ _08549_ _08555_ VGND VGND VPWR VPWR _08556_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_151_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15239_ _05441_ _05432_ VGND VGND VPWR VPWR _05526_ sky130_fd_sc_hd__and2b_1
XFILLER_0_1_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09800_ _07145_ _07178_ VGND VGND VPWR VPWR _07330_ sky130_fd_sc_hd__nand2_1
X_09731_ _05224_ _06062_ VGND VGND VPWR VPWR _06580_ sky130_fd_sc_hd__nand2_1
X_18929_ clknet_4_12_0_clk _00083_ VGND VGND VPWR VPWR ApproximateM_inst.lob_16.lob2.genblk2.mux_final.sel
+ sky130_fd_sc_hd__dfxtp_1
X_09662_ _05235_ VGND VGND VPWR VPWR _05834_ sky130_fd_sc_hd__buf_4
X_09593_ _04427_ _04569_ _04384_ _04635_ VGND VGND VPWR VPWR _05083_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_147_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_830 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_143_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09929_ _08724_ _05975_ VGND VGND VPWR VPWR _08735_ sky130_fd_sc_hd__nand2_1
X_12940_ _02983_ _03032_ VGND VGND VPWR VPWR _03033_ sky130_fd_sc_hd__or2_1
XTAP_2400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12871_ _00908_ _02963_ _00906_ VGND VGND VPWR VPWR _02964_ sky130_fd_sc_hd__a21o_1
XTAP_2411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_101 _09395_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_112 net43 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14610_ _01521_ _07015_ _04837_ _04838_ VGND VGND VPWR VPWR _04840_ sky130_fd_sc_hd__a22o_1
XANTENNA_123 _02783_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_134 _05279_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11822_ _04001_ _09219_ _01813_ _01914_ VGND VGND VPWR VPWR _01915_ sky130_fd_sc_hd__o2bb2a_1
XTAP_2444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15590_ _05855_ _05907_ VGND VGND VPWR VPWR _05908_ sky130_fd_sc_hd__xnor2_1
XTAP_1710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_145 _08674_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_156 _08762_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_167 _02646_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14541_ _01504_ _00461_ _04634_ _04633_ VGND VGND VPWR VPWR _04765_ sky130_fd_sc_hd__a31o_1
X_11753_ _01081_ ApproximateM_inst.lob_16.lob1.genblk1\[13\].genblk1.mux.sel ApproximateM_inst.lob_16.lob1.genblk1\[12\].genblk1.mux.sel
+ _01082_ VGND VGND VPWR VPWR _01846_ sky130_fd_sc_hd__a22o_1
XFILLER_0_83_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_178 _02646_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10704_ _00779_ _00794_ _00795_ _00796_ VGND VGND VPWR VPWR _00797_ sky130_fd_sc_hd__a211oi_4
XTAP_1787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17260_ _06657_ net145 _07598_ _07597_ VGND VGND VPWR VPWR _07720_ sky130_fd_sc_hd__a31o_1
X_14472_ _04688_ _04689_ VGND VGND VPWR VPWR _04691_ sky130_fd_sc_hd__xnor2_2
X_11684_ _01733_ _01772_ _01775_ VGND VGND VPWR VPWR _01777_ sky130_fd_sc_hd__nor3_1
XTAP_1798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16211_ _06578_ VGND VGND VPWR VPWR _06579_ sky130_fd_sc_hd__buf_2
X_10635_ _00726_ _00727_ VGND VGND VPWR VPWR _00728_ sky130_fd_sc_hd__nor2_1
XFILLER_0_102_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13423_ _03543_ VGND VGND VPWR VPWR _03544_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_125_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17191_ _07643_ _07644_ VGND VGND VPWR VPWR _07645_ sky130_fd_sc_hd__nor2_1
XFILLER_0_36_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13354_ _03434_ _03435_ _03466_ VGND VGND VPWR VPWR _03468_ sky130_fd_sc_hd__o21ai_2
X_16142_ _06494_ _06503_ _03080_ VGND VGND VPWR VPWR _06505_ sky130_fd_sc_hd__mux2_1
X_10566_ _00634_ _00635_ _00657_ _00658_ VGND VGND VPWR VPWR _00659_ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12305_ _02397_ VGND VGND VPWR VPWR _02398_ sky130_fd_sc_hd__inv_2
X_13285_ _03214_ _03220_ _03213_ VGND VGND VPWR VPWR _03392_ sky130_fd_sc_hd__a21bo_1
X_16073_ _06427_ _06429_ VGND VGND VPWR VPWR _06430_ sky130_fd_sc_hd__nor2_1
X_10497_ _00589_ VGND VGND VPWR VPWR _00590_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15024_ _05184_ _05185_ VGND VGND VPWR VPWR _05293_ sky130_fd_sc_hd__and2b_1
X_12236_ _02327_ _02328_ VGND VGND VPWR VPWR _02329_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_122_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12167_ _01106_ _01113_ _02259_ _00398_ VGND VGND VPWR VPWR _02260_ sky130_fd_sc_hd__or4b_4
X_11118_ _05595_ _04395_ _04886_ _05573_ VGND VGND VPWR VPWR _01211_ sky130_fd_sc_hd__a22o_1
X_12098_ _02086_ _02084_ VGND VGND VPWR VPWR _02191_ sky130_fd_sc_hd__or2_1
X_16975_ _00398_ _07311_ VGND VGND VPWR VPWR _07410_ sky130_fd_sc_hd__nand2_4
X_18714_ _09209_ _09241_ VGND VGND VPWR VPWR _09242_ sky130_fd_sc_hd__and2_1
XFILLER_0_36_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11049_ _01138_ _01140_ _01141_ VGND VGND VPWR VPWR _01142_ sky130_fd_sc_hd__and3_1
X_15926_ _06200_ _03011_ _06246_ _03154_ VGND VGND VPWR VPWR _06271_ sky130_fd_sc_hd__nand4_1
XFILLER_0_127_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput7 i_wb_addr[14] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__clkbuf_1
X_18645_ _06427_ _09190_ _09191_ VGND VGND VPWR VPWR _09192_ sky130_fd_sc_hd__a21oi_1
X_15857_ _03016_ _05652_ VGND VGND VPWR VPWR _06197_ sky130_fd_sc_hd__and2_1
X_14808_ _05034_ _05035_ _05055_ VGND VGND VPWR VPWR _05057_ sky130_fd_sc_hd__o21ai_1
X_18576_ _09097_ VGND VGND VPWR VPWR _09140_ sky130_fd_sc_hd__buf_2
X_15788_ _06121_ _06122_ VGND VGND VPWR VPWR _06123_ sky130_fd_sc_hd__and2_1
XFILLER_0_98_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17527_ _07887_ _07889_ _07885_ VGND VGND VPWR VPWR _08012_ sky130_fd_sc_hd__o21ba_1
X_14739_ _04979_ _04980_ VGND VGND VPWR VPWR _04981_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_87_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17458_ _06800_ _07934_ _07935_ VGND VGND VPWR VPWR _07936_ sky130_fd_sc_hd__a21o_1
X_16409_ _02974_ _03119_ _03534_ _06788_ _06794_ VGND VGND VPWR VPWR _06795_ sky130_fd_sc_hd__o311a_1
XFILLER_0_55_772 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17389_ _03107_ _07592_ VGND VGND VPWR VPWR _07861_ sky130_fd_sc_hd__nand2_4
XFILLER_0_27_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_125_660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_112_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09714_ _04690_ _05388_ VGND VGND VPWR VPWR _06395_ sky130_fd_sc_hd__nand2_1
X_09645_ _05638_ VGND VGND VPWR VPWR _05649_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_96_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09576_ _04088_ _03892_ _04886_ _03903_ VGND VGND VPWR VPWR _04897_ sky130_fd_sc_hd__and4_1
XTAP_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10420_ _09256_ VGND VGND VPWR VPWR _00513_ sky130_fd_sc_hd__buf_4
XFILLER_0_116_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10351_ _03728_ _00443_ VGND VGND VPWR VPWR _00444_ sky130_fd_sc_hd__nand2_1
XFILLER_0_131_630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13070_ _00517_ _03024_ VGND VGND VPWR VPWR _03162_ sky130_fd_sc_hd__and2_1
X_10282_ _00336_ _00372_ _00373_ _00374_ VGND VGND VPWR VPWR _00375_ sky130_fd_sc_hd__and4b_2
X_12021_ _02112_ _02113_ ApproximateM_inst.lob_16.lob2.genblk1\[5\].genblk1.mux.sel
+ _03432_ VGND VGND VPWR VPWR _02114_ sky130_fd_sc_hd__and4bb_1
X_16760_ _02533_ _06592_ _06551_ VGND VGND VPWR VPWR _07176_ sky130_fd_sc_hd__a21o_1
X_13972_ _04123_ _04124_ _04142_ VGND VGND VPWR VPWR _04144_ sky130_fd_sc_hd__o21a_1
X_15711_ _02991_ _03071_ _06037_ VGND VGND VPWR VPWR _06039_ sky130_fd_sc_hd__nand3_1
X_12923_ _03015_ VGND VGND VPWR VPWR _03016_ sky130_fd_sc_hd__clkbuf_4
X_16691_ _07081_ _07082_ _07100_ VGND VGND VPWR VPWR _07101_ sky130_fd_sc_hd__nand3_1
X_18430_ _06409_ _07274_ _08992_ _06720_ VGND VGND VPWR VPWR _08993_ sky130_fd_sc_hd__o211a_1
X_15642_ _05961_ _05963_ VGND VGND VPWR VPWR _05965_ sky130_fd_sc_hd__or2_1
XTAP_2230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12854_ _02945_ _02946_ VGND VGND VPWR VPWR _02947_ sky130_fd_sc_hd__and2_1
XTAP_2241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_706 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11805_ _01756_ _01896_ _01892_ _01895_ VGND VGND VPWR VPWR _01898_ sky130_fd_sc_hd__a211o_1
XTAP_2274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18361_ _08802_ _08870_ VGND VGND VPWR VPWR _08918_ sky130_fd_sc_hd__nor2_1
X_15573_ _05882_ _05889_ VGND VGND VPWR VPWR _05890_ sky130_fd_sc_hd__or2_1
XFILLER_0_69_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12785_ _02873_ _02877_ VGND VGND VPWR VPWR _02878_ sky130_fd_sc_hd__xnor2_1
XTAP_2296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17312_ _07772_ _07774_ _07775_ VGND VGND VPWR VPWR _07778_ sky130_fd_sc_hd__or3_1
X_14524_ _04745_ _04746_ VGND VGND VPWR VPWR _04747_ sky130_fd_sc_hd__nand2_1
XTAP_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11736_ ApproximateM_inst.lob_16.lob2.genblk1\[8\].genblk1.mux.sel _00210_ VGND VGND
+ VPWR VPWR _01829_ sky130_fd_sc_hd__and2_2
X_18292_ _00786_ _00787_ _07743_ _08774_ VGND VGND VPWR VPWR _08844_ sky130_fd_sc_hd__o31a_1
XFILLER_0_139_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_125_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17243_ _07666_ _07663_ VGND VGND VPWR VPWR _07702_ sky130_fd_sc_hd__or2b_1
XFILLER_0_154_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14455_ _04484_ _04670_ _04671_ VGND VGND VPWR VPWR _04672_ sky130_fd_sc_hd__or3_2
XFILLER_0_37_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11667_ _01757_ _01758_ _01201_ _01759_ VGND VGND VPWR VPWR _01760_ sky130_fd_sc_hd__o211a_1
XFILLER_0_153_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13406_ _03367_ _03369_ _03523_ _03524_ VGND VGND VPWR VPWR _03525_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_141_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10618_ _00709_ _00710_ VGND VGND VPWR VPWR _00711_ sky130_fd_sc_hd__xnor2_1
X_17174_ _07622_ _07625_ _07626_ VGND VGND VPWR VPWR _07627_ sky130_fd_sc_hd__and3_1
X_14386_ _04584_ _04585_ _04595_ VGND VGND VPWR VPWR _04596_ sky130_fd_sc_hd__o21ai_2
X_11598_ _01687_ _01688_ _01689_ VGND VGND VPWR VPWR _01691_ sky130_fd_sc_hd__a21o_1
XFILLER_0_141_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16125_ _03152_ _07766_ _03150_ VGND VGND VPWR VPWR _06486_ sky130_fd_sc_hd__nor3_1
XFILLER_0_141_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10549_ _06711_ _07733_ VGND VGND VPWR VPWR _00642_ sky130_fd_sc_hd__nand2_1
X_13337_ _03447_ _03448_ VGND VGND VPWR VPWR _03449_ sky130_fd_sc_hd__and2_1
XFILLER_0_122_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16056_ _03013_ _03073_ VGND VGND VPWR VPWR _06411_ sky130_fd_sc_hd__or2_1
X_13268_ net131 _03266_ _03291_ VGND VGND VPWR VPWR _03373_ sky130_fd_sc_hd__nor3_2
X_15007_ _01745_ _03142_ VGND VGND VPWR VPWR _05274_ sky130_fd_sc_hd__nand2_1
XFILLER_0_110_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12219_ _02308_ _02311_ VGND VGND VPWR VPWR _02312_ sky130_fd_sc_hd__and2b_1
X_13199_ _03298_ _03299_ VGND VGND VPWR VPWR _03300_ sky130_fd_sc_hd__nor2_1
XFILLER_0_138_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16958_ _06937_ _07332_ _07390_ _06542_ VGND VGND VPWR VPWR _07391_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_154_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15909_ _06251_ _06252_ VGND VGND VPWR VPWR _06253_ sky130_fd_sc_hd__nand2_1
X_16889_ _07124_ _07042_ _07313_ _06561_ VGND VGND VPWR VPWR _07316_ sky130_fd_sc_hd__o22a_1
X_09430_ _03281_ _03206_ _03260_ _03292_ VGND VGND VPWR VPWR _00001_ sky130_fd_sc_hd__a22o_1
XFILLER_0_149_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18628_ net314 _09097_ _09175_ _09176_ VGND VGND VPWR VPWR _00034_ sky130_fd_sc_hd__o211a_1
XFILLER_0_154_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18559_ net301 _09098_ _09129_ _09126_ VGND VGND VPWR VPWR _00005_ sky130_fd_sc_hd__o211a_1
XFILLER_0_19_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_12 _00644_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_23 _01115_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_644 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_34 _01355_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_45 _02917_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_56 _03760_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_67 _04649_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_78 _07123_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_89 _08880_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_466 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_112_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09628_ _05355_ VGND VGND VPWR VPWR _05464_ sky130_fd_sc_hd__buf_4
XFILLER_0_97_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09559_ _04690_ _04700_ VGND VGND VPWR VPWR _04711_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12570_ _02622_ _02659_ _02662_ VGND VGND VPWR VPWR _02663_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_65_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11521_ _01174_ _01612_ _01611_ VGND VGND VPWR VPWR _01614_ sky130_fd_sc_hd__a21o_1
XFILLER_0_108_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14240_ _04132_ _07015_ _07123_ _04099_ VGND VGND VPWR VPWR _04436_ sky130_fd_sc_hd__a22oi_1
X_11452_ _04548_ _00211_ _01541_ _01542_ VGND VGND VPWR VPWR _01545_ sky130_fd_sc_hd__a22o_1
XFILLER_0_34_775 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10403_ _00494_ _00495_ _00344_ _00343_ VGND VGND VPWR VPWR _00496_ sky130_fd_sc_hd__a31o_1
X_14171_ _09350_ _08409_ _00715_ _00112_ VGND VGND VPWR VPWR _04361_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_1_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11383_ _00877_ _00223_ _01428_ VGND VGND VPWR VPWR _01476_ sky130_fd_sc_hd__and3_1
XFILLER_0_21_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13122_ _05845_ _03215_ _03216_ VGND VGND VPWR VPWR _03218_ sky130_fd_sc_hd__a21bo_1
X_10334_ _09348_ _00273_ _00424_ _00426_ VGND VGND VPWR VPWR _00427_ sky130_fd_sc_hd__a211oi_4
XTAP_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13053_ _00861_ _03144_ _03023_ VGND VGND VPWR VPWR _03145_ sky130_fd_sc_hd__o21ai_1
X_17930_ _08366_ _08377_ VGND VGND VPWR VPWR _08450_ sky130_fd_sc_hd__or2_1
X_10265_ cla_inst.in2\[30\] VGND VGND VPWR VPWR _00358_ sky130_fd_sc_hd__buf_2
X_12004_ _02093_ _02096_ _02094_ VGND VGND VPWR VPWR _02097_ sky130_fd_sc_hd__o21ai_1
X_17861_ _08373_ _08374_ VGND VGND VPWR VPWR _08375_ sky130_fd_sc_hd__nor2_1
X_10196_ _00281_ _00287_ _00286_ VGND VGND VPWR VPWR _00289_ sky130_fd_sc_hd__a21o_1
X_16812_ _07133_ _07136_ VGND VGND VPWR VPWR _07233_ sky130_fd_sc_hd__and2b_1
X_17792_ _07207_ _07780_ _07623_ _06947_ VGND VGND VPWR VPWR _08301_ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16743_ _07154_ _07157_ VGND VGND VPWR VPWR _07158_ sky130_fd_sc_hd__xnor2_2
X_13955_ _03456_ VGND VGND VPWR VPWR _04125_ sky130_fd_sc_hd__buf_4
XFILLER_0_88_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12906_ _01745_ VGND VGND VPWR VPWR _02999_ sky130_fd_sc_hd__clkbuf_4
X_16674_ _06343_ _06997_ _06342_ VGND VGND VPWR VPWR _07083_ sky130_fd_sc_hd__a21oi_1
X_13886_ _04004_ _04005_ _04048_ _04049_ VGND VGND VPWR VPWR _04050_ sky130_fd_sc_hd__or4_4
X_18413_ _08840_ _08972_ _08974_ VGND VGND VPWR VPWR _08975_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_29_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15625_ _05945_ _05946_ VGND VGND VPWR VPWR _05947_ sky130_fd_sc_hd__nand2_1
XTAP_2060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12837_ _02928_ _02929_ VGND VGND VPWR VPWR _02930_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18344_ _08848_ _08899_ VGND VGND VPWR VPWR _08900_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_127_700 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15556_ _05781_ _05782_ _05784_ VGND VGND VPWR VPWR _05872_ sky130_fd_sc_hd__o21a_1
XTAP_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12768_ _02858_ _02859_ _01795_ _02854_ VGND VGND VPWR VPWR _02861_ sky130_fd_sc_hd__o211a_1
XFILLER_0_56_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14507_ _02188_ cla_inst.in1\[31\] VGND VGND VPWR VPWR _04728_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_686 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18275_ _01359_ _06593_ _06594_ VGND VGND VPWR VPWR _08826_ sky130_fd_sc_hd__a21o_1
X_11719_ _01783_ _01786_ _01751_ _01785_ VGND VGND VPWR VPWR _01812_ sky130_fd_sc_hd__a211o_1
XFILLER_0_126_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15487_ _05789_ _05796_ VGND VGND VPWR VPWR _05797_ sky130_fd_sc_hd__or2_1
XFILLER_0_25_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12699_ _02758_ _02791_ VGND VGND VPWR VPWR _02792_ sky130_fd_sc_hd__xor2_1
XFILLER_0_127_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17226_ _07680_ _07681_ _07682_ VGND VGND VPWR VPWR _07684_ sky130_fd_sc_hd__nand3_1
XFILLER_0_116_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_154_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput10 i_wb_addr[17] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__clkbuf_1
X_14438_ _00115_ _05921_ _04519_ _04518_ VGND VGND VPWR VPWR _04653_ sky130_fd_sc_hd__a31o_1
XFILLER_0_142_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput21 i_wb_addr[27] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_140_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput32 i_wb_addr[8] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput43 i_wb_data[17] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_114_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput54 i_wb_data[27] VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__buf_1
X_17157_ _07290_ VGND VGND VPWR VPWR _07608_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_142_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput65 i_wb_data[8] VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__buf_2
X_14369_ _04575_ _04576_ _04984_ _00498_ VGND VGND VPWR VPWR _04577_ sky130_fd_sc_hd__and4bb_2
X_16108_ _06466_ VGND VGND VPWR VPWR _06467_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_141_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17088_ _07507_ _07531_ _07532_ VGND VGND VPWR VPWR _07533_ sky130_fd_sc_hd__and3_1
XFILLER_0_12_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16039_ _03000_ _03044_ VGND VGND VPWR VPWR _06392_ sky130_fd_sc_hd__or2_1
XFILLER_0_110_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_118_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_140_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10050_ _08202_ _08148_ _08213_ _08235_ VGND VGND VPWR VPWR _00143_ sky130_fd_sc_hd__nor4_1
XFILLER_0_98_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13740_ _03507_ _03510_ _03718_ _03719_ VGND VGND VPWR VPWR _03890_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_97_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10952_ _04416_ _00949_ _03421_ _04340_ VGND VGND VPWR VPWR _01045_ sky130_fd_sc_hd__a22o_1
X_13671_ _03660_ _03665_ _03813_ VGND VGND VPWR VPWR _03814_ sky130_fd_sc_hd__a21bo_1
X_10883_ _00974_ _00975_ VGND VGND VPWR VPWR _00976_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_97_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15410_ _05711_ _05712_ _04238_ VGND VGND VPWR VPWR _05713_ sky130_fd_sc_hd__a21oi_1
X_12622_ _02677_ _02714_ VGND VGND VPWR VPWR _02715_ sky130_fd_sc_hd__xnor2_1
X_16390_ _06771_ _06773_ VGND VGND VPWR VPWR _06774_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_39_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15341_ _01356_ _00322_ _05633_ _05634_ VGND VGND VPWR VPWR _05637_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12553_ ApproximateM_inst.lob_16.lob2.mux.sel _00774_ VGND VGND VPWR VPWR _02646_
+ sky130_fd_sc_hd__and2_2
X_11504_ _05595_ _03903_ _03914_ _06019_ VGND VGND VPWR VPWR _01597_ sky130_fd_sc_hd__a22o_1
XFILLER_0_80_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18060_ _08586_ _08589_ _08591_ VGND VGND VPWR VPWR _08592_ sky130_fd_sc_hd__a21oi_2
X_15272_ _05446_ _05448_ _05561_ VGND VGND VPWR VPWR _05563_ sky130_fd_sc_hd__o21a_1
X_12484_ _02568_ _02569_ VGND VGND VPWR VPWR _02577_ sky130_fd_sc_hd__xor2_1
XFILLER_0_22_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17011_ _07447_ _07448_ VGND VGND VPWR VPWR _07449_ sky130_fd_sc_hd__and2b_1
X_14223_ _03539_ _04417_ VGND VGND VPWR VPWR _04418_ sky130_fd_sc_hd__nor2_1
X_11435_ _04362_ _00774_ _00909_ _04340_ VGND VGND VPWR VPWR _01528_ sky130_fd_sc_hd__a22o_1
XFILLER_0_124_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_734 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_767 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11366_ net142 _01457_ _01389_ _01387_ VGND VGND VPWR VPWR _01459_ sky130_fd_sc_hd__o211a_1
X_14154_ _01504_ _05888_ VGND VGND VPWR VPWR _04343_ sky130_fd_sc_hd__nand2_1
X_10317_ _00408_ _00409_ VGND VGND VPWR VPWR _00410_ sky130_fd_sc_hd__xor2_1
X_13105_ _03198_ VGND VGND VPWR VPWR _03199_ sky130_fd_sc_hd__clkbuf_4
X_14085_ _04097_ _04098_ VGND VGND VPWR VPWR _04267_ sky130_fd_sc_hd__and2b_1
XTAP_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11297_ _01387_ _01388_ _01383_ _01384_ VGND VGND VPWR VPWR _01390_ sky130_fd_sc_hd__a211o_1
X_18962_ clknet_4_6_0_clk _09392_ VGND VGND VPWR VPWR salida\[15\] sky130_fd_sc_hd__dfxtp_1
XTAP_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10248_ _08832_ _08854_ VGND VGND VPWR VPWR _00341_ sky130_fd_sc_hd__or2_1
XTAP_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17913_ _08427_ _08429_ _08430_ VGND VGND VPWR VPWR _08433_ sky130_fd_sc_hd__nand3_1
X_13036_ _03026_ _01503_ _02805_ VGND VGND VPWR VPWR _03128_ sky130_fd_sc_hd__a21o_1
X_18893_ clknet_4_11_0_clk _00047_ VGND VGND VPWR VPWR ApproximateM_inst.lob_16.lob1.genblk1\[11\].genblk1.mux.sel
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_119_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17844_ _06961_ _06957_ _07706_ _08260_ VGND VGND VPWR VPWR _08357_ sky130_fd_sc_hd__or4_1
X_10179_ _09344_ _09347_ _06938_ _08311_ VGND VGND VPWR VPWR _00272_ sky130_fd_sc_hd__o211ai_4
X_17775_ _07194_ _07318_ _07290_ _07313_ VGND VGND VPWR VPWR _08282_ sky130_fd_sc_hd__or4_2
X_14987_ _09352_ _05986_ _05249_ _05250_ VGND VGND VPWR VPWR _05252_ sky130_fd_sc_hd__o2bb2a_1
X_16726_ _07103_ _07138_ VGND VGND VPWR VPWR _07139_ sky130_fd_sc_hd__xnor2_1
X_13938_ _04100_ _04105_ VGND VGND VPWR VPWR _04106_ sky130_fd_sc_hd__xor2_1
XFILLER_0_135_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16657_ _06976_ _06978_ VGND VGND VPWR VPWR _07064_ sky130_fd_sc_hd__and2_1
X_13869_ _09349_ _03815_ _03837_ cla_inst.in2\[27\] VGND VGND VPWR VPWR _04031_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_29_300 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15608_ _05914_ _05926_ VGND VGND VPWR VPWR _05928_ sky130_fd_sc_hd__or2_1
XFILLER_0_60_10 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_147_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16588_ _02728_ _06509_ _03169_ VGND VGND VPWR VPWR _06989_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_57_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18327_ _03198_ _06152_ VGND VGND VPWR VPWR _08882_ sky130_fd_sc_hd__nand2_1
X_15539_ _05449_ _00119_ _05852_ _05849_ VGND VGND VPWR VPWR _05853_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_72_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18258_ _08804_ _08806_ VGND VGND VPWR VPWR _08807_ sky130_fd_sc_hd__nand2_1
XFILLER_0_60_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17209_ _07664_ VGND VGND VPWR VPWR _07665_ sky130_fd_sc_hd__buf_4
XFILLER_0_13_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18189_ _08654_ _08657_ _08652_ VGND VGND VPWR VPWR _08732_ sky130_fd_sc_hd__o21a_1
XFILLER_0_13_745 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_74 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09962_ _07363_ _07733_ VGND VGND VPWR VPWR _09091_ sky130_fd_sc_hd__nand2_1
XFILLER_0_110_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09893_ _03465_ _03815_ VGND VGND VPWR VPWR _08344_ sky130_fd_sc_hd__and2_1
XTAP_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_200 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_146_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_145_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11220_ _01093_ _01103_ VGND VGND VPWR VPWR _01313_ sky130_fd_sc_hd__or2b_1
XFILLER_0_105_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11151_ _01242_ VGND VGND VPWR VPWR _01244_ sky130_fd_sc_hd__inv_2
XFILLER_0_101_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10102_ _00184_ VGND VGND VPWR VPWR _00195_ sky130_fd_sc_hd__clkbuf_4
X_11082_ _01172_ _01174_ VGND VGND VPWR VPWR _01175_ sky130_fd_sc_hd__and2_1
X_14910_ _05038_ _05042_ _05040_ VGND VGND VPWR VPWR _05168_ sky130_fd_sc_hd__o21ba_1
X_10033_ _00109_ _00125_ _09212_ _09188_ VGND VGND VPWR VPWR _00126_ sky130_fd_sc_hd__and4_1
X_15890_ _06076_ _06079_ _06185_ _06231_ VGND VGND VPWR VPWR _06232_ sky130_fd_sc_hd__a211o_1
X_14841_ _05080_ _05081_ _05086_ _03125_ _05092_ VGND VGND VPWR VPWR _09358_ sky130_fd_sc_hd__a221o_1
X_17560_ _02124_ _07825_ VGND VGND VPWR VPWR _08047_ sky130_fd_sc_hd__nand2_1
X_14772_ _04910_ _04911_ VGND VGND VPWR VPWR _05018_ sky130_fd_sc_hd__or2_1
XFILLER_0_98_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11984_ _02073_ _02075_ _02076_ VGND VGND VPWR VPWR _02077_ sky130_fd_sc_hd__nor3_1
X_16511_ _02826_ _02827_ VGND VGND VPWR VPWR _06905_ sky130_fd_sc_hd__nor2_1
X_13723_ _03863_ _03871_ VGND VGND VPWR VPWR _03872_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_14_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10935_ _01026_ _01027_ VGND VGND VPWR VPWR _01028_ sky130_fd_sc_hd__xnor2_2
X_17491_ _07866_ _07873_ VGND VGND VPWR VPWR _07972_ sky130_fd_sc_hd__or2b_1
XFILLER_0_85_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16442_ _06654_ _06665_ _06829_ VGND VGND VPWR VPWR _06831_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_129_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13654_ _05508_ _05464_ _07722_ _08169_ VGND VGND VPWR VPWR _03796_ sky130_fd_sc_hd__nand4_2
X_10866_ _00957_ VGND VGND VPWR VPWR _00959_ sky130_fd_sc_hd__inv_2
XFILLER_0_66_450 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12605_ _02547_ _02546_ VGND VGND VPWR VPWR _02698_ sky130_fd_sc_hd__and2b_1
XPHY_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16373_ _06755_ VGND VGND VPWR VPWR _06756_ sky130_fd_sc_hd__clkbuf_4
XPHY_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13585_ _03718_ _03719_ _03507_ _03510_ VGND VGND VPWR VPWR _03721_ sky130_fd_sc_hd__o211ai_2
XPHY_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10797_ _08311_ _00855_ _00823_ _00854_ VGND VGND VPWR VPWR _00890_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_53_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18112_ _08646_ _08647_ VGND VGND VPWR VPWR _08649_ sky130_fd_sc_hd__or2_1
XPHY_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15324_ _05614_ _05618_ _04823_ VGND VGND VPWR VPWR _05620_ sky130_fd_sc_hd__o21a_1
XPHY_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12536_ _02593_ _02627_ VGND VGND VPWR VPWR _02629_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_121_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18043_ _08565_ _08571_ VGND VGND VPWR VPWR _08574_ sky130_fd_sc_hd__or2_1
X_15255_ _05541_ _05543_ VGND VGND VPWR VPWR _05544_ sky130_fd_sc_hd__or2_1
X_12467_ _02502_ _02559_ VGND VGND VPWR VPWR _02560_ sky130_fd_sc_hd__nor2_1
XFILLER_0_112_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14206_ _04228_ _04230_ VGND VGND VPWR VPWR _04400_ sky130_fd_sc_hd__nor2_2
XFILLER_0_111_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11418_ _09188_ _01509_ _01510_ VGND VGND VPWR VPWR _01511_ sky130_fd_sc_hd__a21bo_1
X_15186_ _09352_ _00318_ _05466_ _05467_ VGND VGND VPWR VPWR _05469_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_22_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12398_ _02421_ _02488_ _02490_ VGND VGND VPWR VPWR _02491_ sky130_fd_sc_hd__nor3_1
XFILLER_0_1_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14137_ _03014_ _00557_ _04321_ _04323_ VGND VGND VPWR VPWR _04324_ sky130_fd_sc_hd__a22oi_1
X_11349_ _01337_ _01377_ _01440_ _01441_ VGND VGND VPWR VPWR _01442_ sky130_fd_sc_hd__o211a_1
XFILLER_0_39_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18945_ clknet_4_2_0_clk _00099_ VGND VGND VPWR VPWR cla_inst.in2\[31\] sky130_fd_sc_hd__dfxtp_2
X_14068_ _03541_ _03545_ _03099_ VGND VGND VPWR VPWR _04249_ sky130_fd_sc_hd__mux2_1
X_13019_ _03026_ _03111_ _01963_ VGND VGND VPWR VPWR _03112_ sky130_fd_sc_hd__a21o_1
X_18876_ clknet_4_14_0_clk net315 VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_146_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17827_ _02985_ _06547_ _06550_ VGND VGND VPWR VPWR _08339_ sky130_fd_sc_hd__a21o_1
XFILLER_0_55_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17758_ _08261_ _08262_ VGND VGND VPWR VPWR _08263_ sky130_fd_sc_hd__nor2_1
XFILLER_0_77_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16709_ _07028_ _07029_ VGND VGND VPWR VPWR _07120_ sky130_fd_sc_hd__and2b_1
X_17689_ _07038_ _07745_ VGND VGND VPWR VPWR _08188_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_658 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_135_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_128_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_cap140 _01380_ VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__buf_1
XFILLER_0_41_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09945_ _08854_ _08897_ VGND VGND VPWR VPWR _08908_ sky130_fd_sc_hd__nor2_1
XFILLER_0_96_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09876_ _07015_ VGND VGND VPWR VPWR _08158_ sky130_fd_sc_hd__clkbuf_8
XTAP_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10720_ _05617_ VGND VGND VPWR VPWR _00813_ sky130_fd_sc_hd__inv_4
XTAP_1947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_623 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10651_ _00741_ _00742_ _00555_ _00698_ VGND VGND VPWR VPWR _00744_ sky130_fd_sc_hd__o211a_1
XFILLER_0_76_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10582_ _00666_ _00674_ VGND VGND VPWR VPWR _00675_ sky130_fd_sc_hd__xnor2_1
X_13370_ _03302_ _03303_ VGND VGND VPWR VPWR _03485_ sky130_fd_sc_hd__or2b_1
XFILLER_0_35_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12321_ _02401_ _02413_ VGND VGND VPWR VPWR _02414_ sky130_fd_sc_hd__or2_1
XFILLER_0_63_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15040_ _05304_ _05305_ _05309_ VGND VGND VPWR VPWR _09360_ sky130_fd_sc_hd__o21ai_1
X_12252_ _02343_ _02336_ _02342_ VGND VGND VPWR VPWR _02345_ sky130_fd_sc_hd__and3_1
XFILLER_0_31_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11203_ _00808_ _00807_ VGND VGND VPWR VPWR _01296_ sky130_fd_sc_hd__and2b_1
X_12183_ _02271_ _02273_ _02274_ _02270_ VGND VGND VPWR VPWR _02276_ sky130_fd_sc_hd__o31ai_1
X_11134_ _01222_ _01225_ _01226_ VGND VGND VPWR VPWR _01227_ sky130_fd_sc_hd__or3_1
X_16991_ _07426_ VGND VGND VPWR VPWR _07427_ sky130_fd_sc_hd__inv_2
XFILLER_0_101_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11065_ _01034_ _01033_ _01032_ VGND VGND VPWR VPWR _01158_ sky130_fd_sc_hd__a21o_1
X_18730_ _03161_ net46 _09251_ VGND VGND VPWR VPWR _09254_ sky130_fd_sc_hd__mux2_1
X_15942_ _06265_ _06269_ _06287_ VGND VGND VPWR VPWR _06289_ sky130_fd_sc_hd__or3_1
X_10016_ cla_inst.in2\[27\] VGND VGND VPWR VPWR _00109_ sky130_fd_sc_hd__buf_2
X_18661_ _09176_ _09203_ VGND VGND VPWR VPWR _09204_ sky130_fd_sc_hd__and2_1
X_15873_ _06171_ _06214_ VGND VGND VPWR VPWR _06215_ sky130_fd_sc_hd__xor2_1
X_17612_ _07974_ _07992_ _07991_ VGND VGND VPWR VPWR _08105_ sky130_fd_sc_hd__a21oi_1
X_14824_ _05071_ _05073_ _04961_ _04939_ VGND VGND VPWR VPWR _05075_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_99_862 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_116_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18592_ net291 _09140_ _09151_ _09144_ VGND VGND VPWR VPWR _00019_ sky130_fd_sc_hd__o211a_1
X_17543_ _06379_ _06377_ _06378_ VGND VGND VPWR VPWR _08030_ sky130_fd_sc_hd__nand3_1
X_14755_ _04862_ _04969_ _04997_ _04998_ VGND VGND VPWR VPWR _04999_ sky130_fd_sc_hd__o211ai_1
X_11967_ _02059_ _00357_ _07613_ _04034_ VGND VGND VPWR VPWR _02060_ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_759 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13706_ _03850_ _03852_ VGND VGND VPWR VPWR _03853_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_58_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17474_ _07950_ _07953_ VGND VGND VPWR VPWR _07954_ sky130_fd_sc_hd__xor2_1
X_10918_ _05497_ _01009_ _01010_ VGND VGND VPWR VPWR _01011_ sky130_fd_sc_hd__a21bo_1
X_14686_ _04884_ _04922_ _04923_ VGND VGND VPWR VPWR _04924_ sky130_fd_sc_hd__nand3_2
XFILLER_0_86_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11898_ _01987_ _01990_ VGND VGND VPWR VPWR _01991_ sky130_fd_sc_hd__and2b_1
X_16425_ sel_op\[0\] VGND VGND VPWR VPWR _06812_ sky130_fd_sc_hd__inv_4
XFILLER_0_117_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13637_ _04635_ _04427_ cla_inst.in1\[25\] cla_inst.in1\[24\] VGND VGND VPWR VPWR
+ _03777_ sky130_fd_sc_hd__and4_1
Xsplit70 _05311_ VGND VGND VPWR VPWR net233 sky130_fd_sc_hd__clkbuf_2
X_10849_ _03990_ _00211_ _00928_ _00927_ VGND VGND VPWR VPWR _00942_ sky130_fd_sc_hd__a31o_1
XFILLER_0_6_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16356_ _03027_ _00593_ _02373_ _02982_ VGND VGND VPWR VPWR _06737_ sky130_fd_sc_hd__a211o_1
X_13568_ _03440_ _03442_ VGND VGND VPWR VPWR _03702_ sky130_fd_sc_hd__or2_1
XFILLER_0_14_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15307_ _05459_ _05501_ _05457_ VGND VGND VPWR VPWR _05601_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_42_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12519_ _02609_ _02610_ _02611_ VGND VGND VPWR VPWR _02612_ sky130_fd_sc_hd__nand3_1
X_16287_ _00644_ net213 _06517_ VGND VGND VPWR VPWR _06662_ sky130_fd_sc_hd__or3_1
X_13499_ _06029_ _05649_ cla_inst.in1\[30\] _07755_ VGND VGND VPWR VPWR _03626_ sky130_fd_sc_hd__and4_1
XFILLER_0_2_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18026_ _08553_ _08554_ VGND VGND VPWR VPWR _08555_ sky130_fd_sc_hd__xor2_2
X_15238_ _05510_ _05511_ _05514_ VGND VGND VPWR VPWR _05525_ sky130_fd_sc_hd__or3b_1
XFILLER_0_41_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15169_ _05449_ _03044_ _05447_ VGND VGND VPWR VPWR _05450_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_10_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_4_7_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_7_0_clk sky130_fd_sc_hd__clkbuf_8
X_09730_ _05126_ _05115_ VGND VGND VPWR VPWR _06569_ sky130_fd_sc_hd__or2b_1
X_18928_ clknet_4_8_0_clk _00082_ VGND VGND VPWR VPWR ApproximateM_inst.lob_16.lob2.genblk1\[14\].genblk1.mux.sel
+ sky130_fd_sc_hd__dfxtp_1
X_09661_ _05192_ _05203_ _05802_ VGND VGND VPWR VPWR _05823_ sky130_fd_sc_hd__and3_1
X_18859_ clknet_4_4_0_clk net258 VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__dfxtp_1
X_09592_ _04635_ _04427_ _04569_ _04449_ VGND VGND VPWR VPWR _05072_ sky130_fd_sc_hd__and4_1
XFILLER_0_96_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_119_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_842 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_114 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_131_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_591 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09928_ _08713_ VGND VGND VPWR VPWR _08724_ sky130_fd_sc_hd__clkbuf_8
X_09859_ ApproximateM_inst.lob_16.lob2.genblk1\[3\].genblk1.mux.sel VGND VGND VPWR
+ VPWR _07973_ sky130_fd_sc_hd__buf_6
X_12870_ _02959_ _02962_ VGND VGND VPWR VPWR _02963_ sky130_fd_sc_hd__nand2_2
XFILLER_0_99_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_102 _09398_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_113 net49 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11821_ _01814_ VGND VGND VPWR VPWR _01914_ sky130_fd_sc_hd__inv_2
XFILLER_0_96_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_124 _02987_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_135 _05856_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_146 _08674_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_157 _08762_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14540_ _04762_ _04763_ VGND VGND VPWR VPWR _04764_ sky130_fd_sc_hd__xnor2_1
XTAP_1733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11752_ _01658_ _01666_ VGND VGND VPWR VPWR _01845_ sky130_fd_sc_hd__xnor2_1
XTAP_1744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_168 _05410_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_179 _02646_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10703_ _04318_ _04755_ _04744_ VGND VGND VPWR VPWR _00796_ sky130_fd_sc_hd__a21oi_2
XTAP_1777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14471_ _04544_ _04546_ VGND VGND VPWR VPWR _04689_ sky130_fd_sc_hd__nor2_1
XTAP_1788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11683_ _01733_ _01772_ _01775_ VGND VGND VPWR VPWR _01776_ sky130_fd_sc_hd__o21a_1
XTAP_1799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16210_ _06573_ _06577_ _01106_ VGND VGND VPWR VPWR _06578_ sky130_fd_sc_hd__a21o_1
XFILLER_0_138_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13422_ _03540_ _03541_ _03061_ VGND VGND VPWR VPWR _03543_ sky130_fd_sc_hd__mux2_1
X_10634_ _00109_ _09349_ _03618_ _00171_ VGND VGND VPWR VPWR _00727_ sky130_fd_sc_hd__and4_1
X_17190_ _07484_ _07506_ _07533_ VGND VGND VPWR VPWR _07644_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_36_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16141_ _03099_ _06498_ _06502_ VGND VGND VPWR VPWR _06503_ sky130_fd_sc_hd__a21oi_1
X_13353_ _03434_ _03435_ _03466_ VGND VGND VPWR VPWR _03467_ sky130_fd_sc_hd__or3_4
X_10565_ _00655_ _00656_ _00636_ _00637_ VGND VGND VPWR VPWR _00658_ sky130_fd_sc_hd__a211o_1
XFILLER_0_107_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12304_ _02392_ _02395_ _02311_ _02396_ VGND VGND VPWR VPWR _02397_ sky130_fd_sc_hd__o211a_1
XFILLER_0_133_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16072_ _07646_ _09354_ VGND VGND VPWR VPWR _06429_ sky130_fd_sc_hd__nand2_1
XFILLER_0_106_385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13284_ _03382_ _03383_ _03389_ VGND VGND VPWR VPWR _03391_ sky130_fd_sc_hd__a21o_1
X_10496_ _00427_ _00430_ _00587_ _00588_ VGND VGND VPWR VPWR _00589_ sky130_fd_sc_hd__o211a_1
XFILLER_0_122_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15023_ _05180_ _05291_ VGND VGND VPWR VPWR _05292_ sky130_fd_sc_hd__xnor2_2
X_12235_ _02163_ _02161_ VGND VGND VPWR VPWR _02328_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_121_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12166_ _04864_ VGND VGND VPWR VPWR _02259_ sky130_fd_sc_hd__clkinv_4
X_11117_ _07352_ _05322_ _01127_ _01128_ VGND VGND VPWR VPWR _01210_ sky130_fd_sc_hd__a22o_1
X_12097_ _02189_ VGND VGND VPWR VPWR _02190_ sky130_fd_sc_hd__inv_2
X_16974_ _07196_ _07197_ _07294_ VGND VGND VPWR VPWR _07409_ sky130_fd_sc_hd__and3_1
X_18713_ net55 _06408_ _09182_ VGND VGND VPWR VPWR _09241_ sky130_fd_sc_hd__mux2_1
X_11048_ _01109_ _01137_ VGND VGND VPWR VPWR _01141_ sky130_fd_sc_hd__or2_1
X_15925_ _03011_ _06246_ _03154_ _06200_ VGND VGND VPWR VPWR _06270_ sky130_fd_sc_hd__a22o_1
Xinput8 i_wb_addr[15] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__clkbuf_1
X_18644_ net69 VGND VGND VPWR VPWR _09191_ sky130_fd_sc_hd__buf_2
X_15856_ _06194_ _06195_ VGND VGND VPWR VPWR _06196_ sky130_fd_sc_hd__nand2_1
XFILLER_0_99_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14807_ _05034_ _05035_ _05055_ VGND VGND VPWR VPWR _05056_ sky130_fd_sc_hd__or3_2
XFILLER_0_99_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15787_ _06053_ _06055_ _06120_ VGND VGND VPWR VPWR _06122_ sky130_fd_sc_hd__or3_1
X_18575_ net277 _09098_ _09139_ _09126_ VGND VGND VPWR VPWR _00013_ sky130_fd_sc_hd__o211a_1
X_12999_ _03025_ _00881_ _02646_ VGND VGND VPWR VPWR _03092_ sky130_fd_sc_hd__a21o_1
X_17526_ _08009_ _08010_ VGND VGND VPWR VPWR _08011_ sky130_fd_sc_hd__or2_1
X_14738_ _02059_ _03455_ VGND VGND VPWR VPWR _04980_ sky130_fd_sc_hd__nand2_1
XFILLER_0_143_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_146_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17457_ _06755_ _07621_ _07933_ net331 VGND VGND VPWR VPWR _07935_ sky130_fd_sc_hd__o22a_1
X_14669_ _04780_ _04787_ VGND VGND VPWR VPWR _04905_ sky130_fd_sc_hd__and2_1
XFILLER_0_145_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16408_ _03083_ _06789_ _06793_ VGND VGND VPWR VPWR _06794_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_116_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17388_ _07038_ _07649_ _07859_ _06527_ VGND VGND VPWR VPWR _07860_ sky130_fd_sc_hd__a22o_1
X_16339_ _03539_ _06705_ _06712_ _06718_ _06484_ VGND VGND VPWR VPWR _06719_ sky130_fd_sc_hd__o221a_1
XFILLER_0_42_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18009_ _07390_ _07650_ VGND VGND VPWR VPWR _08536_ sky130_fd_sc_hd__nand2_1
XFILLER_0_140_664 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_74 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09713_ _04853_ _04875_ _04897_ VGND VGND VPWR VPWR _06384_ sky130_fd_sc_hd__o21ba_1
X_09644_ ApproximateM_inst.lob_16.lob2.genblk1\[6\].genblk1.mux.sel VGND VGND VPWR
+ VPWR _05638_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_97_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09575_ _03739_ VGND VGND VPWR VPWR _04886_ sky130_fd_sc_hd__clkbuf_4
XTAP_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_879 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10350_ _05333_ VGND VGND VPWR VPWR _00443_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_5_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10281_ _00333_ _00335_ _08681_ _09005_ VGND VGND VPWR VPWR _00374_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_130_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12020_ _05638_ _04220_ _00217_ _00992_ VGND VGND VPWR VPWR _02113_ sky130_fd_sc_hd__a22oi_1
X_13971_ _04127_ _04141_ VGND VGND VPWR VPWR _04142_ sky130_fd_sc_hd__xnor2_2
X_15710_ _02991_ _00495_ _06037_ VGND VGND VPWR VPWR _06038_ sky130_fd_sc_hd__a21o_1
X_12922_ _03014_ VGND VGND VPWR VPWR _03015_ sky130_fd_sc_hd__buf_2
X_16690_ _07083_ _07085_ _07093_ _07099_ VGND VGND VPWR VPWR _07100_ sky130_fd_sc_hd__o211a_1
X_15641_ _03015_ _03067_ _05962_ _05959_ VGND VGND VPWR VPWR _05963_ sky130_fd_sc_hd__o2bb2a_1
X_12853_ _02943_ _02944_ _02926_ _02928_ VGND VGND VPWR VPWR _02946_ sky130_fd_sc_hd__o211ai_2
XTAP_2220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11804_ _01892_ _01895_ _01756_ _01896_ VGND VGND VPWR VPWR _01897_ sky130_fd_sc_hd__o211ai_2
XTAP_2264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18360_ _08915_ _08916_ VGND VGND VPWR VPWR _08917_ sky130_fd_sc_hd__and2_1
X_15572_ _05885_ _05887_ VGND VGND VPWR VPWR _05889_ sky130_fd_sc_hd__or2_1
XTAP_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12784_ _02875_ _02876_ VGND VGND VPWR VPWR _02877_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_84_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17311_ _07772_ _07774_ _07775_ VGND VGND VPWR VPWR _07776_ sky130_fd_sc_hd__o21a_1
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14523_ _00679_ _00678_ _01575_ _00715_ VGND VGND VPWR VPWR _04746_ sky130_fd_sc_hd__nand4_1
XFILLER_0_68_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11735_ _01820_ _01826_ _01827_ VGND VGND VPWR VPWR _01828_ sky130_fd_sc_hd__a21o_2
XFILLER_0_127_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18291_ _08797_ _08796_ VGND VGND VPWR VPWR _08842_ sky130_fd_sc_hd__or2b_1
XFILLER_0_154_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17242_ _07662_ _07661_ VGND VGND VPWR VPWR _07701_ sky130_fd_sc_hd__or2b_1
X_14454_ _04667_ _04669_ _04649_ VGND VGND VPWR VPWR _04671_ sky130_fd_sc_hd__o21a_1
XFILLER_0_22_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11666_ _01198_ _01199_ _01200_ _01181_ VGND VGND VPWR VPWR _01759_ sky130_fd_sc_hd__a22o_1
XFILLER_0_36_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13405_ _03521_ _03522_ _03370_ _03347_ VGND VGND VPWR VPWR _03524_ sky130_fd_sc_hd__o211a_1
X_10617_ _00204_ _00557_ VGND VGND VPWR VPWR _00710_ sky130_fd_sc_hd__nand2_1
X_17173_ _06581_ _07511_ VGND VGND VPWR VPWR _07626_ sky130_fd_sc_hd__nor2_1
X_14385_ _04586_ _04594_ VGND VGND VPWR VPWR _04595_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_153_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11597_ _01687_ _01688_ _01689_ VGND VGND VPWR VPWR _01690_ sky130_fd_sc_hd__nand3_1
XFILLER_0_24_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16124_ _00517_ _03156_ VGND VGND VPWR VPWR _06485_ sky130_fd_sc_hd__nor2_1
X_13336_ _03439_ _03446_ VGND VGND VPWR VPWR _03448_ sky130_fd_sc_hd__nand2_1
X_10548_ _00639_ _00640_ VGND VGND VPWR VPWR _00641_ sky130_fd_sc_hd__nor2_1
XFILLER_0_106_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16055_ _06330_ _06407_ _06409_ _06024_ VGND VGND VPWR VPWR _06410_ sky130_fd_sc_hd__a211oi_2
X_13267_ _03341_ VGND VGND VPWR VPWR _03372_ sky130_fd_sc_hd__inv_2
X_10479_ _00560_ _00561_ _00571_ VGND VGND VPWR VPWR _00572_ sky130_fd_sc_hd__o21ai_1
X_15006_ _05271_ _05272_ VGND VGND VPWR VPWR _05273_ sky130_fd_sc_hd__nand2_1
X_12218_ _02309_ _02308_ _02310_ VGND VGND VPWR VPWR _02311_ sky130_fd_sc_hd__or3_1
XFILLER_0_20_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13198_ _00189_ _00191_ _04045_ _04067_ VGND VGND VPWR VPWR _03299_ sky130_fd_sc_hd__and4_1
XFILLER_0_20_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12149_ _07036_ _07069_ _00210_ _03607_ VGND VGND VPWR VPWR _02242_ sky130_fd_sc_hd__and4_1
XFILLER_0_138_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16957_ _07389_ VGND VGND VPWR VPWR _07390_ sky130_fd_sc_hd__clkbuf_4
X_15908_ _03007_ _03072_ _06249_ _06250_ VGND VGND VPWR VPWR _06252_ sky130_fd_sc_hd__a211o_1
XFILLER_0_154_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16888_ _06561_ _07124_ _07042_ _07314_ VGND VGND VPWR VPWR _07315_ sky130_fd_sc_hd__nor4_1
X_18627_ _09124_ VGND VGND VPWR VPWR _09176_ sky130_fd_sc_hd__buf_4
X_15839_ _06121_ _06124_ _06177_ VGND VGND VPWR VPWR _06178_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_63_87 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18558_ salida\[1\] _09114_ _09118_ salida\[33\] _09128_ VGND VGND VPWR VPWR _09129_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_86_161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17509_ _07975_ _07976_ _07990_ VGND VGND VPWR VPWR _07992_ sky130_fd_sc_hd__or3b_1
XFILLER_0_47_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18489_ _09018_ _09021_ _09052_ _09053_ _09019_ VGND VGND VPWR VPWR _09056_ sky130_fd_sc_hd__o2111a_1
XANTENNA_13 _00813_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_24 _01115_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_35 _01355_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_656 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_46 _02917_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_57 _04074_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_68 _04679_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_79 _07591_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_112_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09627_ _05279_ VGND VGND VPWR VPWR _05453_ sky130_fd_sc_hd__buf_4
XFILLER_0_69_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09558_ _04384_ VGND VGND VPWR VPWR _04700_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_84_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09489_ _03760_ _03935_ VGND VGND VPWR VPWR _03946_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_66_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11520_ _01174_ _01611_ _01612_ VGND VGND VPWR VPWR _01613_ sky130_fd_sc_hd__and3_1
XFILLER_0_93_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11451_ _03990_ _00146_ _01515_ _01509_ _00197_ VGND VGND VPWR VPWR _01544_ sky130_fd_sc_hd__a32o_1
XFILLER_0_34_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10402_ _09311_ VGND VGND VPWR VPWR _00495_ sky130_fd_sc_hd__buf_4
X_14170_ net219 _04155_ VGND VGND VPWR VPWR _04360_ sky130_fd_sc_hd__nor2_1
XFILLER_0_34_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11382_ _01426_ _01427_ VGND VGND VPWR VPWR _01475_ sky130_fd_sc_hd__and2b_1
XFILLER_0_21_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13121_ _04121_ _05322_ _05333_ _04088_ VGND VGND VPWR VPWR _03216_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10333_ _00421_ _00422_ _00425_ _00378_ VGND VGND VPWR VPWR _00426_ sky130_fd_sc_hd__o2bb2a_1
X_13052_ _03025_ _03143_ VGND VGND VPWR VPWR _03144_ sky130_fd_sc_hd__and2_1
X_10264_ _07570_ VGND VGND VPWR VPWR _00357_ sky130_fd_sc_hd__buf_6
X_12003_ _02094_ _02095_ VGND VGND VPWR VPWR _02096_ sky130_fd_sc_hd__nand2_1
X_10195_ _00281_ _00286_ _00287_ VGND VGND VPWR VPWR _00288_ sky130_fd_sc_hd__nand3_1
X_17860_ _08269_ _08271_ _08372_ VGND VGND VPWR VPWR _08374_ sky130_fd_sc_hd__and3_1
XFILLER_0_100_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16811_ _07229_ _07230_ VGND VGND VPWR VPWR _07231_ sky130_fd_sc_hd__nand2_1
XFILLER_0_108_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17791_ _07302_ _07303_ _07511_ _07621_ VGND VGND VPWR VPWR _08299_ sky130_fd_sc_hd__or4_1
XFILLER_0_17_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13954_ _04120_ _04122_ _03949_ _04091_ VGND VGND VPWR VPWR _04124_ sky130_fd_sc_hd__a211oi_4
X_16742_ _06973_ net205 _07155_ VGND VGND VPWR VPWR _07157_ sky130_fd_sc_hd__a21oi_2
X_12905_ _01505_ VGND VGND VPWR VPWR _02998_ sky130_fd_sc_hd__clkbuf_4
X_16673_ _02975_ _03916_ _03120_ _04243_ VGND VGND VPWR VPWR _07082_ sky130_fd_sc_hd__or4_1
X_13885_ _04046_ _04047_ _04006_ _03877_ VGND VGND VPWR VPWR _04049_ sky130_fd_sc_hd__o211a_1
XFILLER_0_88_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18412_ _08917_ _08918_ _08921_ _08893_ VGND VGND VPWR VPWR _08974_ sky130_fd_sc_hd__a22o_1
X_12836_ _02926_ _02927_ _02901_ _02922_ VGND VGND VPWR VPWR _02929_ sky130_fd_sc_hd__a211o_1
X_15624_ _05866_ _05870_ _05944_ VGND VGND VPWR VPWR _05946_ sky130_fd_sc_hd__or3_1
XTAP_2050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15555_ _05868_ _05869_ _05752_ VGND VGND VPWR VPWR _05871_ sky130_fd_sc_hd__a21oi_1
XTAP_2094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18343_ _07592_ _08896_ _08898_ VGND VGND VPWR VPWR _08899_ sky130_fd_sc_hd__nand3_1
XTAP_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12767_ _01795_ _02854_ _02858_ _02859_ VGND VGND VPWR VPWR _02860_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_29_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_712 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14506_ _04515_ cla_inst.in1\[30\] VGND VGND VPWR VPWR _04727_ sky130_fd_sc_hd__nand2_1
XTAP_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11718_ _01751_ _01785_ _01783_ _01786_ VGND VGND VPWR VPWR _01811_ sky130_fd_sc_hd__o211ai_2
X_18274_ _03056_ _06447_ VGND VGND VPWR VPWR _08825_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_154_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15486_ _05416_ _05793_ _05795_ VGND VGND VPWR VPWR _05796_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_84_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12698_ _02759_ _02789_ _02790_ VGND VGND VPWR VPWR _02791_ sky130_fd_sc_hd__and3_1
XFILLER_0_154_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14437_ _04514_ _04522_ VGND VGND VPWR VPWR _04652_ sky130_fd_sc_hd__and2_1
X_17225_ _07680_ _07681_ _07682_ VGND VGND VPWR VPWR _07683_ sky130_fd_sc_hd__a21o_1
Xinput11 i_wb_addr[18] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__clkbuf_1
X_11649_ _00164_ _01357_ _01680_ VGND VGND VPWR VPWR _01742_ sky130_fd_sc_hd__and3_1
Xinput22 i_wb_addr[28] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_114_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_142_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput33 i_wb_addr[9] VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput44 i_wb_data[18] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__clkbuf_2
X_17156_ _06969_ _07109_ VGND VGND VPWR VPWR _07607_ sky130_fd_sc_hd__nand2_1
X_14368_ _03881_ _03892_ cla_inst.in1\[27\] _07004_ VGND VGND VPWR VPWR _04576_ sky130_fd_sc_hd__and4_4
Xinput55 i_wb_data[28] VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__buf_1
Xinput66 i_wb_data[9] VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__buf_2
XFILLER_0_141_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16107_ _02728_ _03022_ VGND VGND VPWR VPWR _06466_ sky130_fd_sc_hd__and2b_1
X_13319_ _03428_ VGND VGND VPWR VPWR _03429_ sky130_fd_sc_hd__inv_2
XFILLER_0_40_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17087_ _07508_ _07509_ _07530_ VGND VGND VPWR VPWR _07532_ sky130_fd_sc_hd__or3_1
XFILLER_0_150_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14299_ _04499_ _04500_ VGND VGND VPWR VPWR _04501_ sky130_fd_sc_hd__or2b_1
X_16038_ _06389_ _06390_ _04421_ VGND VGND VPWR VPWR _06391_ sky130_fd_sc_hd__a21o_1
XFILLER_0_58_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17989_ _08512_ _08513_ _08514_ VGND VGND VPWR VPWR _08515_ sky130_fd_sc_hd__nand3_1
XFILLER_0_74_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_358 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_643 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_114_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_420 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_117_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_90 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_98_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10951_ _01040_ _01043_ VGND VGND VPWR VPWR _01044_ sky130_fd_sc_hd__xor2_2
XFILLER_0_98_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13670_ _03661_ _03664_ VGND VGND VPWR VPWR _03813_ sky130_fd_sc_hd__nand2_1
XFILLER_0_57_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10882_ _08615_ _00557_ _00945_ _00944_ VGND VGND VPWR VPWR _00975_ sky130_fd_sc_hd__a31o_2
X_12621_ _07602_ _02676_ _02678_ VGND VGND VPWR VPWR _02714_ sky130_fd_sc_hd__a21bo_1
X_15340_ _05635_ VGND VGND VPWR VPWR _05636_ sky130_fd_sc_hd__inv_2
XFILLER_0_109_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12552_ _02635_ _02642_ _02641_ VGND VGND VPWR VPWR _02645_ sky130_fd_sc_hd__a21o_1
XFILLER_0_66_687 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_136_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11503_ _05573_ _05595_ _03903_ VGND VGND VPWR VPWR _01596_ sky130_fd_sc_hd__and3_1
X_15271_ _05557_ _05560_ VGND VGND VPWR VPWR _05561_ sky130_fd_sc_hd__xor2_1
X_12483_ _02574_ _02575_ VGND VGND VPWR VPWR _02576_ sky130_fd_sc_hd__and2_1
XFILLER_0_80_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17010_ _07445_ _07446_ _07379_ _07380_ VGND VGND VPWR VPWR _07448_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_123_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14222_ _03063_ _03115_ _03916_ VGND VGND VPWR VPWR _04417_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11434_ _04504_ _04427_ _00217_ _00909_ VGND VGND VPWR VPWR _01527_ sky130_fd_sc_hd__nand4_2
XFILLER_0_22_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14153_ _04339_ _04341_ VGND VGND VPWR VPWR _04342_ sky130_fd_sc_hd__nor2_1
X_11365_ _01387_ _01389_ _01457_ net142 VGND VGND VPWR VPWR _01458_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_132_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_779 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13104_ _03197_ VGND VGND VPWR VPWR _03198_ sky130_fd_sc_hd__clkbuf_4
X_10316_ _00253_ _00213_ _00256_ _00255_ VGND VGND VPWR VPWR _00409_ sky130_fd_sc_hd__a31o_1
X_14084_ _04107_ _04108_ _04119_ VGND VGND VPWR VPWR _04266_ sky130_fd_sc_hd__nor3_1
X_18961_ clknet_4_6_0_clk _09391_ VGND VGND VPWR VPWR salida\[14\] sky130_fd_sc_hd__dfxtp_1
X_11296_ _01383_ _01384_ _01387_ _01388_ VGND VGND VPWR VPWR _01389_ sky130_fd_sc_hd__o211ai_4
XTAP_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17912_ _08427_ _08429_ _08430_ VGND VGND VPWR VPWR _08432_ sky130_fd_sc_hd__a21o_1
X_13035_ _03023_ _03126_ VGND VGND VPWR VPWR _03127_ sky130_fd_sc_hd__nand2_1
X_10247_ _06993_ _00339_ _09112_ _09101_ VGND VGND VPWR VPWR _00340_ sky130_fd_sc_hd__a31o_1
X_18892_ clknet_4_11_0_clk _00046_ VGND VGND VPWR VPWR ApproximateM_inst.lob_16.lob1.genblk1\[10\].genblk1.mux.sel
+ sky130_fd_sc_hd__dfxtp_1
X_17843_ _08353_ _08355_ VGND VGND VPWR VPWR _08356_ sky130_fd_sc_hd__xor2_1
X_10178_ _00268_ _00269_ _00161_ _00231_ VGND VGND VPWR VPWR _00271_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_89_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17774_ net146 _07604_ _07664_ _07394_ VGND VGND VPWR VPWR _08281_ sky130_fd_sc_hd__a22o_1
X_14986_ _05249_ _05250_ _09352_ _05975_ VGND VGND VPWR VPWR _05251_ sky130_fd_sc_hd__and4bb_1
X_16725_ _07111_ _07137_ VGND VGND VPWR VPWR _07138_ sky130_fd_sc_hd__xor2_1
X_13937_ _04103_ _04104_ VGND VGND VPWR VPWR _04105_ sky130_fd_sc_hd__xnor2_1
X_13868_ _03818_ _03820_ VGND VGND VPWR VPWR _04030_ sky130_fd_sc_hd__nor2_1
X_16656_ _06973_ _07062_ VGND VGND VPWR VPWR _07063_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_76_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_312 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12819_ _02909_ _02910_ _02896_ _02897_ VGND VGND VPWR VPWR _02912_ sky130_fd_sc_hd__o211ai_2
X_15607_ _05914_ _05926_ VGND VGND VPWR VPWR _05927_ sky130_fd_sc_hd__nand2_1
XFILLER_0_146_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13799_ _04340_ _04416_ cla_inst.in1\[26\] cla_inst.in1\[25\] VGND VGND VPWR VPWR
+ _03954_ sky130_fd_sc_hd__and4_2
X_16587_ _03169_ _06673_ VGND VGND VPWR VPWR _06988_ sky130_fd_sc_hd__nor2_1
XFILLER_0_60_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18326_ _03056_ _06447_ _03143_ VGND VGND VPWR VPWR _08881_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_139_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_151_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15538_ _05850_ VGND VGND VPWR VPWR _05852_ sky130_fd_sc_hd__inv_2
XTAP_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15469_ _05774_ _05775_ _05716_ _05695_ VGND VGND VPWR VPWR _05777_ sky130_fd_sc_hd__o211a_1
X_18257_ _08655_ _08733_ _08805_ VGND VGND VPWR VPWR _08806_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_4_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17208_ _00247_ _07311_ _07312_ VGND VGND VPWR VPWR _07664_ sky130_fd_sc_hd__and3_2
XFILLER_0_13_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18188_ _08729_ _08730_ VGND VGND VPWR VPWR _08731_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_130_707 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17139_ _07496_ _07505_ VGND VGND VPWR VPWR _07588_ sky130_fd_sc_hd__nor2_1
XFILLER_0_69_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09961_ _06678_ _06743_ VGND VGND VPWR VPWR _09080_ sky130_fd_sc_hd__or2_2
XFILLER_0_0_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09892_ _03629_ _03596_ _04657_ _03837_ VGND VGND VPWR VPWR _08333_ sky130_fd_sc_hd__nand4_2
XTAP_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_142 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_827 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_304 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_359 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_247 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_121_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11150_ _01241_ _01242_ cla_inst.in2\[21\] _09219_ VGND VGND VPWR VPWR _01243_ sky130_fd_sc_hd__and4b_1
XFILLER_0_101_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10101_ _00178_ VGND VGND VPWR VPWR _00194_ sky130_fd_sc_hd__buf_6
X_11081_ _05017_ _00165_ _01172_ _01173_ VGND VGND VPWR VPWR _01174_ sky130_fd_sc_hd__nand4_1
X_10032_ cla_inst.in2\[26\] VGND VGND VPWR VPWR _00125_ sky130_fd_sc_hd__clkbuf_4
X_14840_ _05090_ _05091_ _03199_ VGND VGND VPWR VPWR _05092_ sky130_fd_sc_hd__o21a_1
X_14771_ _04750_ _04915_ VGND VGND VPWR VPWR _05016_ sky130_fd_sc_hd__nor2_1
X_11983_ _02071_ _02072_ _02067_ _02070_ VGND VGND VPWR VPWR _02076_ sky130_fd_sc_hd__o211a_1
X_13722_ _03864_ _03869_ VGND VGND VPWR VPWR _03871_ sky130_fd_sc_hd__xor2_1
XFILLER_0_86_716 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16510_ _06834_ _06901_ _06903_ _06559_ VGND VGND VPWR VPWR _06904_ sky130_fd_sc_hd__a211o_1
XFILLER_0_58_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10934_ _03990_ _03618_ VGND VGND VPWR VPWR _01027_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17490_ _07872_ _07871_ VGND VGND VPWR VPWR _07971_ sky130_fd_sc_hd__or2b_1
X_13653_ _05366_ cla_inst.in1\[28\] _07374_ _05410_ VGND VGND VPWR VPWR _03795_ sky130_fd_sc_hd__a22o_1
X_16441_ _06771_ _06773_ VGND VGND VPWR VPWR _06829_ sky130_fd_sc_hd__or2b_1
X_10865_ _00956_ _00957_ _03717_ _03410_ VGND VGND VPWR VPWR _00958_ sky130_fd_sc_hd__and4b_1
XFILLER_0_128_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12604_ _08865_ _01503_ VGND VGND VPWR VPWR _02697_ sky130_fd_sc_hd__nand2_1
XPHY_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_602 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_109_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16372_ _02977_ _06753_ VGND VGND VPWR VPWR _06755_ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_164 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13584_ _03507_ _03510_ _03718_ _03719_ VGND VGND VPWR VPWR _03720_ sky130_fd_sc_hd__a211o_1
X_10796_ _00859_ _00888_ VGND VGND VPWR VPWR _00889_ sky130_fd_sc_hd__xnor2_2
XPHY_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15323_ _05614_ _05618_ VGND VGND VPWR VPWR _05619_ sky130_fd_sc_hd__nand2_1
XFILLER_0_93_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18111_ _08635_ _08645_ VGND VGND VPWR VPWR _08647_ sky130_fd_sc_hd__nor2_1
XPHY_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12535_ _02593_ _02627_ VGND VGND VPWR VPWR _02628_ sky130_fd_sc_hd__or2b_1
XPHY_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15254_ _05449_ _01139_ _05542_ _05538_ VGND VGND VPWR VPWR _05543_ sky130_fd_sc_hd__o2bb2a_1
X_18042_ _08565_ _08571_ VGND VGND VPWR VPWR _08573_ sky130_fd_sc_hd__nand2_1
X_12466_ _07700_ _07799_ _00212_ _00206_ VGND VGND VPWR VPWR _02559_ sky130_fd_sc_hd__and4_2
XFILLER_0_81_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14205_ _04397_ _04398_ VGND VGND VPWR VPWR _04399_ sky130_fd_sc_hd__nand2_2
XFILLER_0_124_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11417_ _01151_ _01031_ _09179_ _04078_ VGND VGND VPWR VPWR _01510_ sky130_fd_sc_hd__a22o_1
X_15185_ _05466_ _05467_ _09352_ _07134_ VGND VGND VPWR VPWR _05468_ sky130_fd_sc_hd__and4bb_1
X_12397_ _02489_ _02214_ _02419_ _02420_ VGND VGND VPWR VPWR _02490_ sky130_fd_sc_hd__o22a_1
X_14136_ _04320_ VGND VGND VPWR VPWR _04323_ sky130_fd_sc_hd__inv_2
XFILLER_0_39_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11348_ _01415_ _01439_ _01438_ VGND VGND VPWR VPWR _01441_ sky130_fd_sc_hd__o21ai_2
X_18944_ clknet_4_2_0_clk _00098_ VGND VGND VPWR VPWR cla_inst.in2\[30\] sky130_fd_sc_hd__dfxtp_1
X_14067_ _04245_ _04246_ _04247_ VGND VGND VPWR VPWR _04248_ sky130_fd_sc_hd__mux2_1
X_11279_ _01251_ _01270_ VGND VGND VPWR VPWR _01372_ sky130_fd_sc_hd__nand2_1
X_13018_ _01866_ VGND VGND VPWR VPWR _03111_ sky130_fd_sc_hd__clkbuf_4
X_18875_ clknet_4_14_0_clk net316 VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__dfxtp_1
X_17826_ _03041_ _06443_ _08337_ VGND VGND VPWR VPWR _08338_ sky130_fd_sc_hd__o21a_1
XFILLER_0_55_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17757_ _02200_ _06891_ _06969_ _08150_ VGND VGND VPWR VPWR _08262_ sky130_fd_sc_hd__and4_1
X_14969_ _03008_ _00678_ _05878_ _06471_ VGND VGND VPWR VPWR _05232_ sky130_fd_sc_hd__and4_1
X_16708_ _07117_ _07118_ VGND VGND VPWR VPWR _07119_ sky130_fd_sc_hd__nor2_1
X_17688_ _07038_ _07623_ _08095_ _08186_ VGND VGND VPWR VPWR _08187_ sky130_fd_sc_hd__a31o_1
XFILLER_0_147_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16639_ _07041_ _07043_ VGND VGND VPWR VPWR _07044_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_18_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18309_ _08785_ _08791_ _08861_ VGND VGND VPWR VPWR _08862_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_127_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_710 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_143_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_143_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_142_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_cap130 _02071_ VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__buf_1
XFILLER_0_130_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap141 net325 VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__buf_1
XFILLER_0_111_740 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09944_ _08865_ _08876_ _08887_ _08843_ VGND VGND VPWR VPWR _08897_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_110_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09875_ _07635_ _07657_ VGND VGND VPWR VPWR _08148_ sky130_fd_sc_hd__nand2_2
XTAP_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10650_ _00555_ _00698_ _00741_ _00742_ VGND VGND VPWR VPWR _00743_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_35_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10581_ _00672_ _00673_ VGND VGND VPWR VPWR _00674_ sky130_fd_sc_hd__nor2_1
XFILLER_0_119_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12320_ _02411_ _02412_ VGND VGND VPWR VPWR _02413_ sky130_fd_sc_hd__or2_1
XFILLER_0_23_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12251_ _02336_ _02342_ _02343_ VGND VGND VPWR VPWR _02344_ sky130_fd_sc_hd__a21oi_1
X_11202_ _05224_ _05050_ VGND VGND VPWR VPWR _01295_ sky130_fd_sc_hd__nand2_1
X_12182_ _02270_ _02271_ _02273_ _02274_ VGND VGND VPWR VPWR _02275_ sky130_fd_sc_hd__or4_4
X_11133_ _01137_ _01221_ VGND VGND VPWR VPWR _01226_ sky130_fd_sc_hd__and2_1
X_16990_ _07408_ _07323_ _07425_ VGND VGND VPWR VPWR _07426_ sky130_fd_sc_hd__a21oi_2
X_11064_ _01034_ _01032_ _01033_ VGND VGND VPWR VPWR _01157_ sky130_fd_sc_hd__nand3_1
X_15941_ _06284_ _06286_ VGND VGND VPWR VPWR _06287_ sky130_fd_sc_hd__xnor2_2
X_10015_ _09219_ VGND VGND VPWR VPWR _00108_ sky130_fd_sc_hd__clkbuf_4
X_18660_ net64 _00881_ _09193_ VGND VGND VPWR VPWR _09203_ sky130_fd_sc_hd__mux2_1
X_15872_ _06211_ _06212_ VGND VGND VPWR VPWR _06214_ sky130_fd_sc_hd__nor2_1
X_17611_ _08101_ _08102_ VGND VGND VPWR VPWR _08103_ sky130_fd_sc_hd__nand2_1
X_14823_ _04961_ _04939_ _05071_ _05073_ VGND VGND VPWR VPWR _05074_ sky130_fd_sc_hd__o211ai_2
X_18591_ salida\[15\] _09141_ _09142_ salida\[47\] _09146_ VGND VGND VPWR VPWR _09151_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_99_874 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17542_ _08025_ _08026_ VGND VGND VPWR VPWR _08029_ sky130_fd_sc_hd__or2_1
X_14754_ _04992_ _04993_ _04996_ VGND VGND VPWR VPWR _04998_ sky130_fd_sc_hd__nand3_2
X_11966_ _03728_ VGND VGND VPWR VPWR _02059_ sky130_fd_sc_hd__buf_8
XFILLER_0_58_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10917_ _05638_ _05377_ _05028_ _00992_ VGND VGND VPWR VPWR _01010_ sky130_fd_sc_hd__a22o_1
X_13705_ _03851_ _03687_ VGND VGND VPWR VPWR _03852_ sky130_fd_sc_hd__nand2_1
X_14685_ _04920_ _04921_ _04902_ VGND VGND VPWR VPWR _04923_ sky130_fd_sc_hd__a21o_1
X_17473_ _07833_ _07838_ _07952_ VGND VGND VPWR VPWR _07953_ sky130_fd_sc_hd__o21ai_2
X_11897_ _01988_ _01987_ _01989_ VGND VGND VPWR VPWR _01990_ sky130_fd_sc_hd__or3_4
X_13636_ _00294_ _07102_ cla_inst.in1\[24\] _04351_ VGND VGND VPWR VPWR _03776_ sky130_fd_sc_hd__a22oi_1
X_16424_ _00210_ _06528_ _06530_ _06810_ sel_op\[0\] VGND VGND VPWR VPWR _06811_ sky130_fd_sc_hd__o32a_1
X_10848_ _00925_ _00926_ _00940_ VGND VGND VPWR VPWR _00941_ sky130_fd_sc_hd__nor3b_1
XFILLER_0_66_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13567_ _00115_ _00247_ _03500_ _03499_ VGND VGND VPWR VPWR _03701_ sky130_fd_sc_hd__a31o_1
XFILLER_0_109_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_137_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16355_ _03049_ _06622_ _06735_ _06626_ VGND VGND VPWR VPWR _06736_ sky130_fd_sc_hd__o211a_1
XFILLER_0_41_79 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10779_ cla_inst.in2\[24\] _00174_ _00196_ _00871_ VGND VGND VPWR VPWR _00872_ sky130_fd_sc_hd__nand4_1
XFILLER_0_125_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15306_ _05598_ _05599_ VGND VGND VPWR VPWR _05600_ sky130_fd_sc_hd__nand2_1
X_12518_ _02559_ _02608_ VGND VGND VPWR VPWR _02611_ sky130_fd_sc_hd__or2b_1
XFILLER_0_81_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16286_ _03281_ _03003_ _06520_ VGND VGND VPWR VPWR _06661_ sky130_fd_sc_hd__a21o_1
XFILLER_0_125_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13498_ _05649_ _09256_ _09303_ _06029_ VGND VGND VPWR VPWR _03625_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_54_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18025_ _07108_ _07745_ VGND VGND VPWR VPWR _08554_ sky130_fd_sc_hd__nand2_1
X_15237_ _05428_ _05396_ _05509_ VGND VGND VPWR VPWR _05524_ sky130_fd_sc_hd__a21o_1
X_12449_ _02540_ _02541_ VGND VGND VPWR VPWR _02542_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_124_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15168_ _07635_ VGND VGND VPWR VPWR _05449_ sky130_fd_sc_hd__buf_2
XFILLER_0_10_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14119_ _00644_ _02476_ _03455_ _00513_ VGND VGND VPWR VPWR _04304_ sky130_fd_sc_hd__and4_1
X_15099_ _05265_ _05269_ _05266_ VGND VGND VPWR VPWR _05374_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_5_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18927_ clknet_4_13_0_clk _00081_ VGND VGND VPWR VPWR ApproximateM_inst.lob_16.lob2.genblk1\[13\].genblk1.mux.sel
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09660_ _05192_ _05203_ _05802_ VGND VGND VPWR VPWR _05812_ sky130_fd_sc_hd__a21oi_4
X_18858_ clknet_4_7_0_clk net280 VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__dfxtp_1
X_17809_ _08208_ _08210_ _08206_ VGND VGND VPWR VPWR _08319_ sky130_fd_sc_hd__a21o_1
X_09591_ _05017_ _05050_ VGND VGND VPWR VPWR _05061_ sky130_fd_sc_hd__nand2_1
X_18789_ _09300_ VGND VGND VPWR VPWR _00087_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_900 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_903 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_128_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_122_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_854 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_130_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09927_ _05213_ VGND VGND VPWR VPWR _08713_ sky130_fd_sc_hd__buf_4
X_09858_ cla_inst.in1\[24\] VGND VGND VPWR VPWR _07962_ sky130_fd_sc_hd__clkbuf_4
XTAP_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09789_ _07178_ _07189_ _07199_ VGND VGND VPWR VPWR _07210_ sky130_fd_sc_hd__nand3_4
XTAP_2402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11820_ _01908_ _01912_ VGND VGND VPWR VPWR _01913_ sky130_fd_sc_hd__xor2_1
XANTENNA_103 _09399_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_114 net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_125 _02987_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_136 _05856_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_147 _08762_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_158 _08762_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11751_ _01828_ _01841_ _01842_ net138 VGND VGND VPWR VPWR _01844_ sky130_fd_sc_hd__a211oi_2
XANTENNA_169 _06555_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10702_ _04318_ _04744_ _04755_ VGND VGND VPWR VPWR _00795_ sky130_fd_sc_hd__and3_1
XTAP_1767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14470_ _04686_ _04687_ VGND VGND VPWR VPWR _04688_ sky130_fd_sc_hd__or2b_1
XTAP_1778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_154_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11682_ _01729_ _01774_ VGND VGND VPWR VPWR _01775_ sky130_fd_sc_hd__xnor2_1
XTAP_1789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_730 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13421_ _03058_ _03070_ _03049_ VGND VGND VPWR VPWR _03541_ sky130_fd_sc_hd__mux2_1
X_10633_ _00149_ _00206_ _00172_ _00151_ VGND VGND VPWR VPWR _00726_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_36_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16140_ _00494_ _06470_ _06501_ VGND VGND VPWR VPWR _06502_ sky130_fd_sc_hd__and3_1
X_13352_ _03437_ _03464_ VGND VGND VPWR VPWR _03466_ sky130_fd_sc_hd__xor2_1
XFILLER_0_63_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10564_ _00636_ _00637_ _00655_ _00656_ VGND VGND VPWR VPWR _00657_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_107_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12303_ _02308_ _02310_ _02309_ VGND VGND VPWR VPWR _02396_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_122_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16071_ _00127_ VGND VGND VPWR VPWR _06427_ sky130_fd_sc_hd__clkinv_4
X_13283_ _03382_ _03383_ _03389_ VGND VGND VPWR VPWR _03390_ sky130_fd_sc_hd__nand3_1
X_10495_ _00585_ _00586_ _00418_ _00421_ VGND VGND VPWR VPWR _00588_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_106_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15022_ _05288_ _05289_ VGND VGND VPWR VPWR _05291_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_133_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12234_ _02324_ _02323_ VGND VGND VPWR VPWR _02327_ sky130_fd_sc_hd__and2b_1
XFILLER_0_32_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_570 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12165_ _07853_ _00557_ _02257_ VGND VGND VPWR VPWR _02258_ sky130_fd_sc_hd__and3_2
X_11116_ _01206_ _01208_ VGND VGND VPWR VPWR _01209_ sky130_fd_sc_hd__nand2_1
X_12096_ _02188_ _05017_ _07559_ _07602_ VGND VGND VPWR VPWR _02189_ sky130_fd_sc_hd__and4_1
X_16973_ _07307_ _07309_ VGND VGND VPWR VPWR _07408_ sky130_fd_sc_hd__nand2_1
X_18712_ _09239_ VGND VGND VPWR VPWR _00063_ sky130_fd_sc_hd__clkbuf_1
X_11047_ _00845_ _01139_ _01108_ VGND VGND VPWR VPWR _01140_ sky130_fd_sc_hd__a21o_2
X_15924_ _06260_ _06261_ VGND VGND VPWR VPWR _06269_ sky130_fd_sc_hd__nor2_1
Xinput9 i_wb_addr[16] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__clkbuf_1
X_18643_ _09183_ VGND VGND VPWR VPWR _09190_ sky130_fd_sc_hd__buf_2
X_15855_ _03010_ _03013_ _03154_ _03072_ VGND VGND VPWR VPWR _06195_ sky130_fd_sc_hd__nand4_2
XFILLER_0_87_800 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14806_ _05053_ _05054_ VGND VGND VPWR VPWR _05055_ sky130_fd_sc_hd__xnor2_2
X_18574_ salida\[9\] _09114_ _09118_ salida\[41\] _09128_ VGND VGND VPWR VPWR _09139_
+ sky130_fd_sc_hd__a221o_1
X_15786_ _06053_ _06055_ _06120_ VGND VGND VPWR VPWR _06121_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_87_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12998_ _03085_ _03088_ _03090_ VGND VGND VPWR VPWR _03091_ sky130_fd_sc_hd__mux2_1
X_17525_ _07881_ _07891_ _08008_ VGND VGND VPWR VPWR _08010_ sky130_fd_sc_hd__and3_1
XFILLER_0_59_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14737_ _04977_ _04978_ VGND VGND VPWR VPWR _04979_ sky130_fd_sc_hd__nor2_1
X_11949_ _02028_ _02041_ VGND VGND VPWR VPWR _02042_ sky130_fd_sc_hd__or2_1
XFILLER_0_74_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_143_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17456_ _02127_ _07933_ VGND VGND VPWR VPWR _07934_ sky130_fd_sc_hd__nor2_1
XFILLER_0_129_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14668_ _04781_ _04786_ VGND VGND VPWR VPWR _04904_ sky130_fd_sc_hd__and2b_1
XFILLER_0_74_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16407_ _06336_ _06790_ _06792_ _06543_ _06461_ VGND VGND VPWR VPWR _06793_ sky130_fd_sc_hd__a221o_1
X_13619_ _03454_ _05311_ VGND VGND VPWR VPWR _03757_ sky130_fd_sc_hd__and2_1
XFILLER_0_116_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17387_ _02044_ _07743_ VGND VGND VPWR VPWR _07859_ sky130_fd_sc_hd__nor2_4
X_14599_ _04827_ _04828_ _03538_ VGND VGND VPWR VPWR _04829_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16338_ _03547_ _06717_ _03117_ VGND VGND VPWR VPWR _06718_ sky130_fd_sc_hd__a21o_1
X_16269_ _03547_ _06642_ VGND VGND VPWR VPWR _06643_ sky130_fd_sc_hd__nor2_1
XFILLER_0_140_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18008_ _08533_ _08534_ VGND VGND VPWR VPWR _08535_ sky130_fd_sc_hd__nor2_1
XFILLER_0_11_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_20 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_86 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09712_ _06340_ _06351_ _06362_ VGND VGND VPWR VPWR _06373_ sky130_fd_sc_hd__nand3_4
X_09643_ _05573_ _05595_ _05606_ _05617_ VGND VGND VPWR VPWR _05627_ sky130_fd_sc_hd__and4_1
XFILLER_0_93_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09574_ _04121_ _04657_ _04864_ _04088_ VGND VGND VPWR VPWR _04875_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_117_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10280_ _09152_ _09338_ _00370_ _00371_ VGND VGND VPWR VPWR _00373_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_131_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13970_ _04139_ _04140_ VGND VGND VPWR VPWR _04141_ sky130_fd_sc_hd__nor2_1
X_12921_ _00362_ VGND VGND VPWR VPWR _03014_ sky130_fd_sc_hd__buf_2
XFILLER_0_69_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15640_ _05960_ VGND VGND VPWR VPWR _05962_ sky130_fd_sc_hd__inv_2
XTAP_2210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12852_ _02926_ _02928_ _02943_ _02944_ VGND VGND VPWR VPWR _02945_ sky130_fd_sc_hd__a211o_1
XTAP_2221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11803_ _01741_ _01755_ _01754_ VGND VGND VPWR VPWR _01896_ sky130_fd_sc_hd__a21o_1
XTAP_2254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15571_ _03015_ _03142_ _05886_ _05883_ VGND VGND VPWR VPWR _05887_ sky130_fd_sc_hd__o2bb2a_1
XTAP_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12783_ _02858_ _02860_ VGND VGND VPWR VPWR _02876_ sky130_fd_sc_hd__nor2_1
XTAP_2265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17310_ _07625_ _07626_ _07622_ VGND VGND VPWR VPWR _07775_ sky130_fd_sc_hd__a21bo_1
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14522_ _00678_ _08409_ _00715_ _00679_ VGND VGND VPWR VPWR _04745_ sky130_fd_sc_hd__a22o_1
X_11734_ _01594_ _01599_ VGND VGND VPWR VPWR _01827_ sky130_fd_sc_hd__xnor2_1
XTAP_2298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18290_ _08736_ _08809_ _08749_ VGND VGND VPWR VPWR _08841_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_139_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17241_ _02127_ _06723_ _07675_ _07699_ VGND VGND VPWR VPWR _09390_ sky130_fd_sc_hd__o22a_1
X_14453_ _04649_ _04667_ _04669_ VGND VGND VPWR VPWR _04670_ sky130_fd_sc_hd__nor3_1
X_11665_ _01710_ _01716_ _01717_ _01718_ VGND VGND VPWR VPWR _01758_ sky130_fd_sc_hd__and4_1
Xclkbuf_4_6_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_6_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_154_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13404_ _03370_ _03347_ _03521_ _03522_ VGND VGND VPWR VPWR _03523_ sky130_fd_sc_hd__a211oi_4
X_10616_ _00707_ _00708_ VGND VGND VPWR VPWR _00709_ sky130_fd_sc_hd__xor2_2
X_14384_ _04587_ _04593_ VGND VGND VPWR VPWR _04594_ sky130_fd_sc_hd__xor2_1
XFILLER_0_52_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17172_ _07038_ net146 _07623_ _06527_ VGND VGND VPWR VPWR _07625_ sky130_fd_sc_hd__a22o_1
X_11596_ _01646_ _01653_ _01652_ VGND VGND VPWR VPWR _01689_ sky130_fd_sc_hd__a21o_1
XFILLER_0_3_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13335_ _03439_ _03446_ VGND VGND VPWR VPWR _03447_ sky130_fd_sc_hd__or2_1
XFILLER_0_51_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16123_ _06483_ VGND VGND VPWR VPWR _06484_ sky130_fd_sc_hd__clkbuf_4
X_10547_ _06029_ _06051_ _07384_ _07015_ VGND VGND VPWR VPWR _00640_ sky130_fd_sc_hd__and4_1
XFILLER_0_134_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13266_ _00661_ net327 _03293_ _03294_ VGND VGND VPWR VPWR _03371_ sky130_fd_sc_hd__o211a_1
X_16054_ _03016_ _06408_ VGND VGND VPWR VPWR _06409_ sky130_fd_sc_hd__nor2_1
X_10478_ _00562_ _00570_ VGND VGND VPWR VPWR _00571_ sky130_fd_sc_hd__xnor2_1
X_15005_ _05270_ _05264_ VGND VGND VPWR VPWR _05272_ sky130_fd_sc_hd__or2b_1
X_12217_ _02306_ _02307_ _02295_ _02299_ VGND VGND VPWR VPWR _02310_ sky130_fd_sc_hd__a211oi_1
X_13197_ _00191_ _00398_ _00247_ _00189_ VGND VGND VPWR VPWR _03298_ sky130_fd_sc_hd__a22oi_1
X_12148_ _07069_ _00210_ _03607_ _07036_ VGND VGND VPWR VPWR _02241_ sky130_fd_sc_hd__a22o_1
XFILLER_0_138_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12079_ _01810_ _01903_ _02171_ VGND VGND VPWR VPWR _02172_ sky130_fd_sc_hd__a21o_1
X_16956_ _04034_ _03324_ _06814_ _07386_ VGND VGND VPWR VPWR _07389_ sky130_fd_sc_hd__a211oi_2
X_15907_ _06249_ _06250_ _06200_ _03072_ VGND VGND VPWR VPWR _06251_ sky130_fd_sc_hd__o211ai_1
X_16887_ _07313_ VGND VGND VPWR VPWR _07314_ sky130_fd_sc_hd__buf_4
XFILLER_0_78_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18626_ salida\[30\] _09113_ _09117_ salida\[62\] _09163_ VGND VGND VPWR VPWR _09175_
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_154_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15838_ _06175_ _06176_ VGND VGND VPWR VPWR _06177_ sky130_fd_sc_hd__or2_1
XFILLER_0_63_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18557_ _09127_ VGND VGND VPWR VPWR _09128_ sky130_fd_sc_hd__buf_2
X_15769_ _01417_ _04125_ VGND VGND VPWR VPWR _06102_ sky130_fd_sc_hd__nand2_1
XFILLER_0_63_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17508_ _07975_ _07976_ _07990_ VGND VGND VPWR VPWR _07991_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_86_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18488_ _09052_ _09053_ _09054_ VGND VGND VPWR VPWR _09055_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_7_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_14 _01108_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17439_ _03108_ _06440_ VGND VGND VPWR VPWR _07916_ sky130_fd_sc_hd__nor2_1
XANTENNA_25 _01115_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_36 _01503_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_47 _02969_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_58 _04241_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_284 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_69 _05625_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_654 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput110 net110 VGND VGND VPWR VPWR o_wb_data[5] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_112_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09626_ _05268_ _05431_ VGND VGND VPWR VPWR _05442_ sky130_fd_sc_hd__xnor2_2
X_09557_ ApproximateM_inst.lob_16.lob2.genblk1\[11\].genblk1.mux.sel VGND VGND VPWR
+ VPWR _04690_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_77_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09488_ _03870_ _03925_ VGND VGND VPWR VPWR _03935_ sky130_fd_sc_hd__nor2_1
XFILLER_0_38_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_108_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11450_ _04690_ _00211_ _01541_ _01542_ VGND VGND VPWR VPWR _01543_ sky130_fd_sc_hd__nand4_2
XFILLER_0_92_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10401_ _06993_ VGND VGND VPWR VPWR _00494_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_150_215 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11381_ _00163_ _00881_ VGND VGND VPWR VPWR _01474_ sky130_fd_sc_hd__nand2_2
XFILLER_0_6_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13120_ _04088_ _04121_ _05333_ VGND VGND VPWR VPWR _03215_ sky130_fd_sc_hd__and3_1
XFILLER_0_104_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10332_ net338 _00377_ _09346_ _00274_ VGND VGND VPWR VPWR _00425_ sky130_fd_sc_hd__o211a_1
XFILLER_0_61_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13051_ _03142_ VGND VGND VPWR VPWR _03143_ sky130_fd_sc_hd__clkbuf_4
X_10263_ _00353_ _00354_ _09271_ VGND VGND VPWR VPWR _00356_ sky130_fd_sc_hd__o21ai_1
X_12002_ _05301_ _00180_ _00130_ _05279_ VGND VGND VPWR VPWR _02095_ sky130_fd_sc_hd__a22o_1
X_10194_ _00278_ _00279_ _00280_ VGND VGND VPWR VPWR _00287_ sky130_fd_sc_hd__a21o_1
XFILLER_0_100_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16810_ _07193_ _07228_ VGND VGND VPWR VPWR _07230_ sky130_fd_sc_hd__nand2_1
X_17790_ _08173_ _08178_ _08297_ VGND VGND VPWR VPWR _08298_ sky130_fd_sc_hd__a21oi_1
X_16741_ _07059_ _07061_ VGND VGND VPWR VPWR _07155_ sky130_fd_sc_hd__and2b_1
X_13953_ _03949_ _04091_ _04120_ _04122_ VGND VGND VPWR VPWR _04123_ sky130_fd_sc_hd__o211a_4
X_12904_ _02996_ VGND VGND VPWR VPWR _02997_ sky130_fd_sc_hd__buf_2
X_16672_ _06426_ _06435_ _07076_ _07079_ VGND VGND VPWR VPWR _07081_ sky130_fd_sc_hd__o31a_1
X_13884_ _04006_ _03877_ _04046_ _04047_ VGND VGND VPWR VPWR _04048_ sky130_fd_sc_hd__a211oi_2
X_18411_ _08872_ _08921_ VGND VGND VPWR VPWR _08972_ sky130_fd_sc_hd__or2b_1
X_15623_ _05866_ _05870_ _05944_ VGND VGND VPWR VPWR _05945_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_69_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12835_ _02901_ _02922_ _02926_ _02927_ VGND VGND VPWR VPWR _02928_ sky130_fd_sc_hd__o211ai_4
XTAP_2051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18342_ _06374_ _00558_ _04995_ VGND VGND VPWR VPWR _08898_ sky130_fd_sc_hd__a21o_1
X_15554_ _05752_ _05868_ _05869_ VGND VGND VPWR VPWR _05870_ sky130_fd_sc_hd__and3_1
XTAP_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12766_ _02856_ _02857_ _01790_ _02855_ VGND VGND VPWR VPWR _02859_ sky130_fd_sc_hd__a211oi_1
XTAP_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14505_ _08615_ _03456_ _04589_ _04588_ _04725_ VGND VGND VPWR VPWR _04726_ sky130_fd_sc_hd__a32o_2
XTAP_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18273_ _07084_ _08821_ _08823_ VGND VGND VPWR VPWR _08824_ sky130_fd_sc_hd__or3_1
XFILLER_0_83_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11717_ _01808_ _01809_ VGND VGND VPWR VPWR _01810_ sky130_fd_sc_hd__nor2_4
X_15485_ _05612_ _05708_ _05709_ _05794_ VGND VGND VPWR VPWR _05795_ sky130_fd_sc_hd__o211a_1
X_12697_ _02756_ _02757_ _02758_ _02754_ VGND VGND VPWR VPWR _02790_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_83_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17224_ _07566_ _07567_ _07565_ VGND VGND VPWR VPWR _07682_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_37_582 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14436_ _04516_ _04521_ VGND VGND VPWR VPWR _04651_ sky130_fd_sc_hd__and2b_1
X_11648_ _01642_ net125 _01739_ _01740_ VGND VGND VPWR VPWR _01741_ sky130_fd_sc_hd__o211ai_4
Xinput12 i_wb_addr[19] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput23 i_wb_addr[29] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__clkbuf_1
Xinput34 i_wb_cyc VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__buf_2
XFILLER_0_126_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput45 i_wb_data[19] VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__clkbuf_2
X_17155_ _06891_ _07109_ _07499_ _07605_ VGND VGND VPWR VPWR _07606_ sky130_fd_sc_hd__a31o_1
XFILLER_0_142_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14367_ _03793_ _07374_ _07406_ _03859_ VGND VGND VPWR VPWR _04575_ sky130_fd_sc_hd__a22oi_1
X_11579_ _07799_ _05845_ VGND VGND VPWR VPWR _01672_ sky130_fd_sc_hd__and2_2
XFILLER_0_24_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput56 i_wb_data[29] VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__buf_1
Xinput67 i_wb_stb VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__clkbuf_4
X_16106_ _03121_ _06454_ VGND VGND VPWR VPWR _06465_ sky130_fd_sc_hd__nor2_1
X_13318_ _03254_ _03256_ _03426_ _03427_ VGND VGND VPWR VPWR _03428_ sky130_fd_sc_hd__a211oi_4
X_14298_ _04339_ _04343_ _04341_ VGND VGND VPWR VPWR _04500_ sky130_fd_sc_hd__o21ba_1
X_17086_ _07508_ _07509_ _07530_ VGND VGND VPWR VPWR _07531_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_110_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16037_ _00592_ _04336_ VGND VGND VPWR VPWR _06390_ sky130_fd_sc_hd__or2_2
XFILLER_0_149_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13249_ _03351_ _03352_ VGND VGND VPWR VPWR _03353_ sky130_fd_sc_hd__xor2_1
XFILLER_0_58_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17988_ _08429_ _08430_ _08427_ VGND VGND VPWR VPWR _08514_ sky130_fd_sc_hd__a21bo_1
X_16939_ _03079_ _06698_ VGND VGND VPWR VPWR _07371_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18609_ net257 _09157_ _09164_ _09162_ VGND VGND VPWR VPWR _00025_ sky130_fd_sc_hd__o211a_1
XFILLER_0_149_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_114_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_418 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_117_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10950_ _01041_ _01042_ VGND VGND VPWR VPWR _01043_ sky130_fd_sc_hd__xnor2_2
X_09609_ _05246_ VGND VGND VPWR VPWR _05257_ sky130_fd_sc_hd__buf_4
X_10881_ _00968_ _00973_ VGND VGND VPWR VPWR _00974_ sky130_fd_sc_hd__xor2_1
XFILLER_0_97_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12620_ _07091_ _07363_ _07570_ _07602_ VGND VGND VPWR VPWR _02713_ sky130_fd_sc_hd__and4_1
X_12551_ _02635_ _02641_ _02642_ VGND VGND VPWR VPWR _02644_ sky130_fd_sc_hd__nand3_1
XFILLER_0_108_223 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_474 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11502_ _06711_ _00715_ VGND VGND VPWR VPWR _01595_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15270_ _01317_ _05558_ _05559_ VGND VGND VPWR VPWR _05560_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_108_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12482_ _02504_ _02571_ _02573_ VGND VGND VPWR VPWR _02575_ sky130_fd_sc_hd__nand3_1
XFILLER_0_62_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11433_ _01514_ _01524_ VGND VGND VPWR VPWR _01526_ sky130_fd_sc_hd__xor2_1
X_14221_ _03078_ VGND VGND VPWR VPWR _04415_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14152_ _00190_ _00192_ _06482_ _04591_ VGND VGND VPWR VPWR _04341_ sky130_fd_sc_hd__and4_1
X_11364_ _00123_ _00848_ _00849_ VGND VGND VPWR VPWR _01457_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_61_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10315_ _00404_ _00407_ VGND VGND VPWR VPWR _00408_ sky130_fd_sc_hd__xnor2_1
X_13103_ _03036_ _03123_ VGND VGND VPWR VPWR _03197_ sky130_fd_sc_hd__nor2_2
XFILLER_0_132_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14083_ _04261_ _04264_ _03539_ VGND VGND VPWR VPWR _04265_ sky130_fd_sc_hd__mux2_1
X_18960_ clknet_4_6_0_clk _09390_ VGND VGND VPWR VPWR salida\[13\] sky130_fd_sc_hd__dfxtp_1
X_11295_ _01385_ _01284_ _01386_ VGND VGND VPWR VPWR _01388_ sky130_fd_sc_hd__nand3_2
XFILLER_0_131_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17911_ _08330_ _08331_ _08329_ VGND VGND VPWR VPWR _08430_ sky130_fd_sc_hd__o21bai_2
X_13034_ _03028_ _02779_ VGND VGND VPWR VPWR _03126_ sky130_fd_sc_hd__nor2_1
X_10246_ _07744_ VGND VGND VPWR VPWR _00339_ sky130_fd_sc_hd__buf_4
XFILLER_0_28_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18891_ clknet_4_11_0_clk _00045_ VGND VGND VPWR VPWR ApproximateM_inst.lob_16.lob1.genblk1\[9\].genblk1.mux.sel
+ sky130_fd_sc_hd__dfxtp_2
X_17842_ net146 net145 VGND VGND VPWR VPWR _08355_ sky130_fd_sc_hd__nand2_1
X_10177_ _00161_ _00231_ _00268_ _00269_ VGND VGND VPWR VPWR _00270_ sky130_fd_sc_hd__a211o_2
X_17773_ _08162_ _08163_ _08161_ VGND VGND VPWR VPWR _08280_ sky130_fd_sc_hd__o21ai_2
X_14985_ _00148_ _00149_ _06062_ _05257_ VGND VGND VPWR VPWR _05250_ sky130_fd_sc_hd__and4_1
X_16724_ _07133_ _07136_ VGND VGND VPWR VPWR _07137_ sky130_fd_sc_hd__xor2_1
X_13936_ _04001_ _07123_ VGND VGND VPWR VPWR _04104_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16655_ _07059_ _07061_ VGND VGND VPWR VPWR _07062_ sky130_fd_sc_hd__xnor2_1
X_13867_ _00107_ _04012_ _03867_ _03866_ VGND VGND VPWR VPWR _04029_ sky130_fd_sc_hd__a31o_1
X_15606_ _05924_ _05925_ VGND VGND VPWR VPWR _05926_ sky130_fd_sc_hd__nor2_1
XFILLER_0_29_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12818_ _02896_ _02897_ _02909_ _02910_ VGND VGND VPWR VPWR _02911_ sky130_fd_sc_hd__a211o_1
X_16586_ _03206_ _06986_ VGND VGND VPWR VPWR _06987_ sky130_fd_sc_hd__nor2_1
X_13798_ _00294_ _07004_ _07102_ _04504_ VGND VGND VPWR VPWR _03953_ sky130_fd_sc_hd__a22oi_1
X_18325_ _03201_ _08878_ _08879_ VGND VGND VPWR VPWR _08880_ sky130_fd_sc_hd__and3_2
X_15537_ _05849_ _00119_ _05449_ _05850_ VGND VGND VPWR VPWR _05851_ sky130_fd_sc_hd__and4b_1
XTAP_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12749_ _02751_ _02836_ _02839_ _02841_ VGND VGND VPWR VPWR _02842_ sky130_fd_sc_hd__o31a_1
XFILLER_0_151_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18256_ _08732_ _08731_ VGND VGND VPWR VPWR _08805_ sky130_fd_sc_hd__or2b_1
X_15468_ _05716_ _05695_ _05774_ _05775_ VGND VGND VPWR VPWR _05776_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_60_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17207_ _07661_ _07662_ VGND VGND VPWR VPWR _07663_ sky130_fd_sc_hd__xnor2_1
X_14419_ _00702_ _05486_ _05878_ _00195_ VGND VGND VPWR VPWR _04632_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_53_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18187_ _08636_ _08644_ _08646_ VGND VGND VPWR VPWR _08730_ sky130_fd_sc_hd__a21oi_1
X_15399_ _05499_ _05602_ VGND VGND VPWR VPWR _05701_ sky130_fd_sc_hd__or2_1
XFILLER_0_130_719 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17138_ _07552_ _07553_ VGND VGND VPWR VPWR _07587_ sky130_fd_sc_hd__and2_1
XFILLER_0_40_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_122_270 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09960_ _06993_ _09059_ _07428_ _07417_ VGND VGND VPWR VPWR _09070_ sky130_fd_sc_hd__a31o_1
X_17069_ _07124_ _07126_ _07511_ _06561_ VGND VGND VPWR VPWR _07512_ sky130_fd_sc_hd__o22a_1
XFILLER_0_110_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09891_ _06373_ _06504_ _06515_ VGND VGND VPWR VPWR _08322_ sky130_fd_sc_hd__nand3_2
XFILLER_0_0_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_149_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_839 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_118_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10100_ _00147_ VGND VGND VPWR VPWR _00193_ sky130_fd_sc_hd__buf_4
X_11080_ _00294_ _00210_ _00205_ _04504_ VGND VGND VPWR VPWR _01173_ sky130_fd_sc_hd__a22o_1
X_10031_ _00110_ _00114_ VGND VGND VPWR VPWR _00124_ sky130_fd_sc_hd__or2_1
XFILLER_0_98_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14770_ _05012_ _05013_ _04867_ _04968_ VGND VGND VPWR VPWR _05015_ sky130_fd_sc_hd__o211ai_2
X_11982_ _02053_ _02074_ VGND VGND VPWR VPWR _02075_ sky130_fd_sc_hd__nand2_1
X_13721_ _03867_ _03868_ VGND VGND VPWR VPWR _03869_ sky130_fd_sc_hd__xnor2_1
X_10933_ _01024_ _01025_ VGND VGND VPWR VPWR _01026_ sky130_fd_sc_hd__and2b_1
XFILLER_0_86_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16440_ _06824_ _06827_ VGND VGND VPWR VPWR _06828_ sky130_fd_sc_hd__xnor2_1
X_13652_ _03791_ _03792_ VGND VGND VPWR VPWR _03794_ sky130_fd_sc_hd__nor2_1
X_10864_ ApproximateM_inst.lob_16.lob2.genblk2.mux_final.sel ApproximateM_inst.lob_16.lob1.genblk1\[9\].genblk1.mux.sel
+ ApproximateM_inst.lob_16.lob1.genblk1\[8\].genblk1.mux.sel cla_inst.in2\[16\] VGND
+ VGND VPWR VPWR _00957_ sky130_fd_sc_hd__a22o_1
XFILLER_0_128_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12603_ _02672_ _02673_ _02692_ VGND VGND VPWR VPWR _02696_ sky130_fd_sc_hd__a21oi_1
XPHY_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16371_ _03324_ _06752_ net343 VGND VGND VPWR VPWR _06753_ sky130_fd_sc_hd__o21ai_2
XPHY_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13583_ _03715_ _03716_ _03676_ _03677_ VGND VGND VPWR VPWR _03719_ sky130_fd_sc_hd__a211oi_2
X_10795_ _00860_ _00865_ _00867_ _00887_ VGND VGND VPWR VPWR _00888_ sky130_fd_sc_hd__a22o_1
XFILLER_0_54_614 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18110_ _08635_ _08645_ VGND VGND VPWR VPWR _08646_ sky130_fd_sc_hd__and2_1
X_15322_ _05416_ _05615_ _05616_ VGND VGND VPWR VPWR _05618_ sky130_fd_sc_hd__a21oi_1
XPHY_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12534_ _02618_ _02625_ _02626_ VGND VGND VPWR VPWR _02627_ sky130_fd_sc_hd__o21ai_1
XPHY_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18041_ _08490_ _08570_ VGND VGND VPWR VPWR _08571_ sky130_fd_sc_hd__xnor2_1
X_15253_ _05539_ VGND VGND VPWR VPWR _05542_ sky130_fd_sc_hd__inv_2
X_12465_ _02544_ _02557_ VGND VGND VPWR VPWR _02558_ sky130_fd_sc_hd__xnor2_1
X_14204_ _04393_ _04394_ _04396_ VGND VGND VPWR VPWR _04398_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_62_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11416_ _04078_ _01151_ _00871_ VGND VGND VPWR VPWR _01509_ sky130_fd_sc_hd__and3_1
X_15184_ _00148_ _00149_ _00308_ _05964_ VGND VGND VPWR VPWR _05467_ sky130_fd_sc_hd__and4_1
XFILLER_0_22_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12396_ ApproximateM_inst.lob_16.lob2.genblk1\[2\].genblk1.mux.sel VGND VGND VPWR
+ VPWR _02489_ sky130_fd_sc_hd__inv_4
XFILLER_0_111_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14135_ _04320_ _04012_ _00362_ _04321_ VGND VGND VPWR VPWR _04322_ sky130_fd_sc_hd__and4b_1
XFILLER_0_10_717 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11347_ _01415_ _01438_ _01439_ VGND VGND VPWR VPWR _01440_ sky130_fd_sc_hd__or3_4
XFILLER_0_39_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18943_ clknet_4_2_0_clk _00097_ VGND VGND VPWR VPWR cla_inst.in2\[29\] sky130_fd_sc_hd__dfxtp_2
X_11278_ _01252_ _01269_ VGND VGND VPWR VPWR _01371_ sky130_fd_sc_hd__or2b_1
X_14066_ _03079_ VGND VGND VPWR VPWR _04247_ sky130_fd_sc_hd__clkbuf_4
X_10229_ _07025_ VGND VGND VPWR VPWR _00322_ sky130_fd_sc_hd__buf_4
X_13017_ _03040_ _03109_ VGND VGND VPWR VPWR _03110_ sky130_fd_sc_hd__nand2_1
X_18874_ clknet_4_15_0_clk net249 VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__dfxtp_1
X_17825_ _03041_ _06443_ _06424_ VGND VGND VPWR VPWR _08337_ sky130_fd_sc_hd__a21oi_1
X_17756_ _06961_ _07706_ _08260_ _07018_ VGND VGND VPWR VPWR _08261_ sky130_fd_sc_hd__o22a_1
X_14968_ _05230_ VGND VGND VPWR VPWR _05231_ sky130_fd_sc_hd__inv_2
X_16707_ _06766_ _06875_ _07114_ _07116_ VGND VGND VPWR VPWR _07118_ sky130_fd_sc_hd__o22a_1
X_13919_ _03538_ _03124_ _04076_ _04085_ _03199_ VGND VGND VPWR VPWR _04086_ sky130_fd_sc_hd__a32o_1
X_17687_ _08094_ _08092_ VGND VGND VPWR VPWR _08186_ sky130_fd_sc_hd__and2b_1
X_14899_ _05018_ _05027_ _05025_ VGND VGND VPWR VPWR _05156_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_9_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16638_ _06579_ _07042_ VGND VGND VPWR VPWR _07043_ sky130_fd_sc_hd__nor2_1
XFILLER_0_119_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16569_ _06878_ _06879_ _00194_ VGND VGND VPWR VPWR _06968_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_85_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18308_ _08859_ _08860_ VGND VGND VPWR VPWR _08861_ sky130_fd_sc_hd__or2_1
XFILLER_0_127_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18239_ _08784_ _08785_ VGND VGND VPWR VPWR _08786_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_cap120 net319 VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__buf_1
XFILLER_0_20_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09943_ _08832_ VGND VGND VPWR VPWR _08887_ sky130_fd_sc_hd__inv_2
XFILLER_0_111_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_96_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09874_ _07319_ _07940_ _08115_ VGND VGND VPWR VPWR _08137_ sky130_fd_sc_hd__a21o_1
XTAP_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_536 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_107 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10580_ _00670_ _00671_ _00667_ VGND VGND VPWR VPWR _00673_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_91_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12250_ _02218_ _02220_ VGND VGND VPWR VPWR _02343_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_50_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11201_ _00974_ _00975_ VGND VGND VPWR VPWR _01294_ sky130_fd_sc_hd__nand2_1
XFILLER_0_133_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12181_ _02128_ _02258_ VGND VGND VPWR VPWR _02274_ sky130_fd_sc_hd__and2_1
X_11132_ _07853_ _01223_ _01224_ VGND VGND VPWR VPWR _01225_ sky130_fd_sc_hd__a21oi_4
X_11063_ _01154_ _01155_ VGND VGND VPWR VPWR _01156_ sky130_fd_sc_hd__xnor2_1
X_15940_ _06258_ _06285_ VGND VGND VPWR VPWR _06286_ sky130_fd_sc_hd__nand2_1
X_10014_ _00106_ VGND VGND VPWR VPWR _00107_ sky130_fd_sc_hd__clkbuf_4
X_15871_ _06209_ _06210_ VGND VGND VPWR VPWR _06212_ sky130_fd_sc_hd__and2_1
X_17610_ _08099_ _08100_ VGND VGND VPWR VPWR _08102_ sky130_fd_sc_hd__nand2_1
X_14822_ _05069_ _05070_ _04896_ _04963_ VGND VGND VPWR VPWR _05073_ sky130_fd_sc_hd__a211o_1
X_18590_ net285 _09140_ _09150_ _09144_ VGND VGND VPWR VPWR _00018_ sky130_fd_sc_hd__o211a_1
XFILLER_0_25_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_26 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17541_ _08025_ _08026_ VGND VGND VPWR VPWR _08027_ sky130_fd_sc_hd__nand2_1
X_14753_ _04992_ _04993_ _04996_ VGND VGND VPWR VPWR _04997_ sky130_fd_sc_hd__a21o_1
XFILLER_0_98_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11965_ _02007_ _02057_ VGND VGND VPWR VPWR _02058_ sky130_fd_sc_hd__and2_1
XFILLER_0_99_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13704_ _03682_ _03683_ VGND VGND VPWR VPWR _03851_ sky130_fd_sc_hd__or2b_1
X_10916_ _00992_ _05638_ net235 VGND VGND VPWR VPWR _01009_ sky130_fd_sc_hd__and3_1
X_17472_ _07707_ _07832_ VGND VGND VPWR VPWR _07952_ sky130_fd_sc_hd__or2_1
X_14684_ _04902_ _04920_ _04921_ VGND VGND VPWR VPWR _04922_ sky130_fd_sc_hd__nand3_1
X_11896_ _01986_ _01980_ _01984_ VGND VGND VPWR VPWR _01989_ sky130_fd_sc_hd__and3_1
X_16423_ ApproximateM_inst.lob_16.lob1.genblk2.mux_final.sel ApproximateM_inst.lob_16.lob1.genblk1\[14\].genblk1.mux.sel
+ ApproximateM_inst.lob_16.lob1.genblk1\[13\].genblk1.mux.sel ApproximateM_inst.lob_16.lob1.genblk1\[12\].genblk1.mux.sel
+ _03184_ VGND VGND VPWR VPWR _06810_ sky130_fd_sc_hd__o41a_1
X_13635_ _03600_ _03601_ _03599_ VGND VGND VPWR VPWR _03775_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_132_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10847_ _00931_ _00938_ _00939_ VGND VGND VPWR VPWR _00940_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_67_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16354_ _01677_ _06637_ VGND VGND VPWR VPWR _06735_ sky130_fd_sc_hd__or2_1
X_13566_ _03495_ _03503_ _03699_ VGND VGND VPWR VPWR _03700_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_66_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10778_ ApproximateM_inst.lob_16.lob1.genblk1\[2\].genblk1.mux.sel VGND VGND VPWR
+ VPWR _00871_ sky130_fd_sc_hd__buf_4
XFILLER_0_109_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15305_ _05596_ _05597_ _05552_ VGND VGND VPWR VPWR _05599_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_82_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12517_ _00120_ _00213_ _00207_ _07711_ VGND VGND VPWR VPWR _02610_ sky130_fd_sc_hd__a22o_1
XFILLER_0_124_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16285_ _02728_ net344 VGND VGND VPWR VPWR _06660_ sky130_fd_sc_hd__nor2_1
X_13497_ _03395_ _03403_ _03402_ VGND VGND VPWR VPWR _03624_ sky130_fd_sc_hd__a21o_1
XFILLER_0_125_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18024_ _08551_ _08552_ VGND VGND VPWR VPWR _08553_ sky130_fd_sc_hd__nand2_2
X_15236_ _03082_ _05307_ _05425_ _03039_ _05523_ VGND VGND VPWR VPWR _09362_ sky130_fd_sc_hd__o221ai_2
XFILLER_0_124_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12448_ _02501_ _02507_ VGND VGND VPWR VPWR _02541_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_140_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15167_ _03014_ _01223_ _05447_ VGND VGND VPWR VPWR _05448_ sky130_fd_sc_hd__and3_1
XFILLER_0_10_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12379_ _02458_ _02459_ _02452_ VGND VGND VPWR VPWR _02472_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_50_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14118_ _02476_ _03456_ _00665_ _00644_ VGND VGND VPWR VPWR _04303_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_10_558 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15098_ _05371_ _05372_ VGND VGND VPWR VPWR _05373_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_120_571 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14049_ _04225_ _04226_ _04227_ VGND VGND VPWR VPWR _04228_ sky130_fd_sc_hd__and3_2
X_18926_ clknet_4_13_0_clk _00080_ VGND VGND VPWR VPWR ApproximateM_inst.lob_16.lob2.genblk1\[12\].genblk1.mux.sel
+ sky130_fd_sc_hd__dfxtp_2
X_18857_ clknet_4_4_0_clk net266 VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__dfxtp_1
X_17808_ _08316_ _08317_ VGND VGND VPWR VPWR _08318_ sky130_fd_sc_hd__xor2_1
X_09590_ _05039_ VGND VGND VPWR VPWR _05050_ sky130_fd_sc_hd__clkbuf_8
X_18788_ _09298_ _09299_ VGND VGND VPWR VPWR _09300_ sky130_fd_sc_hd__and2_1
XFILLER_0_77_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17739_ _02973_ _06645_ VGND VGND VPWR VPWR _08243_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_122_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09926_ _06493_ _06450_ VGND VGND VPWR VPWR _08702_ sky130_fd_sc_hd__or2b_1
XTAP_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09857_ _07036_ _07069_ _05693_ cla_inst.in1\[22\] VGND VGND VPWR VPWR _07951_ sky130_fd_sc_hd__nand4_2
XTAP_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09788_ _06993_ _07025_ _07145_ _07167_ VGND VGND VPWR VPWR _07199_ sky130_fd_sc_hd__a22o_1
XTAP_2403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_104 _09402_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_115 net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_126 _03201_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_137 _05856_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_148 _08762_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11750_ _01670_ _01676_ _01679_ _01680_ VGND VGND VPWR VPWR _01843_ sky130_fd_sc_hd__nor4_1
XTAP_2469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_159 _08762_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_366 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10701_ _00779_ _00792_ _00793_ VGND VGND VPWR VPWR _00794_ sky130_fd_sc_hd__nand3_4
XTAP_1757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11681_ _01507_ _01773_ VGND VGND VPWR VPWR _01774_ sky130_fd_sc_hd__or2b_1
XTAP_1779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13420_ _03046_ _03054_ _03049_ VGND VGND VPWR VPWR _03540_ sky130_fd_sc_hd__mux2_1
X_10632_ _07537_ _00147_ _00520_ _00359_ _00132_ VGND VGND VPWR VPWR _00725_ sky130_fd_sc_hd__a32o_1
XFILLER_0_64_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10563_ _00653_ _00654_ _00638_ VGND VGND VPWR VPWR _00656_ sky130_fd_sc_hd__a21bo_1
X_13351_ _03438_ _03463_ VGND VGND VPWR VPWR _03464_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_64_786 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_146_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_594 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_107_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12302_ _02393_ _02392_ _02394_ VGND VGND VPWR VPWR _02395_ sky130_fd_sc_hd__nor3_1
X_16070_ _06425_ VGND VGND VPWR VPWR _06426_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_106_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13282_ _03386_ _03387_ VGND VGND VPWR VPWR _03389_ sky130_fd_sc_hd__xor2_2
X_10494_ _00418_ _00421_ _00585_ _00586_ VGND VGND VPWR VPWR _00587_ sky130_fd_sc_hd__a211o_1
XFILLER_0_122_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15021_ _05139_ _05183_ _05136_ VGND VGND VPWR VPWR _05289_ sky130_fd_sc_hd__a21oi_2
X_12233_ _02321_ _02325_ VGND VGND VPWR VPWR _02326_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_122_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12164_ _00515_ _02127_ VGND VGND VPWR VPWR _02257_ sky130_fd_sc_hd__nor2_2
XFILLER_0_20_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11115_ _06982_ _00443_ _01206_ _01207_ VGND VGND VPWR VPWR _01208_ sky130_fd_sc_hd__nand4_2
X_12095_ _04373_ VGND VGND VPWR VPWR _02188_ sky130_fd_sc_hd__clkbuf_8
X_16972_ _07385_ _07405_ VGND VGND VPWR VPWR _07407_ sky130_fd_sc_hd__xnor2_1
X_11046_ _05986_ VGND VGND VPWR VPWR _01139_ sky130_fd_sc_hd__clkbuf_4
X_18711_ _09209_ _09238_ VGND VGND VPWR VPWR _09239_ sky130_fd_sc_hd__and2_1
X_15923_ _02969_ _06264_ _06265_ _06268_ VGND VGND VPWR VPWR _09374_ sky130_fd_sc_hd__o31ai_4
X_18642_ _09183_ VGND VGND VPWR VPWR _09189_ sky130_fd_sc_hd__buf_2
X_15854_ _03012_ _03154_ _03072_ _03010_ VGND VGND VPWR VPWR _06194_ sky130_fd_sc_hd__a22o_1
X_14805_ _01873_ _03055_ VGND VGND VPWR VPWR _05054_ sky130_fd_sc_hd__nand2_1
XFILLER_0_59_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18573_ net271 _09098_ _09138_ _09126_ VGND VGND VPWR VPWR _00012_ sky130_fd_sc_hd__o211a_1
X_15785_ _06118_ _06119_ VGND VGND VPWR VPWR _06120_ sky130_fd_sc_hd__and2_1
X_12997_ _03089_ VGND VGND VPWR VPWR _03090_ sky130_fd_sc_hd__clkbuf_4
X_17524_ _07881_ _07891_ _08008_ VGND VGND VPWR VPWR _08009_ sky130_fd_sc_hd__a21oi_2
X_14736_ _04099_ _04034_ _00502_ _09248_ VGND VGND VPWR VPWR _04978_ sky130_fd_sc_hd__and4_1
XFILLER_0_86_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11948_ _02031_ _02039_ _02040_ VGND VGND VPWR VPWR _02041_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_129_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17455_ _04034_ _06889_ VGND VGND VPWR VPWR _07933_ sky130_fd_sc_hd__nand2_1
X_14667_ _04619_ _04789_ VGND VGND VPWR VPWR _04903_ sky130_fd_sc_hd__or2_1
XFILLER_0_86_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11879_ _01869_ _01970_ _01938_ _01969_ VGND VGND VPWR VPWR _01972_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_117_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16406_ _06431_ _06791_ VGND VGND VPWR VPWR _06792_ sky130_fd_sc_hd__nor2_1
X_13618_ _03531_ _03509_ _06613_ net223 VGND VGND VPWR VPWR _03756_ sky130_fd_sc_hd__nand4_2
XFILLER_0_6_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17386_ _07856_ _07857_ VGND VGND VPWR VPWR _07858_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14598_ _03916_ _03546_ VGND VGND VPWR VPWR _04828_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16337_ _03164_ _06470_ _06713_ _06716_ VGND VGND VPWR VPWR _06717_ sky130_fd_sc_hd__a31o_1
X_13549_ _00169_ _08409_ VGND VGND VPWR VPWR _03681_ sky130_fd_sc_hd__nand2_1
XFILLER_0_109_192 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16268_ _06639_ _06641_ _03061_ VGND VGND VPWR VPWR _06642_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18007_ _07665_ _07596_ _08453_ VGND VGND VPWR VPWR _08534_ sky130_fd_sc_hd__and3_1
X_15219_ _05503_ _05504_ VGND VGND VPWR VPWR _05505_ sky130_fd_sc_hd__and2_1
XFILLER_0_2_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16199_ _03410_ _03673_ _06529_ _06565_ VGND VGND VPWR VPWR _06566_ sky130_fd_sc_hd__or4_4
XFILLER_0_77_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09711_ _04919_ _04930_ _04842_ VGND VGND VPWR VPWR _06362_ sky130_fd_sc_hd__a21bo_1
X_18909_ clknet_4_10_0_clk _00063_ VGND VGND VPWR VPWR cla_inst.in1\[27\] sky130_fd_sc_hd__dfxtp_4
X_09642_ cla_inst.in1\[21\] VGND VGND VPWR VPWR _05617_ sky130_fd_sc_hd__buf_4
XFILLER_0_96_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09573_ _03804_ VGND VGND VPWR VPWR _04864_ sky130_fd_sc_hd__buf_6
XFILLER_0_96_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_148_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09909_ _06319_ _06329_ _06267_ VGND VGND VPWR VPWR _08518_ sky130_fd_sc_hd__a21bo_1
X_12920_ _03012_ VGND VGND VPWR VPWR _03013_ sky130_fd_sc_hd__clkbuf_4
XTAP_2200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12851_ _00893_ _00897_ _00895_ VGND VGND VPWR VPWR _02944_ sky130_fd_sc_hd__a21oi_1
XTAP_2211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11802_ _01892_ _01893_ _01894_ VGND VGND VPWR VPWR _01895_ sky130_fd_sc_hd__nor3_1
XTAP_2244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15570_ _05884_ VGND VGND VPWR VPWR _05886_ sky130_fd_sc_hd__inv_2
XTAP_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12782_ _01374_ _02874_ VGND VGND VPWR VPWR _02875_ sky130_fd_sc_hd__nor2_1
XFILLER_0_68_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer90 _00925_ VGND VGND VPWR VPWR net337 sky130_fd_sc_hd__dlygate4sd1_1
XTAP_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14521_ _03005_ _00557_ VGND VGND VPWR VPWR _04743_ sky130_fd_sc_hd__nand2_1
XTAP_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11733_ _01824_ _01825_ VGND VGND VPWR VPWR _01826_ sky130_fd_sc_hd__or2b_1
XTAP_2299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17240_ _07678_ _07685_ _07696_ _07698_ VGND VGND VPWR VPWR _07699_ sky130_fd_sc_hd__or4b_1
X_14452_ _04650_ _04525_ _04666_ VGND VGND VPWR VPWR _04669_ sky130_fd_sc_hd__and3_1
XTAP_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11664_ _01610_ _01619_ _01708_ _01709_ VGND VGND VPWR VPWR _01757_ sky130_fd_sc_hd__o211a_1
XFILLER_0_154_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13403_ _03518_ _03519_ _03337_ _03339_ VGND VGND VPWR VPWR _03522_ sky130_fd_sc_hd__o211a_1
XFILLER_0_154_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10615_ _00564_ _00567_ _00565_ VGND VGND VPWR VPWR _00708_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_107_630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17171_ _02127_ _06814_ VGND VGND VPWR VPWR _07623_ sky130_fd_sc_hd__nor2_4
XFILLER_0_37_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14383_ _04590_ _04592_ VGND VGND VPWR VPWR _04593_ sky130_fd_sc_hd__xor2_1
X_11595_ _01684_ _01686_ _01685_ VGND VGND VPWR VPWR _01688_ sky130_fd_sc_hd__a21o_1
XFILLER_0_91_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16122_ _08865_ _02965_ _06422_ VGND VGND VPWR VPWR _06483_ sky130_fd_sc_hd__nor3_1
X_13334_ _03442_ _03445_ VGND VGND VPWR VPWR _03446_ sky130_fd_sc_hd__or2_1
X_10546_ _06084_ _07384_ _08158_ _06040_ VGND VGND VPWR VPWR _00639_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_51_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16053_ _03149_ VGND VGND VPWR VPWR _06408_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_106_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13265_ _00696_ net320 _03341_ _03342_ VGND VGND VPWR VPWR _03370_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_51_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10477_ _00568_ _00569_ VGND VGND VPWR VPWR _00570_ sky130_fd_sc_hd__xor2_1
XFILLER_0_121_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15004_ _05264_ _05270_ VGND VGND VPWR VPWR _05271_ sky130_fd_sc_hd__or2b_1
XFILLER_0_121_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12216_ _02277_ _02279_ _02274_ VGND VGND VPWR VPWR _02309_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_122_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13196_ _00737_ _00739_ VGND VGND VPWR VPWR _03297_ sky130_fd_sc_hd__or2b_1
XFILLER_0_20_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12147_ _02234_ _02239_ VGND VGND VPWR VPWR _02240_ sky130_fd_sc_hd__xnor2_1
X_12078_ _01995_ _01996_ _01999_ _02170_ VGND VGND VPWR VPWR _02171_ sky130_fd_sc_hd__o22ai_1
X_16955_ _06563_ _06756_ _07332_ _07387_ VGND VGND VPWR VPWR _07388_ sky130_fd_sc_hd__or4_1
X_11029_ _08039_ _04449_ _04471_ _00992_ VGND VGND VPWR VPWR _01122_ sky130_fd_sc_hd__a22o_1
X_15906_ _03013_ _06246_ _06248_ VGND VGND VPWR VPWR _06250_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_2_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16886_ _00247_ _07311_ _07312_ VGND VGND VPWR VPWR _07313_ sky130_fd_sc_hd__nand3_4
X_15837_ _06161_ _06174_ VGND VGND VPWR VPWR _06176_ sky130_fd_sc_hd__nor2_1
X_18625_ net303 _09157_ _09174_ _09162_ VGND VGND VPWR VPWR _00033_ sky130_fd_sc_hd__o211a_1
X_15768_ _02991_ _03153_ VGND VGND VPWR VPWR _06101_ sky130_fd_sc_hd__nand2_1
X_18556_ net68 _09096_ VGND VGND VPWR VPWR _09127_ sky130_fd_sc_hd__or2_2
XFILLER_0_86_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14719_ _03121_ _04959_ VGND VGND VPWR VPWR _04960_ sky130_fd_sc_hd__nor2_1
X_17507_ _07979_ _07989_ VGND VGND VPWR VPWR _07990_ sky130_fd_sc_hd__xnor2_1
X_18487_ _09018_ _09021_ _09019_ VGND VGND VPWR VPWR _09054_ sky130_fd_sc_hd__o21a_1
X_15699_ _03009_ _03012_ _09059_ _00322_ VGND VGND VPWR VPWR _06026_ sky130_fd_sc_hd__and4_1
X_17438_ _07910_ _07914_ _07912_ VGND VGND VPWR VPWR _07915_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_6_102 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_15 _01115_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_26 _01115_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_37 _01697_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_48 _02989_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17369_ _07833_ _07838_ VGND VGND VPWR VPWR _07839_ sky130_fd_sc_hd__xnor2_2
XANTENNA_59 _04406_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_734 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_144_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput100 net100 VGND VGND VPWR VPWR o_wb_data[25] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_30_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput111 net111 VGND VGND VPWR VPWR o_wb_data[6] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09625_ _05344_ _05421_ VGND VGND VPWR VPWR _05431_ sky130_fd_sc_hd__and2b_1
X_09556_ _04438_ _04482_ _04657_ _04646_ VGND VGND VPWR VPWR _04679_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_78_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09487_ _03881_ _03892_ _03903_ _03914_ VGND VGND VPWR VPWR _03925_ sky130_fd_sc_hd__and4_1
XFILLER_0_38_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_111 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_148_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_148_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_136_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10400_ _00340_ _00347_ VGND VGND VPWR VPWR _00493_ sky130_fd_sc_hd__nand2_1
XFILLER_0_61_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11380_ _01470_ _01472_ VGND VGND VPWR VPWR _01473_ sky130_fd_sc_hd__xor2_1
XFILLER_0_150_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10331_ _00378_ _00421_ _00422_ _00423_ VGND VGND VPWR VPWR _00424_ sky130_fd_sc_hd__and4b_2
XFILLER_0_103_132 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_104_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10262_ _00353_ _09271_ _00354_ VGND VGND VPWR VPWR _00355_ sky130_fd_sc_hd__or3_1
X_13050_ _00322_ VGND VGND VPWR VPWR _03142_ sky130_fd_sc_hd__buf_2
X_12001_ _05410_ _05301_ _00146_ _00197_ VGND VGND VPWR VPWR _02094_ sky130_fd_sc_hd__nand4_1
X_10193_ _00284_ _00285_ VGND VGND VPWR VPWR _00286_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_100_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16740_ _07152_ _07153_ VGND VGND VPWR VPWR _07154_ sky130_fd_sc_hd__xnor2_2
X_13952_ _04107_ _04108_ _04119_ VGND VGND VPWR VPWR _04122_ sky130_fd_sc_hd__or3_4
X_12903_ _00191_ VGND VGND VPWR VPWR _02996_ sky130_fd_sc_hd__clkbuf_4
X_16671_ _06462_ _07078_ VGND VGND VPWR VPWR _07079_ sky130_fd_sc_hd__nor2_1
X_13883_ _04043_ _04044_ _03828_ _04007_ VGND VGND VPWR VPWR _04047_ sky130_fd_sc_hd__o211a_1
X_15622_ _05941_ _05942_ VGND VGND VPWR VPWR _05944_ sky130_fd_sc_hd__and2_1
X_18410_ _08969_ _08970_ VGND VGND VPWR VPWR _08971_ sky130_fd_sc_hd__or2_1
X_12834_ _02924_ _02925_ _02923_ _02907_ VGND VGND VPWR VPWR _02927_ sky130_fd_sc_hd__a211o_1
XTAP_2030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18341_ _08895_ _04023_ _07743_ VGND VGND VPWR VPWR _08896_ sky130_fd_sc_hd__or3_1
X_15553_ _05864_ _05865_ _05776_ _05778_ VGND VGND VPWR VPWR _05869_ sky130_fd_sc_hd__a211o_1
XTAP_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12765_ _01790_ _02855_ _02856_ _02857_ VGND VGND VPWR VPWR _02858_ sky130_fd_sc_hd__o211a_1
XTAP_2085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_336 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14504_ _04515_ VGND VGND VPWR VPWR _04725_ sky130_fd_sc_hd__buf_4
XTAP_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18272_ _05557_ _06401_ _06400_ VGND VGND VPWR VPWR _08823_ sky130_fd_sc_hd__a21oi_1
X_11716_ _01806_ _01807_ _01507_ VGND VGND VPWR VPWR _01809_ sky130_fd_sc_hd__a21oi_1
XTAP_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15484_ _05616_ _05790_ VGND VGND VPWR VPWR _05794_ sky130_fd_sc_hd__nand2_1
X_12696_ _02782_ _02786_ _02787_ _02788_ VGND VGND VPWR VPWR _02789_ sky130_fd_sc_hd__and4_1
XFILLER_0_126_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17223_ _06368_ _07355_ _04725_ VGND VGND VPWR VPWR _07681_ sky130_fd_sc_hd__or3b_1
X_14435_ _04325_ _04523_ VGND VGND VPWR VPWR _04650_ sky130_fd_sc_hd__or2_1
XFILLER_0_115_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11647_ _01721_ _01738_ _01737_ VGND VGND VPWR VPWR _01740_ sky130_fd_sc_hd__a21o_1
Xinput13 i_wb_addr[1] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput24 i_wb_addr[2] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__buf_2
XFILLER_0_25_756 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17154_ _06657_ _07604_ _07498_ VGND VGND VPWR VPWR _07605_ sky130_fd_sc_hd__and3_1
Xinput35 i_wb_data[0] VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_4_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14366_ _04571_ _04572_ _04567_ net333 VGND VGND VPWR VPWR _04574_ sky130_fd_sc_hd__a211o_1
Xinput46 i_wb_data[1] VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__clkbuf_4
X_11578_ _05878_ VGND VGND VPWR VPWR _01671_ sky130_fd_sc_hd__clkinv_4
XFILLER_0_107_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput57 i_wb_data[2] VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__clkbuf_4
Xinput68 i_wb_we VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__buf_4
XFILLER_0_40_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16105_ _06463_ VGND VGND VPWR VPWR _06464_ sky130_fd_sc_hd__clkbuf_4
X_13317_ _03424_ _03425_ _03411_ VGND VGND VPWR VPWR _03427_ sky130_fd_sc_hd__a21oi_2
X_10529_ _00451_ _00453_ VGND VGND VPWR VPWR _00622_ sky130_fd_sc_hd__nand2_1
X_17085_ _07510_ _07529_ VGND VGND VPWR VPWR _07530_ sky130_fd_sc_hd__xor2_1
X_14297_ _04497_ _04498_ VGND VGND VPWR VPWR _04499_ sky130_fd_sc_hd__xnor2_1
X_16036_ _06386_ _06387_ _06388_ VGND VGND VPWR VPWR _06389_ sky130_fd_sc_hd__a21bo_1
X_13248_ _00713_ _00717_ _00712_ VGND VGND VPWR VPWR _03352_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_149_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13179_ _03276_ _03277_ VGND VGND VPWR VPWR _03278_ sky130_fd_sc_hd__and2_1
X_17987_ _03044_ _08428_ _03000_ VGND VGND VPWR VPWR _08513_ sky130_fd_sc_hd__or3b_2
X_16938_ _06704_ _06710_ _03079_ VGND VGND VPWR VPWR _07370_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_88 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16869_ _07292_ _07293_ VGND VGND VPWR VPWR _07294_ sky130_fd_sc_hd__xnor2_2
X_18608_ salida\[21\] _09159_ _09160_ salida\[53\] _09163_ VGND VGND VPWR VPWR _09164_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_59_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18539_ net148 VGND VGND VPWR VPWR _09109_ sky130_fd_sc_hd__inv_2
XFILLER_0_74_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_118_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_522 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_214 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_141_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_4_5_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_5_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_3_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09608_ cla_inst.in1\[20\] VGND VGND VPWR VPWR _05246_ sky130_fd_sc_hd__clkbuf_8
X_10880_ _00969_ _00972_ VGND VGND VPWR VPWR _00973_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_85_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09539_ ApproximateM_inst.lob_16.lob2.genblk1\[13\].genblk1.mux.sel VGND VGND VPWR
+ VPWR _04493_ sky130_fd_sc_hd__buf_4
XFILLER_0_109_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12550_ _02635_ _02641_ _02642_ VGND VGND VPWR VPWR _02643_ sky130_fd_sc_hd__and3_1
XFILLER_0_19_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11501_ _01589_ _01592_ VGND VGND VPWR VPWR _01594_ sky130_fd_sc_hd__xor2_1
XFILLER_0_93_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_108_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12481_ _02571_ _02573_ _02504_ VGND VGND VPWR VPWR _02574_ sky130_fd_sc_hd__a21o_1
XFILLER_0_62_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14220_ _02975_ _04413_ VGND VGND VPWR VPWR _04414_ sky130_fd_sc_hd__nor2_2
X_11432_ _01514_ _01524_ VGND VGND VPWR VPWR _01525_ sky130_fd_sc_hd__or2_1
XFILLER_0_62_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14151_ _00192_ _06482_ _05921_ _00190_ VGND VGND VPWR VPWR _04339_ sky130_fd_sc_hd__a22oi_1
X_11363_ _01396_ _01404_ _01397_ _01398_ VGND VGND VPWR VPWR _01456_ sky130_fd_sc_hd__or4_1
XFILLER_0_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13102_ _03194_ VGND VGND VPWR VPWR _03196_ sky130_fd_sc_hd__inv_2
X_10314_ _00405_ _00406_ VGND VGND VPWR VPWR _00407_ sky130_fd_sc_hd__and2b_1
X_14082_ _03547_ _04262_ VGND VGND VPWR VPWR _04264_ sky130_fd_sc_hd__nor2_1
X_11294_ _01385_ _01284_ _01386_ VGND VGND VPWR VPWR _01387_ sky130_fd_sc_hd__a21o_2
XFILLER_0_131_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_770 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17910_ _04336_ _08428_ _03368_ VGND VGND VPWR VPWR _08429_ sky130_fd_sc_hd__or3b_1
X_13033_ _03124_ VGND VGND VPWR VPWR _03125_ sky130_fd_sc_hd__clkbuf_4
X_10245_ _09070_ _09137_ VGND VGND VPWR VPWR _00338_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_792 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18890_ clknet_4_13_0_clk _00044_ VGND VGND VPWR VPWR ApproximateM_inst.lob_16.lob1.genblk1\[8\].genblk1.mux.sel
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_28_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10176_ _00267_ _00266_ _08289_ _07919_ VGND VGND VPWR VPWR _00269_ sky130_fd_sc_hd__a211oi_2
X_17841_ _08351_ _08352_ VGND VGND VPWR VPWR _08353_ sky130_fd_sc_hd__nand2_1
X_14984_ _03321_ _06094_ _00460_ _03322_ VGND VGND VPWR VPWR _05249_ sky130_fd_sc_hd__a22oi_1
X_17772_ _08176_ _08177_ _08175_ VGND VGND VPWR VPWR _08279_ sky130_fd_sc_hd__o21ai_1
X_13935_ _04101_ _04102_ VGND VGND VPWR VPWR _04103_ sky130_fd_sc_hd__nand2_1
X_16723_ _07031_ _07044_ _07135_ VGND VGND VPWR VPWR _07136_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_88_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16654_ _06967_ _06975_ _07060_ VGND VGND VPWR VPWR _07061_ sky130_fd_sc_hd__o21ai_1
X_13866_ _03863_ _03871_ _04027_ VGND VGND VPWR VPWR _04028_ sky130_fd_sc_hd__a21bo_1
X_15605_ _05915_ _05923_ VGND VGND VPWR VPWR _05925_ sky130_fd_sc_hd__and2_1
X_12817_ _02907_ _02908_ _01468_ _01490_ VGND VGND VPWR VPWR _02910_ sky130_fd_sc_hd__o211a_1
XFILLER_0_97_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16585_ _06984_ _06985_ VGND VGND VPWR VPWR _06986_ sky130_fd_sc_hd__xor2_1
X_13797_ _05975_ _03763_ _03765_ _03766_ VGND VGND VPWR VPWR _03952_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_96_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15536_ _07668_ _00318_ _05758_ _03009_ VGND VGND VPWR VPWR _05850_ sky130_fd_sc_hd__a22o_1
X_18324_ _02887_ _08877_ VGND VGND VPWR VPWR _08879_ sky130_fd_sc_hd__nand2_1
XFILLER_0_45_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12748_ _02838_ _02840_ _02837_ VGND VGND VPWR VPWR _02841_ sky130_fd_sc_hd__a21o_1
XTAP_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_127_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18255_ _08802_ _08803_ VGND VGND VPWR VPWR _08804_ sky130_fd_sc_hd__and2_1
X_15467_ _05773_ _05757_ _05759_ VGND VGND VPWR VPWR _05775_ sky130_fd_sc_hd__and3_1
XFILLER_0_5_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12679_ _02769_ _02771_ VGND VGND VPWR VPWR _02772_ sky130_fd_sc_hd__and2_1
XFILLER_0_37_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17206_ _07538_ _07545_ _07536_ VGND VGND VPWR VPWR _07662_ sky130_fd_sc_hd__o21ba_1
X_14418_ _01504_ _05856_ _04497_ VGND VGND VPWR VPWR _04631_ sky130_fd_sc_hd__and3_1
XFILLER_0_114_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18186_ _08727_ _08728_ VGND VGND VPWR VPWR _08729_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_154_396 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15398_ _05596_ _05699_ VGND VGND VPWR VPWR _05700_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_8_36 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_558 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_512 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_107_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17137_ _07549_ _07551_ VGND VGND VPWR VPWR _07586_ sky130_fd_sc_hd__and2b_1
X_14349_ _04552_ _04554_ _04555_ VGND VGND VPWR VPWR _04556_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_69_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17068_ _04012_ _06889_ VGND VGND VPWR VPWR _07511_ sky130_fd_sc_hd__nand2_4
XFILLER_0_122_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16019_ _06367_ _06369_ _00786_ VGND VGND VPWR VPWR _06370_ sky130_fd_sc_hd__a21bo_1
XTAP_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09890_ _06949_ _08278_ _08289_ _08300_ VGND VGND VPWR VPWR _08311_ sky130_fd_sc_hd__or4b_4
XTAP_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_83 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_612 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_137_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_103 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10030_ _08191_ _00122_ VGND VGND VPWR VPWR _00123_ sky130_fd_sc_hd__nor2_2
XFILLER_0_98_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11981_ _01967_ _02027_ _02052_ VGND VGND VPWR VPWR _02074_ sky130_fd_sc_hd__or3_1
X_13720_ cla_inst.in2\[25\] _04012_ VGND VGND VPWR VPWR _03868_ sky130_fd_sc_hd__nand2_1
X_10932_ _03771_ _04242_ _00176_ _04078_ VGND VGND VPWR VPWR _01025_ sky130_fd_sc_hd__a22o_1
XFILLER_0_105_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13651_ _06040_ _06084_ _00509_ _00513_ VGND VGND VPWR VPWR _03792_ sky130_fd_sc_hd__and4_1
XFILLER_0_79_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10863_ _04078_ _03771_ _00949_ _03421_ VGND VGND VPWR VPWR _00956_ sky130_fd_sc_hd__and4_1
XFILLER_0_85_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12602_ _02654_ _02660_ _02661_ VGND VGND VPWR VPWR _02695_ sky130_fd_sc_hd__a21oi_1
XPHY_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16370_ net212 _06517_ _06520_ _06751_ VGND VGND VPWR VPWR _06752_ sky130_fd_sc_hd__o22a_1
XFILLER_0_94_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13582_ _03676_ _03677_ _03715_ _03716_ VGND VGND VPWR VPWR _03718_ sky130_fd_sc_hd__o211a_1
X_10794_ _00868_ _00886_ VGND VGND VPWR VPWR _00887_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_94_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15321_ _05520_ _05516_ _05517_ VGND VGND VPWR VPWR _05616_ sky130_fd_sc_hd__o21a_1
XFILLER_0_93_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_330 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_137_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12533_ _02622_ _02624_ VGND VGND VPWR VPWR _02626_ sky130_fd_sc_hd__nand2_1
XPHY_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18040_ _08568_ _08569_ VGND VGND VPWR VPWR _08570_ sky130_fd_sc_hd__nand2_1
X_15252_ _05538_ _01139_ _05449_ _05539_ VGND VGND VPWR VPWR _05541_ sky130_fd_sc_hd__and4b_1
XFILLER_0_109_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12464_ _02550_ _02556_ VGND VGND VPWR VPWR _02557_ sky130_fd_sc_hd__and2_1
XFILLER_0_136_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14203_ _04393_ _04394_ _04396_ VGND VGND VPWR VPWR _04397_ sky130_fd_sc_hd__or3_4
XFILLER_0_35_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11415_ _03662_ _07591_ VGND VGND VPWR VPWR _01508_ sky130_fd_sc_hd__nand2_2
XFILLER_0_124_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15183_ _09350_ _05715_ _05975_ _00112_ VGND VGND VPWR VPWR _05466_ sky130_fd_sc_hd__a22oi_1
X_12395_ _05671_ _00197_ _02486_ _02487_ _09188_ VGND VGND VPWR VPWR _02488_ sky130_fd_sc_hd__a32oi_4
XFILLER_0_105_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14134_ _00678_ _04045_ _04067_ _00679_ VGND VGND VPWR VPWR _04321_ sky130_fd_sc_hd__a22o_1
X_11346_ _01413_ _01414_ _01312_ _01378_ VGND VGND VPWR VPWR _01439_ sky130_fd_sc_hd__o211a_1
XFILLER_0_22_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18942_ clknet_4_2_0_clk _00096_ VGND VGND VPWR VPWR cla_inst.in2\[28\] sky130_fd_sc_hd__dfxtp_1
X_14065_ _03540_ _03554_ _02980_ VGND VGND VPWR VPWR _04246_ sky130_fd_sc_hd__mux2_1
X_11277_ _01238_ _01273_ _01368_ _01369_ VGND VGND VPWR VPWR _01370_ sky130_fd_sc_hd__o211a_1
X_13016_ _03025_ _03108_ _02272_ VGND VGND VPWR VPWR _03109_ sky130_fd_sc_hd__a21o_1
X_10228_ _05747_ _07025_ _00317_ _00320_ VGND VGND VPWR VPWR _00321_ sky130_fd_sc_hd__and4_1
X_18873_ clknet_4_14_0_clk net246 VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__dfxtp_1
X_17824_ _06388_ _06387_ _06386_ VGND VGND VPWR VPWR _08336_ sky130_fd_sc_hd__a21o_1
X_10159_ _00203_ _00166_ VGND VGND VPWR VPWR _00252_ sky130_fd_sc_hd__nand2_1
XFILLER_0_55_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14967_ _00678_ _00443_ _06471_ _00679_ VGND VGND VPWR VPWR _05230_ sky130_fd_sc_hd__a22o_1
X_17755_ _07933_ VGND VGND VPWR VPWR _08260_ sky130_fd_sc_hd__buf_2
XFILLER_0_89_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16706_ _06766_ _06875_ _07114_ _07116_ VGND VGND VPWR VPWR _07117_ sky130_fd_sc_hd__nor4_1
X_13918_ _04080_ _04084_ _03921_ VGND VGND VPWR VPWR _04085_ sky130_fd_sc_hd__mux2_1
X_17686_ _08183_ _08184_ VGND VGND VPWR VPWR _08185_ sky130_fd_sc_hd__or2b_1
X_14898_ _05009_ _05154_ VGND VGND VPWR VPWR _05155_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_77_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13849_ _00173_ _00175_ _04460_ _04482_ VGND VGND VPWR VPWR _04009_ sky130_fd_sc_hd__and4_2
X_16637_ _06957_ VGND VGND VPWR VPWR _07042_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_76_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_147_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_528 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16568_ _06939_ _06966_ VGND VGND VPWR VPWR _06967_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_45_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18307_ _08858_ _08844_ VGND VGND VPWR VPWR _08860_ sky130_fd_sc_hd__and2b_1
XFILLER_0_45_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15519_ _05746_ _05745_ VGND VGND VPWR VPWR _05831_ sky130_fd_sc_hd__or2b_1
X_16499_ _06801_ _06818_ VGND VGND VPWR VPWR _06892_ sky130_fd_sc_hd__nor2_1
XFILLER_0_127_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18238_ _08707_ _08710_ _08783_ VGND VGND VPWR VPWR _08785_ sky130_fd_sc_hd__a21o_1
XFILLER_0_32_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18169_ _08704_ _08708_ VGND VGND VPWR VPWR _08710_ sky130_fd_sc_hd__nand2_1
XFILLER_0_143_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_cap121 _03884_ VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__buf_1
XFILLER_0_20_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_cap143 _00603_ VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__buf_1
X_09942_ _07123_ VGND VGND VPWR VPWR _08876_ sky130_fd_sc_hd__buf_4
XFILLER_0_96_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09873_ _07319_ _07940_ _08115_ VGND VGND VPWR VPWR _08126_ sky130_fd_sc_hd__nand3_4
XTAP_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_118_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_119_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11200_ _00968_ _00973_ VGND VGND VPWR VPWR _01293_ sky130_fd_sc_hd__nand2_1
X_12180_ _00846_ _00716_ _02272_ VGND VGND VPWR VPWR _02273_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_31_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11131_ _00515_ _01136_ VGND VGND VPWR VPWR _01224_ sky130_fd_sc_hd__nor2_4
XFILLER_0_101_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11062_ _04984_ _00218_ VGND VGND VPWR VPWR _01155_ sky130_fd_sc_hd__nand2_1
X_10013_ cla_inst.in2\[25\] VGND VGND VPWR VPWR _00106_ sky130_fd_sc_hd__clkbuf_4
X_15870_ _06209_ _06210_ VGND VGND VPWR VPWR _06211_ sky130_fd_sc_hd__nor2_1
XFILLER_0_99_810 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14821_ _04896_ _04963_ _05069_ _05070_ VGND VGND VPWR VPWR _05071_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_116_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14752_ _04725_ _04125_ _04994_ VGND VGND VPWR VPWR _04996_ sky130_fd_sc_hd__and3_2
X_17540_ _07911_ _07912_ _07910_ VGND VGND VPWR VPWR _08026_ sky130_fd_sc_hd__a21o_1
X_11964_ _02006_ _02001_ _02004_ VGND VGND VPWR VPWR _02057_ sky130_fd_sc_hd__or3_1
XFILLER_0_59_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13703_ _03847_ _03849_ VGND VGND VPWR VPWR _03850_ sky130_fd_sc_hd__nand2_1
X_10915_ _05671_ _05322_ VGND VGND VPWR VPWR _01008_ sky130_fd_sc_hd__nand2_1
XFILLER_0_58_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17471_ _07942_ _07949_ VGND VGND VPWR VPWR _07950_ sky130_fd_sc_hd__xor2_1
X_14683_ _04917_ _04918_ _04903_ _04791_ VGND VGND VPWR VPWR _04921_ sky130_fd_sc_hd__o211ai_1
X_11895_ _01675_ _01864_ _01981_ VGND VGND VPWR VPWR _01988_ sky130_fd_sc_hd__or3_1
XFILLER_0_129_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13634_ _03612_ _03613_ VGND VGND VPWR VPWR _03774_ sky130_fd_sc_hd__nand2_2
X_16422_ _07657_ _06541_ _06807_ VGND VGND VPWR VPWR _06809_ sky130_fd_sc_hd__and3_1
X_10846_ _00932_ _00933_ _00937_ VGND VGND VPWR VPWR _00939_ sky130_fd_sc_hd__nand3_1
XFILLER_0_82_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_650 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16353_ _06727_ _06733_ _03079_ VGND VGND VPWR VPWR _06734_ sky130_fd_sc_hd__mux2_2
X_13565_ _03496_ _03502_ VGND VGND VPWR VPWR _03699_ sky130_fd_sc_hd__nand2_1
Xsplit84 _06571_ VGND VGND VPWR VPWR net331 sky130_fd_sc_hd__dlymetal6s2s_1
X_10777_ _00200_ _00869_ VGND VGND VPWR VPWR _00870_ sky130_fd_sc_hd__or2_1
XFILLER_0_54_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15304_ _05552_ _05596_ _05597_ VGND VGND VPWR VPWR _05598_ sky130_fd_sc_hd__or3_1
XFILLER_0_82_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12516_ _02608_ _02559_ VGND VGND VPWR VPWR _02609_ sky130_fd_sc_hd__or2b_1
XFILLER_0_26_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16284_ _06654_ _06658_ VGND VGND VPWR VPWR _06659_ sky130_fd_sc_hd__and2_1
X_13496_ _03620_ _03621_ _03393_ _03587_ VGND VGND VPWR VPWR _03623_ sky130_fd_sc_hd__a211o_4
XFILLER_0_136_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15235_ _05518_ _05521_ _05522_ VGND VGND VPWR VPWR _05523_ sky130_fd_sc_hd__a21o_1
X_18023_ _07194_ _07290_ _07511_ _07621_ VGND VGND VPWR VPWR _08552_ sky130_fd_sc_hd__or4_1
X_12447_ _02538_ _02539_ VGND VGND VPWR VPWR _02540_ sky130_fd_sc_hd__or2_1
XFILLER_0_125_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15166_ _05445_ _05446_ VGND VGND VPWR VPWR _05447_ sky130_fd_sc_hd__nor2_1
X_12378_ _02400_ _02461_ VGND VGND VPWR VPWR _02471_ sky130_fd_sc_hd__xor2_2
X_14117_ _04115_ _04109_ VGND VGND VPWR VPWR _04302_ sky130_fd_sc_hd__and2b_1
X_11329_ cla_inst.in2\[20\] _00878_ VGND VGND VPWR VPWR _01422_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15097_ _01505_ _00322_ VGND VGND VPWR VPWR _05372_ sky130_fd_sc_hd__nand2_1
XFILLER_0_120_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14048_ _04052_ _04055_ VGND VGND VPWR VPWR _04227_ sky130_fd_sc_hd__or2b_1
X_18925_ clknet_4_11_0_clk _00079_ VGND VGND VPWR VPWR ApproximateM_inst.lob_16.lob2.genblk1\[11\].genblk1.mux.sel
+ sky130_fd_sc_hd__dfxtp_4
X_18856_ clknet_4_4_0_clk net256 VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__dfxtp_1
X_17807_ _08187_ _08200_ _08198_ VGND VGND VPWR VPWR _08317_ sky130_fd_sc_hd__a21o_1
X_18787_ _02985_ net45 _09276_ VGND VGND VPWR VPWR _09299_ sky130_fd_sc_hd__mux2_1
X_15999_ _07058_ _01264_ VGND VGND VPWR VPWR _06348_ sky130_fd_sc_hd__or2_2
XFILLER_0_89_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17738_ _06385_ _06546_ _08241_ _01678_ VGND VGND VPWR VPWR _08242_ sky130_fd_sc_hd__a22o_1
XFILLER_0_82_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17669_ _08159_ _08164_ VGND VGND VPWR VPWR _08166_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_116_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_670 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09925_ _06384_ _06439_ VGND VGND VPWR VPWR _08692_ sky130_fd_sc_hd__or2b_1
XTAP_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09856_ _07210_ _07308_ _07297_ VGND VGND VPWR VPWR _07940_ sky130_fd_sc_hd__a21o_1
XTAP_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09787_ _05736_ _05986_ _06105_ _06073_ VGND VGND VPWR VPWR _07189_ sky130_fd_sc_hd__a31o_1
XTAP_2404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_105 _09403_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_116 _00131_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_127 _03790_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_138 _05888_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_149 _08762_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_139_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10700_ _00762_ _00763_ _00778_ VGND VGND VPWR VPWR _00793_ sky130_fd_sc_hd__a21o_1
XTAP_1747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11680_ cla_inst.in2\[20\] _01503_ _01240_ _01506_ VGND VGND VPWR VPWR _01773_ sky130_fd_sc_hd__a22o_1
XTAP_1769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10631_ _09353_ _00207_ _00548_ _00547_ VGND VGND VPWR VPWR _00724_ sky130_fd_sc_hd__a31o_1
X_13350_ _03449_ _03462_ VGND VGND VPWR VPWR _03463_ sky130_fd_sc_hd__xnor2_1
X_10562_ _00638_ _00653_ _00654_ VGND VGND VPWR VPWR _00655_ sky130_fd_sc_hd__nand3b_2
XFILLER_0_118_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12301_ _02390_ _02391_ _02385_ net123 VGND VGND VPWR VPWR _02394_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_133_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13281_ _03728_ _06062_ VGND VGND VPWR VPWR _03387_ sky130_fd_sc_hd__nand2_1
XFILLER_0_107_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10493_ _00583_ _00584_ net339 _00424_ VGND VGND VPWR VPWR _00586_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_121_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15020_ _05243_ _05287_ VGND VGND VPWR VPWR _05288_ sky130_fd_sc_hd__xor2_2
XFILLER_0_121_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12232_ _02323_ _02324_ VGND VGND VPWR VPWR _02325_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_20_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12163_ _02254_ _02255_ VGND VGND VPWR VPWR _02256_ sky130_fd_sc_hd__nand2_1
XFILLER_0_130_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11114_ _07254_ _05039_ _00439_ _07232_ VGND VGND VPWR VPWR _01207_ sky130_fd_sc_hd__a22o_1
X_12094_ _02185_ _02186_ VGND VGND VPWR VPWR _02187_ sky130_fd_sc_hd__nand2_1
X_16971_ _07392_ _07404_ VGND VGND VPWR VPWR _07405_ sky130_fd_sc_hd__xnor2_1
X_18710_ net54 _03068_ _09182_ VGND VGND VPWR VPWR _09238_ sky130_fd_sc_hd__mux2_1
X_11045_ _01109_ _01137_ VGND VGND VPWR VPWR _01138_ sky130_fd_sc_hd__nand2_1
X_15922_ _04958_ _05307_ _06266_ _03039_ VGND VGND VPWR VPWR _06268_ sky130_fd_sc_hd__o22a_1
X_18641_ _09187_ VGND VGND VPWR VPWR _00037_ sky130_fd_sc_hd__clkbuf_1
X_15853_ _06118_ _06173_ VGND VGND VPWR VPWR _06193_ sky130_fd_sc_hd__and2b_1
X_14804_ _05051_ _05052_ VGND VGND VPWR VPWR _05053_ sky130_fd_sc_hd__nand2_1
X_18572_ salida\[8\] _09114_ _09118_ salida\[40\] _09128_ VGND VGND VPWR VPWR _09138_
+ sky130_fd_sc_hd__a221o_1
X_15784_ _06098_ _06099_ _06117_ VGND VGND VPWR VPWR _06119_ sky130_fd_sc_hd__or3_1
X_12996_ _03047_ VGND VGND VPWR VPWR _03089_ sky130_fd_sc_hd__clkbuf_4
X_17523_ _07999_ _08007_ VGND VGND VPWR VPWR _08008_ sky130_fd_sc_hd__xnor2_1
X_14735_ _04034_ _00502_ _09311_ _04099_ VGND VGND VPWR VPWR _04977_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_52_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11947_ _02035_ _02038_ VGND VGND VPWR VPWR _02040_ sky130_fd_sc_hd__and2b_1
XFILLER_0_52_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17454_ _07896_ _07898_ VGND VGND VPWR VPWR _07932_ sky130_fd_sc_hd__nor2_1
X_14666_ _04899_ _04901_ VGND VGND VPWR VPWR _04902_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_28_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11878_ _01969_ _01938_ _01970_ _01869_ VGND VGND VPWR VPWR _01971_ sky130_fd_sc_hd__o211a_1
XFILLER_0_27_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13617_ _03366_ cla_inst.in1\[20\] _05377_ _03345_ VGND VGND VPWR VPWR _03755_ sky130_fd_sc_hd__a22o_1
X_16405_ _03083_ _06430_ VGND VGND VPWR VPWR _06791_ sky130_fd_sc_hd__nor2_1
X_10829_ _00920_ _00921_ VGND VGND VPWR VPWR _00922_ sky130_fd_sc_hd__and2b_1
X_14597_ _03543_ _03555_ _02979_ VGND VGND VPWR VPWR _04827_ sky130_fd_sc_hd__mux2_1
X_17385_ _07727_ _07719_ VGND VGND VPWR VPWR _07857_ sky130_fd_sc_hd__and2b_1
X_13548_ _03678_ _03679_ VGND VGND VPWR VPWR _03680_ sky130_fd_sc_hd__nor2_1
X_16336_ _03077_ _06715_ VGND VGND VPWR VPWR _06716_ sky130_fd_sc_hd__and2_1
XFILLER_0_42_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_125_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16267_ _06467_ _06640_ VGND VGND VPWR VPWR _06641_ sky130_fd_sc_hd__and2_1
X_13479_ net330 _03597_ _03602_ VGND VGND VPWR VPWR _03604_ sky130_fd_sc_hd__a21o_1
XFILLER_0_70_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15218_ _05429_ _05390_ _05502_ VGND VGND VPWR VPWR _05504_ sky130_fd_sc_hd__or3_1
X_18006_ _07313_ _07487_ _07593_ _07318_ VGND VGND VPWR VPWR _08533_ sky130_fd_sc_hd__o22a_1
XFILLER_0_140_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16198_ ApproximateM_inst.lob_16.lob1.genblk1\[12\].genblk1.mux.sel _03826_ sel_op\[2\]
+ VGND VGND VPWR VPWR _06565_ sky130_fd_sc_hd__or3b_1
X_15149_ _05390_ _05391_ _05394_ VGND VGND VPWR VPWR _05428_ sky130_fd_sc_hd__or3_1
X_09710_ _06267_ _06329_ _06319_ VGND VGND VPWR VPWR _06351_ sky130_fd_sc_hd__a21o_1
X_18908_ clknet_4_10_0_clk _00062_ VGND VGND VPWR VPWR cla_inst.in1\[26\] sky130_fd_sc_hd__dfxtp_1
X_09641_ cla_inst.in1\[22\] VGND VGND VPWR VPWR _05606_ sky130_fd_sc_hd__buf_4
X_18839_ clknet_4_0_0_clk net302 VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__dfxtp_1
X_09572_ _03990_ _04482_ VGND VGND VPWR VPWR _04853_ sky130_fd_sc_hd__nand2_8
XFILLER_0_78_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_94 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_148_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_242 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_116_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_848 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_130_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_358 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_112_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_130_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09908_ _08398_ _08485_ _08474_ VGND VGND VPWR VPWR _08507_ sky130_fd_sc_hd__a21o_1
X_09839_ cla_inst.in1\[29\] VGND VGND VPWR VPWR _07755_ sky130_fd_sc_hd__clkbuf_4
X_12850_ _00893_ _00895_ _00897_ VGND VGND VPWR VPWR _02943_ sky130_fd_sc_hd__and3_1
XTAP_2201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11801_ _01707_ _01891_ _01887_ _01890_ VGND VGND VPWR VPWR _01894_ sky130_fd_sc_hd__o211a_1
XTAP_2234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12781_ _01370_ _01373_ _01371_ _01372_ VGND VGND VPWR VPWR _02874_ sky130_fd_sc_hd__o211a_1
XTAP_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer80 _04683_ VGND VGND VPWR VPWR net243 sky130_fd_sc_hd__clkbuf_1
XTAP_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer91 _00375_ VGND VGND VPWR VPWR net338 sky130_fd_sc_hd__clkbuf_1
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14520_ _04739_ _04740_ _04598_ _04701_ VGND VGND VPWR VPWR _04742_ sky130_fd_sc_hd__o211ai_4
XTAP_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11732_ _01816_ _01819_ VGND VGND VPWR VPWR _01825_ sky130_fd_sc_hd__xnor2_1
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14451_ _04650_ _04525_ _04666_ VGND VGND VPWR VPWR _04667_ sky130_fd_sc_hd__a21oi_2
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11663_ _01741_ _01754_ _01755_ VGND VGND VPWR VPWR _01756_ sky130_fd_sc_hd__nand3_2
XFILLER_0_37_743 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13402_ _03337_ _03339_ _03518_ _03519_ VGND VGND VPWR VPWR _03521_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_153_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10614_ _00705_ _00706_ VGND VGND VPWR VPWR _00707_ sky130_fd_sc_hd__xnor2_2
X_17170_ _06561_ _07124_ _07318_ _07621_ VGND VGND VPWR VPWR _07622_ sky130_fd_sc_hd__or4_1
XFILLER_0_36_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14382_ _06460_ _03455_ VGND VGND VPWR VPWR _04592_ sky130_fd_sc_hd__nand2_1
X_11594_ _01684_ _01685_ _01686_ VGND VGND VPWR VPWR _01687_ sky130_fd_sc_hd__nand3_2
XFILLER_0_36_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16121_ _04241_ _06474_ _06480_ _03117_ VGND VGND VPWR VPWR _06481_ sky130_fd_sc_hd__a211o_1
XFILLER_0_153_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13333_ _00362_ _00207_ _03441_ _03444_ VGND VGND VPWR VPWR _03445_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_24_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10545_ _00457_ _00462_ _00456_ VGND VGND VPWR VPWR _00638_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_52_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16052_ _06404_ _06405_ VGND VGND VPWR VPWR _06407_ sky130_fd_sc_hd__nand2_1
XFILLER_0_134_494 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13264_ _03368_ _03311_ _03310_ VGND VGND VPWR VPWR _03369_ sky130_fd_sc_hd__nand3_2
XFILLER_0_122_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10476_ _00253_ _00166_ _00406_ _00405_ VGND VGND VPWR VPWR _00569_ sky130_fd_sc_hd__a31o_1
XFILLER_0_121_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15003_ _05267_ _05269_ VGND VGND VPWR VPWR _05270_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_122_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12215_ _02295_ _02299_ _02306_ _02307_ VGND VGND VPWR VPWR _02308_ sky130_fd_sc_hd__o211a_1
X_13195_ _03293_ _03294_ _00661_ net327 VGND VGND VPWR VPWR _03296_ sky130_fd_sc_hd__a211o_4
X_12146_ _02235_ _02238_ VGND VGND VPWR VPWR _02239_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_138_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12077_ _02081_ _02167_ _02169_ VGND VGND VPWR VPWR _02170_ sky130_fd_sc_hd__o21ai_1
X_16954_ _06374_ _03324_ _06814_ _07386_ VGND VGND VPWR VPWR _07387_ sky130_fd_sc_hd__a211o_2
X_11028_ _01097_ _01101_ VGND VGND VPWR VPWR _01121_ sky130_fd_sc_hd__xnor2_1
X_15905_ _03013_ _06246_ _06248_ VGND VGND VPWR VPWR _06249_ sky130_fd_sc_hd__and3_1
X_16885_ _02124_ _06871_ VGND VGND VPWR VPWR _07312_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18624_ salida\[29\] _09159_ _09160_ salida\[61\] _09163_ VGND VGND VPWR VPWR _09174_
+ sky130_fd_sc_hd__a221o_1
X_15836_ _06161_ _06174_ VGND VGND VPWR VPWR _06175_ sky130_fd_sc_hd__and2_1
XFILLER_0_154_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18555_ net295 _09098_ _09122_ _09126_ VGND VGND VPWR VPWR _00004_ sky130_fd_sc_hd__o211a_1
X_12979_ _03071_ VGND VGND VPWR VPWR _03072_ sky130_fd_sc_hd__clkbuf_4
X_15767_ _02992_ _03071_ _06037_ _06041_ VGND VGND VPWR VPWR _06100_ sky130_fd_sc_hd__a31o_1
XFILLER_0_75_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17506_ _07987_ _07988_ VGND VGND VPWR VPWR _07989_ sky130_fd_sc_hd__nor2_1
X_14718_ _04957_ _04958_ _03538_ VGND VGND VPWR VPWR _04959_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18486_ _03155_ _08428_ _03011_ VGND VGND VPWR VPWR _09053_ sky130_fd_sc_hd__or3b_1
XTAP_2790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15698_ _03012_ _09059_ _00322_ _03010_ VGND VGND VPWR VPWR _06025_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_59_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17437_ _07911_ VGND VGND VPWR VPWR _07914_ sky130_fd_sc_hd__inv_2
X_14649_ _04880_ _04881_ net196 _04756_ VGND VGND VPWR VPWR _04883_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_28_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_16 _01115_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_27 _01115_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_38 _01697_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_49 _03265_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17368_ _07836_ _07837_ VGND VGND VPWR VPWR _07838_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_12_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16319_ _02489_ _03152_ _06487_ _06485_ VGND VGND VPWR VPWR _06697_ sky130_fd_sc_hd__or4_1
XFILLER_0_125_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17299_ _07739_ _07740_ _07761_ VGND VGND VPWR VPWR _07763_ sky130_fd_sc_hd__nor3_1
XFILLER_0_3_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput101 net101 VGND VGND VPWR VPWR o_wb_data[26] sky130_fd_sc_hd__clkbuf_4
Xoutput112 net112 VGND VGND VPWR VPWR o_wb_data[7] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09624_ _05366_ _05322_ _05388_ _05410_ VGND VGND VPWR VPWR _05421_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_418 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09555_ _04646_ _04373_ _04395_ _04657_ VGND VGND VPWR VPWR _04668_ sky130_fd_sc_hd__and4_4
XFILLER_0_78_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09486_ _03826_ VGND VGND VPWR VPWR _03914_ sky130_fd_sc_hd__buf_6
XFILLER_0_93_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_136_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_135_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10330_ net338 _00377_ _09346_ _00274_ VGND VGND VPWR VPWR _00423_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_103_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10261_ cla_inst.in2\[31\] _07613_ _00351_ _00352_ VGND VGND VPWR VPWR _00354_ sky130_fd_sc_hd__a22oi_1
X_12000_ _05224_ _00178_ VGND VGND VPWR VPWR _02093_ sky130_fd_sc_hd__nand2_2
X_10192_ _03990_ _05497_ VGND VGND VPWR VPWR _00285_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13951_ _04107_ _04108_ _04119_ VGND VGND VPWR VPWR _04120_ sky130_fd_sc_hd__o21ai_2
X_12902_ _02992_ _01417_ _01359_ _02994_ VGND VGND VPWR VPWR _02995_ sky130_fd_sc_hd__or4_1
X_13882_ _03828_ _04007_ _04043_ _04044_ VGND VGND VPWR VPWR _04046_ sky130_fd_sc_hd__a211oi_2
X_16670_ _06341_ _06546_ _07077_ _00881_ VGND VGND VPWR VPWR _07078_ sky130_fd_sc_hd__a22o_1
X_12833_ _02923_ _02907_ _02924_ _02925_ VGND VGND VPWR VPWR _02926_ sky130_fd_sc_hd__o211ai_4
X_15621_ _05841_ _05940_ VGND VGND VPWR VPWR _05942_ sky130_fd_sc_hd__or2_1
XTAP_2020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18340_ _06374_ _06368_ VGND VGND VPWR VPWR _08895_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15552_ _05866_ VGND VGND VPWR VPWR _05868_ sky130_fd_sc_hd__inv_2
XTAP_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12764_ _01238_ _01272_ _01271_ VGND VGND VPWR VPWR _02857_ sky130_fd_sc_hd__o21ai_1
XTAP_2075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14503_ _04719_ _04720_ _04721_ VGND VGND VPWR VPWR _04724_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_68_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11715_ _01507_ _01806_ _01807_ VGND VGND VPWR VPWR _01808_ sky130_fd_sc_hd__and3_1
XFILLER_0_56_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15483_ _05792_ VGND VGND VPWR VPWR _05793_ sky130_fd_sc_hd__inv_2
X_18271_ _05557_ _06400_ _06401_ VGND VGND VPWR VPWR _08821_ sky130_fd_sc_hd__and3_1
XTAP_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12695_ _02755_ _02785_ VGND VGND VPWR VPWR _02788_ sky130_fd_sc_hd__or2_1
XTAP_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17222_ _04725_ _06510_ _02127_ VGND VGND VPWR VPWR _07680_ sky130_fd_sc_hd__a21o_1
XFILLER_0_154_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14434_ _04645_ _04648_ VGND VGND VPWR VPWR _04649_ sky130_fd_sc_hd__xor2_4
X_11646_ _01721_ _01737_ _01738_ VGND VGND VPWR VPWR _01739_ sky130_fd_sc_hd__nand3_4
XFILLER_0_140_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput14 i_wb_addr[20] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__clkbuf_1
Xinput25 i_wb_addr[30] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_154_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_223 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14365_ _04567_ net181 _04571_ _04572_ VGND VGND VPWR VPWR _04573_ sky130_fd_sc_hd__o211ai_4
X_17153_ _07396_ VGND VGND VPWR VPWR _07604_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_141_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput36 i_wb_data[10] VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__buf_2
X_11577_ _01655_ _01668_ VGND VGND VPWR VPWR _01670_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_25_768 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_107_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_228 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput47 i_wb_data[20] VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__clkbuf_2
X_13316_ _03411_ _03424_ _03425_ VGND VGND VPWR VPWR _03426_ sky130_fd_sc_hd__and3_2
Xinput58 i_wb_data[30] VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__buf_1
XFILLER_0_80_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16104_ _06462_ VGND VGND VPWR VPWR _06463_ sky130_fd_sc_hd__buf_4
Xinput69 reset VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__buf_4
X_10528_ _00617_ _00618_ _00619_ VGND VGND VPWR VPWR _00621_ sky130_fd_sc_hd__a21oi_2
X_17084_ _07518_ _07528_ VGND VGND VPWR VPWR _07529_ sky130_fd_sc_hd__xnor2_1
X_14296_ _01504_ _05856_ VGND VGND VPWR VPWR _04498_ sky130_fd_sc_hd__nand2_1
XFILLER_0_149_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13247_ _03349_ _03350_ VGND VGND VPWR VPWR _03351_ sky130_fd_sc_hd__and2_1
XFILLER_0_0_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16035_ _02985_ _01695_ VGND VGND VPWR VPWR _06388_ sky130_fd_sc_hd__nand2_1
X_10459_ _00544_ _00551_ VGND VGND VPWR VPWR _00552_ sky130_fd_sc_hd__xor2_1
XFILLER_0_110_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13178_ _03269_ _03275_ VGND VGND VPWR VPWR _03277_ sky130_fd_sc_hd__nand2_1
X_12129_ _02185_ _02186_ VGND VGND VPWR VPWR _02222_ sky130_fd_sc_hd__or2_1
X_17986_ _03000_ _06511_ _00813_ VGND VGND VPWR VPWR _08512_ sky130_fd_sc_hd__a21o_1
XFILLER_0_74_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16937_ _06360_ _06545_ _07368_ _03101_ VGND VGND VPWR VPWR _07369_ sky130_fd_sc_hd__a22o_1
X_16868_ _06657_ _07108_ VGND VGND VPWR VPWR _07293_ sky130_fd_sc_hd__nand2_1
X_18607_ _09127_ VGND VGND VPWR VPWR _09163_ sky130_fd_sc_hd__clkbuf_4
X_15819_ _06155_ VGND VGND VPWR VPWR _06156_ sky130_fd_sc_hd__inv_2
X_16799_ _03324_ _06529_ _06814_ _02099_ VGND VGND VPWR VPWR _07218_ sky130_fd_sc_hd__a211o_2
XFILLER_0_90_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_816 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18538_ _09099_ _09100_ _09102_ _09107_ VGND VGND VPWR VPWR _09108_ sky130_fd_sc_hd__nor4_2
XFILLER_0_74_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18469_ _07256_ _09022_ _09025_ _09034_ VGND VGND VPWR VPWR _09035_ sky130_fd_sc_hd__a211o_1
XFILLER_0_63_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_126_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_226 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09607_ _05224_ VGND VGND VPWR VPWR _05235_ sky130_fd_sc_hd__buf_4
X_09538_ _04471_ VGND VGND VPWR VPWR _04482_ sky130_fd_sc_hd__buf_12
XFILLER_0_78_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09469_ _03717_ VGND VGND VPWR VPWR _03728_ sky130_fd_sc_hd__buf_4
XFILLER_0_149_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11500_ _01589_ _01592_ VGND VGND VPWR VPWR _01593_ sky130_fd_sc_hd__and2_1
XFILLER_0_65_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12480_ _02572_ VGND VGND VPWR VPWR _02573_ sky130_fd_sc_hd__inv_2
XFILLER_0_93_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_718 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11431_ _01518_ _01523_ VGND VGND VPWR VPWR _01524_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_136_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14150_ _04181_ _04180_ VGND VGND VPWR VPWR _04338_ sky130_fd_sc_hd__or2b_1
X_11362_ _01401_ _01403_ VGND VGND VPWR VPWR _01455_ sky130_fd_sc_hd__or2b_1
X_13101_ _03165_ _03193_ _02975_ VGND VGND VPWR VPWR _03194_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10313_ _00183_ _03432_ _03618_ _00184_ VGND VGND VPWR VPWR _00406_ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14081_ _03568_ _03571_ _03099_ VGND VGND VPWR VPWR _04262_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11293_ _00811_ _00815_ VGND VGND VPWR VPWR _01386_ sky130_fd_sc_hd__xnor2_1
X_13032_ _06765_ _03123_ VGND VGND VPWR VPWR _03124_ sky130_fd_sc_hd__nor2_2
X_10244_ _09080_ _09131_ VGND VGND VPWR VPWR _00337_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17840_ _07035_ _07125_ _07487_ _07593_ VGND VGND VPWR VPWR _08352_ sky130_fd_sc_hd__or4_2
X_10175_ _07919_ _08289_ _00266_ _00267_ VGND VGND VPWR VPWR _00268_ sky130_fd_sc_hd__o211a_2
XFILLER_0_28_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17771_ _08275_ _08276_ VGND VGND VPWR VPWR _08277_ sky130_fd_sc_hd__nor2_1
X_14983_ _07635_ _05888_ _05127_ _05125_ VGND VGND VPWR VPWR _05248_ sky130_fd_sc_hd__a31o_1
X_16722_ _06945_ _07030_ VGND VGND VPWR VPWR _07135_ sky130_fd_sc_hd__or2b_1
X_13934_ _04099_ _04132_ _07962_ _05715_ VGND VGND VPWR VPWR _04102_ sky130_fd_sc_hd__nand4_1
XFILLER_0_88_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16653_ _06939_ _06966_ VGND VGND VPWR VPWR _07060_ sky130_fd_sc_hd__nand2_1
X_13865_ _03864_ _03869_ VGND VGND VPWR VPWR _04027_ sky130_fd_sc_hd__nand2_1
X_15604_ _05915_ _05923_ VGND VGND VPWR VPWR _05924_ sky130_fd_sc_hd__nor2_1
X_12816_ _01468_ _01490_ _02907_ _02908_ VGND VGND VPWR VPWR _02909_ sky130_fd_sc_hd__a211oi_2
X_16584_ _06866_ _06900_ _06902_ VGND VGND VPWR VPWR _06985_ sky130_fd_sc_hd__a21bo_1
X_13796_ _03777_ _03778_ VGND VGND VPWR VPWR _03951_ sky130_fd_sc_hd__or2_1
XFILLER_0_84_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18323_ _02887_ _08877_ VGND VGND VPWR VPWR _08878_ sky130_fd_sc_hd__or2_1
XFILLER_0_139_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15535_ _03009_ _07668_ _01317_ _05758_ VGND VGND VPWR VPWR _05849_ sky130_fd_sc_hd__and4_1
XTAP_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12747_ _02746_ _02750_ VGND VGND VPWR VPWR _02840_ sky130_fd_sc_hd__or2b_1
XFILLER_0_45_819 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18254_ _08798_ _08801_ VGND VGND VPWR VPWR _08803_ sky130_fd_sc_hd__or2_1
XFILLER_0_154_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15466_ _05757_ _05759_ _05773_ VGND VGND VPWR VPWR _05774_ sky130_fd_sc_hd__a21oi_1
X_12678_ _02762_ _02770_ VGND VGND VPWR VPWR _02771_ sky130_fd_sc_hd__nor2_1
XFILLER_0_38_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_142_504 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17205_ _07648_ _07660_ VGND VGND VPWR VPWR _07661_ sky130_fd_sc_hd__xnor2_1
X_11629_ _01215_ _01209_ _01214_ VGND VGND VPWR VPWR _01722_ sky130_fd_sc_hd__nand3_2
X_14417_ _00877_ _03044_ VGND VGND VPWR VPWR _04630_ sky130_fd_sc_hd__nand2_2
XFILLER_0_115_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18185_ _08632_ _08649_ _08633_ VGND VGND VPWR VPWR _08728_ sky130_fd_sc_hd__o21ba_1
X_15397_ _05697_ _05698_ VGND VGND VPWR VPWR _05699_ sky130_fd_sc_hd__nor2_1
XFILLER_0_13_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17136_ _07561_ _07564_ _07585_ _06723_ _02259_ VGND VGND VPWR VPWR _09389_ sky130_fd_sc_hd__o32a_2
XFILLER_0_52_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14348_ _04552_ _04554_ _03202_ VGND VGND VPWR VPWR _04555_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_40_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14279_ _03014_ _00716_ _04476_ _04478_ VGND VGND VPWR VPWR _04479_ sky130_fd_sc_hd__a22oi_1
X_17067_ _07401_ _07403_ VGND VGND VPWR VPWR _07510_ sky130_fd_sc_hd__nand2_1
XFILLER_0_110_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16018_ _04725_ _06368_ VGND VGND VPWR VPWR _06369_ sky130_fd_sc_hd__or2_1
XTAP_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17969_ _08486_ _08492_ VGND VGND VPWR VPWR _08493_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_109_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_218 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_125_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_721 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_120_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11980_ _02067_ _02070_ net130 _02072_ VGND VGND VPWR VPWR _02073_ sky130_fd_sc_hd__a211oi_4
X_10931_ _04078_ _03771_ _04242_ _00772_ VGND VGND VPWR VPWR _01024_ sky130_fd_sc_hd__and4_1
XFILLER_0_14_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13650_ _06084_ _03455_ _00513_ _03790_ VGND VGND VPWR VPWR _03791_ sky130_fd_sc_hd__a22oi_1
X_10862_ net194 _00953_ _00954_ VGND VGND VPWR VPWR _00955_ sky130_fd_sc_hd__nor3_1
XFILLER_0_14_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12601_ _02650_ net203 VGND VGND VPWR VPWR _02694_ sky130_fd_sc_hd__or2b_1
X_13581_ _03713_ _03714_ _03696_ VGND VGND VPWR VPWR _03716_ sky130_fd_sc_hd__o21ai_1
XPHY_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10793_ _00884_ _00885_ VGND VGND VPWR VPWR _00886_ sky130_fd_sc_hd__nor2_1
XPHY_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15320_ _05516_ _05517_ _05407_ VGND VGND VPWR VPWR _05615_ sky130_fd_sc_hd__and3b_1
X_12532_ _02622_ _02624_ VGND VGND VPWR VPWR _02625_ sky130_fd_sc_hd__xnor2_1
XPHY_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15251_ _07668_ _01223_ _00461_ _03009_ VGND VGND VPWR VPWR _05539_ sky130_fd_sc_hd__a22o_1
X_12463_ _02550_ _02554_ _02555_ VGND VGND VPWR VPWR _02556_ sky130_fd_sc_hd__nand3_1
XFILLER_0_124_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_340 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_124_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14202_ _04188_ _04190_ _04186_ VGND VGND VPWR VPWR _04396_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_50_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11414_ cla_inst.in2\[20\] _01503_ _01240_ _01506_ VGND VGND VPWR VPWR _01507_ sky130_fd_sc_hd__and4_2
X_15182_ _07635_ _00461_ _05334_ _05332_ VGND VGND VPWR VPWR _05465_ sky130_fd_sc_hd__a31o_1
XFILLER_0_105_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12394_ _06019_ _08039_ _09212_ VGND VGND VPWR VPWR _02487_ sky130_fd_sc_hd__and3_1
XFILLER_0_50_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14133_ _00679_ _00678_ _04045_ _04154_ VGND VGND VPWR VPWR _04320_ sky130_fd_sc_hd__and4_1
X_11345_ _01362_ _01437_ VGND VGND VPWR VPWR _01438_ sky130_fd_sc_hd__xnor2_1
X_18941_ clknet_4_2_0_clk _00095_ VGND VGND VPWR VPWR cla_inst.in2\[27\] sky130_fd_sc_hd__dfxtp_2
X_14064_ _03550_ _03552_ _03099_ VGND VGND VPWR VPWR _04245_ sky130_fd_sc_hd__mux2_1
X_11276_ _01337_ _01367_ _01366_ VGND VGND VPWR VPWR _01369_ sky130_fd_sc_hd__o21ai_1
X_13015_ _03107_ VGND VGND VPWR VPWR _03108_ sky130_fd_sc_hd__buf_4
X_10227_ _00318_ _00319_ VGND VGND VPWR VPWR _00320_ sky130_fd_sc_hd__nand2_1
X_18872_ clknet_4_14_0_clk net305 VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__dfxtp_1
X_17823_ _06388_ _06386_ _06387_ VGND VGND VPWR VPWR _08335_ sky130_fd_sc_hd__nand3_1
X_10158_ _00204_ _00214_ _00225_ VGND VGND VPWR VPWR _00251_ sky130_fd_sc_hd__and3_1
XFILLER_0_146_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17754_ _08155_ _08157_ VGND VGND VPWR VPWR _08259_ sky130_fd_sc_hd__and2b_1
X_14966_ _03005_ _05921_ VGND VGND VPWR VPWR _05229_ sky130_fd_sc_hd__nand2_1
XFILLER_0_55_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10089_ _00173_ _00175_ _00178_ _00181_ VGND VGND VPWR VPWR _00182_ sky130_fd_sc_hd__nand4_1
X_16705_ _06653_ _06944_ _07115_ _06571_ VGND VGND VPWR VPWR _07116_ sky130_fd_sc_hd__o22a_1
XFILLER_0_89_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13917_ _04082_ _04083_ _02780_ VGND VGND VPWR VPWR _04084_ sky130_fd_sc_hd__mux2_1
X_17685_ _08063_ _08149_ _08182_ VGND VGND VPWR VPWR _08184_ sky130_fd_sc_hd__or3b_1
XFILLER_0_77_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14897_ _05143_ _05153_ VGND VGND VPWR VPWR _05154_ sky130_fd_sc_hd__xor2_1
X_16636_ _07037_ _07040_ VGND VGND VPWR VPWR _07041_ sky130_fd_sc_hd__nand2_1
X_13848_ _00702_ _04700_ _08409_ _00195_ VGND VGND VPWR VPWR _04008_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_85_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16567_ _06940_ _06965_ VGND VGND VPWR VPWR _06966_ sky130_fd_sc_hd__xor2_1
X_13779_ _03509_ _08746_ _08049_ _03531_ VGND VGND VPWR VPWR _03932_ sky130_fd_sc_hd__a22o_1
XFILLER_0_84_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_476 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18306_ _08844_ _08858_ VGND VGND VPWR VPWR _08859_ sky130_fd_sc_hd__and2b_1
X_15518_ _05828_ _05829_ VGND VGND VPWR VPWR _05830_ sky130_fd_sc_hd__nor2_1
XFILLER_0_29_189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16498_ _06890_ VGND VGND VPWR VPWR _06891_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_38_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18237_ _08707_ _08710_ _08783_ VGND VGND VPWR VPWR _08784_ sky130_fd_sc_hd__nand3_1
X_15449_ _05739_ _05754_ VGND VGND VPWR VPWR _05755_ sky130_fd_sc_hd__and2_1
Xclkbuf_4_4_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_4_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_154_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_811 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_362 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18168_ _08704_ _08708_ VGND VGND VPWR VPWR _08709_ sky130_fd_sc_hd__or2_1
XFILLER_0_52_170 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17119_ _07462_ _07463_ _07460_ VGND VGND VPWR VPWR _07567_ sky130_fd_sc_hd__o21bai_2
Xmax_cap122 _02521_ VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_cap144 _01178_ VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__buf_1
X_18099_ _08632_ _08633_ VGND VGND VPWR VPWR _08634_ sky130_fd_sc_hd__or2_1
XFILLER_0_40_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09941_ _05736_ VGND VGND VPWR VPWR _08865_ sky130_fd_sc_hd__buf_4
XFILLER_0_110_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09872_ _08017_ _08093_ _08104_ VGND VGND VPWR VPWR _08115_ sky130_fd_sc_hd__a21o_1
XTAP_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_137_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_118_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11130_ _06094_ VGND VGND VPWR VPWR _01223_ sky130_fd_sc_hd__buf_4
XFILLER_0_102_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11061_ _01152_ _01153_ VGND VGND VPWR VPWR _01154_ sky130_fd_sc_hd__and2b_1
X_10012_ _09351_ _09353_ _07646_ _09354_ VGND VGND VPWR VPWR _00105_ sky130_fd_sc_hd__and4_1
X_14820_ _05067_ _05068_ _04932_ _04964_ VGND VGND VPWR VPWR _05070_ sky130_fd_sc_hd__a211o_2
XFILLER_0_99_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_98_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14751_ _04856_ _04855_ VGND VGND VPWR VPWR _04994_ sky130_fd_sc_hd__nand2_1
X_11963_ _01941_ _02055_ VGND VGND VPWR VPWR _02056_ sky130_fd_sc_hd__nand2_1
X_13702_ _03845_ _03846_ VGND VGND VPWR VPWR _03849_ sky130_fd_sc_hd__nand2_1
X_10914_ _01004_ _01006_ VGND VGND VPWR VPWR _01007_ sky130_fd_sc_hd__xor2_1
XFILLER_0_86_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17470_ _07947_ _07948_ VGND VGND VPWR VPWR _07949_ sky130_fd_sc_hd__or2_1
X_14682_ _04903_ _04791_ _04917_ _04918_ VGND VGND VPWR VPWR _04920_ sky130_fd_sc_hd__a211o_1
XFILLER_0_86_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11894_ _01980_ _01984_ _01986_ VGND VGND VPWR VPWR _01987_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_67_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16421_ _06802_ _06806_ _03535_ VGND VGND VPWR VPWR _06807_ sky130_fd_sc_hd__a21oi_2
X_13633_ _03768_ _03769_ _03770_ VGND VGND VPWR VPWR _03773_ sky130_fd_sc_hd__a21oi_2
X_10845_ _00932_ _00933_ _00937_ VGND VGND VPWR VPWR _00938_ sky130_fd_sc_hd__a21o_1
XFILLER_0_128_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsplit74 _06560_ VGND VGND VPWR VPWR net237 sky130_fd_sc_hd__dlymetal6s2s_1
X_16352_ _06729_ _06731_ _03098_ VGND VGND VPWR VPWR _06733_ sky130_fd_sc_hd__mux2_1
X_13564_ _03494_ _03505_ VGND VGND VPWR VPWR _03698_ sky130_fd_sc_hd__nand2_1
X_10776_ _00253_ _00194_ _00198_ _00199_ VGND VGND VPWR VPWR _00869_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_81_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15303_ _05593_ _05594_ _05478_ _05553_ VGND VGND VPWR VPWR _05597_ sky130_fd_sc_hd__o211a_1
XFILLER_0_82_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_243 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12515_ ApproximateM_inst.lob_16.lob2.genblk1\[1\].genblk1.mux.sel _00218_ _02607_
+ VGND VGND VPWR VPWR _02608_ sky130_fd_sc_hd__and3_1
X_13495_ _03393_ net134 _03620_ _03621_ VGND VGND VPWR VPWR _03622_ sky130_fd_sc_hd__o211ai_4
X_16283_ _06572_ _06581_ _06657_ _06527_ VGND VGND VPWR VPWR _06658_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_136_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18022_ _07396_ _07780_ _07623_ _07394_ VGND VGND VPWR VPWR _08551_ sky130_fd_sc_hd__a22o_1
X_15234_ _05518_ _05521_ _03930_ VGND VGND VPWR VPWR _05522_ sky130_fd_sc_hd__o21ai_1
X_12446_ _02475_ _02478_ VGND VGND VPWR VPWR _02539_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_23_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15165_ _03008_ _07515_ _00460_ _05856_ VGND VGND VPWR VPWR _05446_ sky130_fd_sc_hd__and4_1
XFILLER_0_23_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12377_ _02176_ _02469_ VGND VGND VPWR VPWR _02470_ sky130_fd_sc_hd__and2_4
XFILLER_0_140_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14116_ _04137_ _04136_ VGND VGND VPWR VPWR _04301_ sky130_fd_sc_hd__and2b_1
X_11328_ _01358_ _01420_ VGND VGND VPWR VPWR _01421_ sky130_fd_sc_hd__xor2_1
X_15096_ _05369_ _05370_ VGND VGND VPWR VPWR _05371_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18924_ clknet_4_11_0_clk _00078_ VGND VGND VPWR VPWR ApproximateM_inst.lob_16.lob2.genblk1\[10\].genblk1.mux.sel
+ sky130_fd_sc_hd__dfxtp_2
X_14047_ _04222_ _04223_ _04224_ VGND VGND VPWR VPWR _04226_ sky130_fd_sc_hd__o21ai_1
X_11259_ _01350_ _01339_ _01340_ VGND VGND VPWR VPWR _01352_ sky130_fd_sc_hd__nor3_1
X_18855_ clknet_4_7_0_clk net276 VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__dfxtp_1
X_17806_ _08314_ _08315_ VGND VGND VPWR VPWR _08316_ sky130_fd_sc_hd__and2_1
X_18786_ _09125_ VGND VGND VPWR VPWR _09298_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_89_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15998_ _06343_ _06344_ _06345_ _06346_ VGND VGND VPWR VPWR _06347_ sky130_fd_sc_hd__and4_1
X_17737_ _02987_ _06920_ _06921_ VGND VGND VPWR VPWR _08241_ sky130_fd_sc_hd__a21o_1
X_14949_ _02989_ _03456_ VGND VGND VPWR VPWR _05210_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17668_ _08159_ _08164_ VGND VGND VPWR VPWR _08165_ sky130_fd_sc_hd__and2_1
XFILLER_0_58_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16619_ _06567_ _06570_ _06946_ _00357_ VGND VGND VPWR VPWR _07022_ sky130_fd_sc_hd__o211a_1
X_17599_ _08088_ _08089_ VGND VGND VPWR VPWR _08090_ sky130_fd_sc_hd__nand2_1
XFILLER_0_9_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09924_ _06373_ _08322_ _08659_ _08670_ VGND VGND VPWR VPWR _08681_ sky130_fd_sc_hd__a211o_2
XFILLER_0_0_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09855_ _07908_ _07897_ _06960_ _05812_ VGND VGND VPWR VPWR _07930_ sky130_fd_sc_hd__a211oi_2
XTAP_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09786_ _06993_ _07025_ _07145_ _07167_ VGND VGND VPWR VPWR _07178_ sky130_fd_sc_hd__nand4_2
XTAP_2405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_106 op_code\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_117 _00166_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_128 _04034_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_139 _06765_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10630_ _00512_ _00518_ VGND VGND VPWR VPWR _00723_ sky130_fd_sc_hd__or2_1
XFILLER_0_48_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_119_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10561_ _00651_ _00652_ _00643_ VGND VGND VPWR VPWR _00654_ sky130_fd_sc_hd__a21o_1
XFILLER_0_146_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12300_ _02258_ _02260_ _02386_ VGND VGND VPWR VPWR _02393_ sky130_fd_sc_hd__or3_1
XFILLER_0_118_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13280_ _00459_ _03384_ _03385_ VGND VGND VPWR VPWR _03386_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_63_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10492_ net339 _00424_ _00583_ _00584_ VGND VGND VPWR VPWR _00585_ sky130_fd_sc_hd__o211a_4
XFILLER_0_134_676 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12231_ _02313_ _02318_ _02317_ VGND VGND VPWR VPWR _02324_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_122_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12162_ _02240_ _02253_ VGND VGND VPWR VPWR _02255_ sky130_fd_sc_hd__nand2_1
XFILLER_0_20_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11113_ _07047_ _07254_ _05497_ _04580_ VGND VGND VPWR VPWR _01206_ sky130_fd_sc_hd__nand4_2
XFILLER_0_130_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12093_ _02177_ _02182_ VGND VGND VPWR VPWR _02186_ sky130_fd_sc_hd__xor2_1
X_16970_ _07401_ _07403_ VGND VGND VPWR VPWR _07404_ sky130_fd_sc_hd__xor2_1
X_11044_ _01105_ _00514_ _01136_ _00813_ VGND VGND VPWR VPWR _01137_ sky130_fd_sc_hd__or4_4
X_15921_ _04955_ _04957_ _03536_ VGND VGND VPWR VPWR _06266_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18640_ _09176_ _09186_ VGND VGND VPWR VPWR _09187_ sky130_fd_sc_hd__and2_1
X_15852_ _06183_ _06187_ _06190_ VGND VGND VPWR VPWR _06192_ sky130_fd_sc_hd__o21ai_1
X_14803_ _05036_ _05037_ _05049_ VGND VGND VPWR VPWR _05052_ sky130_fd_sc_hd__nand3_1
X_18571_ net273 _09098_ _09136_ _09126_ VGND VGND VPWR VPWR _00011_ sky130_fd_sc_hd__o211a_1
X_15783_ _06098_ _06099_ _06117_ VGND VGND VPWR VPWR _06118_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_59_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12995_ _03023_ _03087_ VGND VGND VPWR VPWR _03088_ sky130_fd_sc_hd__nand2_1
X_17522_ _08004_ _08005_ VGND VGND VPWR VPWR _08007_ sky130_fd_sc_hd__nor2_1
XFILLER_0_86_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14734_ _04972_ _04974_ _04838_ _04839_ VGND VGND VPWR VPWR _04976_ sky130_fd_sc_hd__o211ai_2
X_11946_ _02035_ _02038_ VGND VGND VPWR VPWR _02039_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_59_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17453_ _07891_ _07892_ _07895_ VGND VGND VPWR VPWR _07931_ sky130_fd_sc_hd__and3_1
X_14665_ _00164_ _04900_ VGND VGND VPWR VPWR _04901_ sky130_fd_sc_hd__nand2_2
X_11877_ _01865_ _01867_ _01868_ _01861_ VGND VGND VPWR VPWR _01970_ sky130_fd_sc_hd__o31ai_2
X_16404_ _06544_ VGND VGND VPWR VPWR _06790_ sky130_fd_sc_hd__clkbuf_4
X_13616_ _03588_ _03589_ _03590_ VGND VGND VPWR VPWR _03754_ sky130_fd_sc_hd__nor3_2
X_17384_ _07726_ _07720_ VGND VGND VPWR VPWR _07856_ sky130_fd_sc_hd__and2b_1
X_10828_ _03771_ ApproximateM_inst.lob_16.lob1.genblk1\[8\].genblk1.mux.sel _04220_
+ cla_inst.in2\[16\] VGND VGND VPWR VPWR _00921_ sky130_fd_sc_hd__a22o_1
X_14596_ _02979_ _03551_ _04825_ VGND VGND VPWR VPWR _04826_ sky130_fd_sc_hd__o21a_1
XFILLER_0_144_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_744 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_116_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16335_ _03050_ _02563_ _03173_ _06470_ _06714_ VGND VGND VPWR VPWR _06715_ sky130_fd_sc_hd__o311a_1
X_13547_ cla_inst.in2\[24\] _00174_ _04886_ _03903_ VGND VGND VPWR VPWR _03679_ sky130_fd_sc_hd__and4_1
X_10759_ _00829_ _00851_ VGND VGND VPWR VPWR _00852_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_42_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16266_ _00167_ _03101_ _00593_ _00558_ _03028_ _02982_ VGND VGND VPWR VPWR _06640_
+ sky130_fd_sc_hd__mux4_1
X_13478_ _03595_ _03597_ _03602_ VGND VGND VPWR VPWR _03603_ sky130_fd_sc_hd__nand3_1
XFILLER_0_112_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18005_ _07039_ _07708_ _08460_ _08357_ VGND VGND VPWR VPWR _08532_ sky130_fd_sc_hd__a31o_1
X_15217_ _05429_ _05390_ _05502_ VGND VGND VPWR VPWR _05503_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_140_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12429_ _02450_ _02455_ _02454_ VGND VGND VPWR VPWR _02522_ sky130_fd_sc_hd__o21ai_1
X_16197_ _03281_ _06529_ _06520_ VGND VGND VPWR VPWR _06564_ sky130_fd_sc_hd__a21o_1
XFILLER_0_124_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15148_ _05402_ _05403_ VGND VGND VPWR VPWR _05427_ sky130_fd_sc_hd__and2b_1
XFILLER_0_50_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15079_ _09350_ _05964_ _06094_ _00112_ VGND VGND VPWR VPWR _05352_ sky130_fd_sc_hd__a22oi_1
X_18907_ clknet_4_10_0_clk _00061_ VGND VGND VPWR VPWR cla_inst.in1\[25\] sky130_fd_sc_hd__dfxtp_1
X_09640_ _05584_ VGND VGND VPWR VPWR _05595_ sky130_fd_sc_hd__clkbuf_4
X_18838_ clknet_4_0_0_clk net296 VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09571_ _04810_ _04821_ _04831_ VGND VGND VPWR VPWR _04842_ sky130_fd_sc_hd__nand3_1
X_18769_ _09273_ _09284_ VGND VGND VPWR VPWR _09285_ sky130_fd_sc_hd__and2_1
XFILLER_0_148_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_418 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09907_ _08398_ _08474_ _08485_ VGND VGND VPWR VPWR _08496_ sky130_fd_sc_hd__nand3_1
X_09838_ _07733_ VGND VGND VPWR VPWR _07744_ sky130_fd_sc_hd__buf_4
XTAP_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09769_ _06982_ VGND VGND VPWR VPWR _06993_ sky130_fd_sc_hd__clkbuf_8
XTAP_2202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11800_ _01872_ _01875_ VGND VGND VPWR VPWR _01893_ sky130_fd_sc_hd__xnor2_1
XTAP_2224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12780_ _00591_ _01264_ _01263_ _01261_ VGND VGND VPWR VPWR _02873_ sky130_fd_sc_hd__a31o_2
XTAP_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer70 _00694_ VGND VGND VPWR VPWR net327 sky130_fd_sc_hd__dlymetal6s4s_1
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xrebuffer81 net243 VGND VGND VPWR VPWR net244 sky130_fd_sc_hd__clkbuf_1
XTAP_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer92 _00378_ VGND VGND VPWR VPWR net339 sky130_fd_sc_hd__dlygate4sd1_1
XTAP_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11731_ _01821_ _01822_ _01823_ VGND VGND VPWR VPWR _01824_ sky130_fd_sc_hd__o21ba_1
XTAP_2279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14450_ _04664_ _04665_ VGND VGND VPWR VPWR _04666_ sky130_fd_sc_hd__nand2_1
XTAP_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11662_ _01739_ _01740_ _01642_ net125 VGND VGND VPWR VPWR _01755_ sky130_fd_sc_hd__a211o_1
XFILLER_0_37_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13401_ _03516_ _03517_ _03371_ _03372_ VGND VGND VPWR VPWR _03519_ sky130_fd_sc_hd__a211oi_2
X_10613_ _00253_ _00398_ VGND VGND VPWR VPWR _00706_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14381_ _04515_ _04588_ _04589_ VGND VGND VPWR VPWR _04590_ sky130_fd_sc_hd__a21bo_1
X_11593_ _01208_ _01683_ _01682_ VGND VGND VPWR VPWR _01686_ sky130_fd_sc_hd__a21o_1
X_16120_ _03164_ _06476_ _06479_ _03547_ VGND VGND VPWR VPWR _06480_ sky130_fd_sc_hd__o211a_1
XFILLER_0_36_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13332_ _03440_ VGND VGND VPWR VPWR _03444_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10544_ _00476_ _00480_ VGND VGND VPWR VPWR _00637_ sky130_fd_sc_hd__and2_1
XFILLER_0_106_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_107_676 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_122_602 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16051_ _02992_ _03068_ VGND VGND VPWR VPWR _06405_ sky130_fd_sc_hd__or2_1
X_10475_ _00566_ _00567_ VGND VGND VPWR VPWR _00568_ sky130_fd_sc_hd__xnor2_1
X_13263_ _00592_ VGND VGND VPWR VPWR _03368_ sky130_fd_sc_hd__buf_4
XFILLER_0_51_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15002_ _01504_ _08876_ VGND VGND VPWR VPWR _05269_ sky130_fd_sc_hd__nand2_1
X_12214_ _02302_ _02305_ _02304_ VGND VGND VPWR VPWR _02307_ sky130_fd_sc_hd__o21ai_1
X_13194_ _00661_ net327 _03293_ _03294_ VGND VGND VPWR VPWR _03295_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_121_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12145_ _02236_ _02237_ VGND VGND VPWR VPWR _02238_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_20_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12076_ _02168_ _01991_ VGND VGND VPWR VPWR _02169_ sky130_fd_sc_hd__xnor2_1
X_16953_ _06460_ VGND VGND VPWR VPWR _07386_ sky130_fd_sc_hd__inv_2
X_11027_ _01118_ _01119_ VGND VGND VPWR VPWR _01120_ sky130_fd_sc_hd__nor2_1
X_15904_ _06247_ VGND VGND VPWR VPWR _06248_ sky130_fd_sc_hd__buf_2
X_16884_ _01962_ _06812_ _06871_ VGND VGND VPWR VPWR _07311_ sky130_fd_sc_hd__o21ai_4
X_18623_ net308 _09157_ _09173_ _09162_ VGND VGND VPWR VPWR _00032_ sky130_fd_sc_hd__o211a_1
XFILLER_0_154_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15835_ _06118_ _06173_ VGND VGND VPWR VPWR _06174_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_99_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18554_ _09125_ VGND VGND VPWR VPWR _09126_ sky130_fd_sc_hd__buf_2
X_15766_ _06047_ _06046_ VGND VGND VPWR VPWR _06099_ sky130_fd_sc_hd__and2b_1
X_12978_ _00495_ VGND VGND VPWR VPWR _03071_ sky130_fd_sc_hd__clkbuf_4
X_17505_ _07985_ _07986_ VGND VGND VPWR VPWR _07988_ sky130_fd_sc_hd__nor2_1
X_14717_ _03547_ _03572_ VGND VGND VPWR VPWR _04958_ sky130_fd_sc_hd__or2_1
XFILLER_0_59_368 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18485_ _03011_ _06512_ _03155_ VGND VGND VPWR VPWR _09052_ sky130_fd_sc_hd__a21bo_1
X_11929_ _02007_ _02008_ VGND VGND VPWR VPWR _02022_ sky130_fd_sc_hd__xor2_1
XTAP_2780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15697_ _03015_ _00339_ VGND VGND VPWR VPWR _06024_ sky130_fd_sc_hd__and2_2
XTAP_2791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_891 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17436_ _07910_ _07911_ _07912_ VGND VGND VPWR VPWR _07913_ sky130_fd_sc_hd__and3b_1
XFILLER_0_137_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14648_ _04741_ _04756_ _04880_ _04881_ VGND VGND VPWR VPWR _04882_ sky130_fd_sc_hd__a211o_1
XFILLER_0_145_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_17 _01115_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_28 _01115_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_39 _01697_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17367_ _07018_ _07387_ VGND VGND VPWR VPWR _07837_ sky130_fd_sc_hd__nor2_1
X_14579_ _04805_ _04806_ VGND VGND VPWR VPWR _04807_ sky130_fd_sc_hd__nor2_2
XFILLER_0_28_799 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_75 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16318_ _02982_ _06490_ _06695_ _06626_ VGND VGND VPWR VPWR _06696_ sky130_fd_sc_hd__o211a_1
XFILLER_0_82_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17298_ _07739_ _07740_ _07761_ VGND VGND VPWR VPWR _07762_ sky130_fd_sc_hd__o21a_1
XFILLER_0_31_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16249_ _06470_ _06620_ VGND VGND VPWR VPWR _06621_ sky130_fd_sc_hd__nand2_1
Xoutput102 net102 VGND VGND VPWR VPWR o_wb_data[27] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_51_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput113 net113 VGND VGND VPWR VPWR o_wb_data[8] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_101_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09623_ _05399_ VGND VGND VPWR VPWR _05410_ sky130_fd_sc_hd__buf_4
X_09554_ _03739_ VGND VGND VPWR VPWR _04657_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_77_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09485_ ApproximateM_inst.lob_16.lob1.genblk1\[12\].genblk1.mux.sel VGND VGND VPWR
+ VPWR _03903_ sky130_fd_sc_hd__buf_4
XFILLER_0_66_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_755 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_135_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_143_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_104_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10260_ cla_inst.in2\[31\] _07613_ _00351_ _00352_ VGND VGND VPWR VPWR _00353_ sky130_fd_sc_hd__and4_1
XFILLER_0_103_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10191_ _00282_ _00283_ VGND VGND VPWR VPWR _00284_ sky130_fd_sc_hd__nor2_1
X_13950_ _04117_ _04118_ VGND VGND VPWR VPWR _04119_ sky130_fd_sc_hd__or2_1
X_12901_ _02993_ VGND VGND VPWR VPWR _02994_ sky130_fd_sc_hd__buf_2
X_13881_ _04041_ _04042_ _04024_ VGND VGND VPWR VPWR _04044_ sky130_fd_sc_hd__o21a_1
XFILLER_0_88_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15620_ _05841_ _05940_ VGND VGND VPWR VPWR _05941_ sky130_fd_sc_hd__nand2_1
XTAP_2010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12832_ _00856_ _00890_ _00889_ VGND VGND VPWR VPWR _02925_ sky130_fd_sc_hd__o21ai_2
XTAP_2021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15551_ _05776_ _05778_ _05864_ _05865_ VGND VGND VPWR VPWR _05866_ sky130_fd_sc_hd__o211a_1
XTAP_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12763_ _01238_ _01271_ _01272_ VGND VGND VPWR VPWR _02856_ sky130_fd_sc_hd__or3_1
XFILLER_0_56_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14502_ _04719_ _04720_ _04721_ VGND VGND VPWR VPWR _04723_ sky130_fd_sc_hd__and3_2
XTAP_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11714_ _01804_ _01805_ _01784_ _01787_ VGND VGND VPWR VPWR _01807_ sky130_fd_sc_hd__a211o_1
X_18270_ _02881_ _08819_ VGND VGND VPWR VPWR _08820_ sky130_fd_sc_hd__xnor2_4
XTAP_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15482_ _05615_ _05790_ VGND VGND VPWR VPWR _05792_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12694_ _02505_ _00134_ _00108_ _00845_ VGND VGND VPWR VPWR _02787_ sky130_fd_sc_hd__a22o_1
XTAP_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17221_ _02633_ _07676_ _07677_ VGND VGND VPWR VPWR _07678_ sky130_fd_sc_hd__a21oi_2
X_14433_ _01873_ _04647_ VGND VGND VPWR VPWR _04648_ sky130_fd_sc_hd__nand2_2
XFILLER_0_126_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11645_ _01719_ _01720_ _01621_ _01640_ VGND VGND VPWR VPWR _01738_ sky130_fd_sc_hd__a211o_1
XFILLER_0_65_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17152_ _07589_ _07601_ VGND VGND VPWR VPWR _07603_ sky130_fd_sc_hd__xnor2_1
Xinput15 i_wb_addr[21] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__clkbuf_1
X_14364_ _02986_ _06732_ _04568_ _04570_ VGND VGND VPWR VPWR _04572_ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput26 i_wb_addr[31] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11576_ _01655_ _01668_ VGND VGND VPWR VPWR _01669_ sky130_fd_sc_hd__or2_1
Xinput37 i_wb_data[11] VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__buf_2
XFILLER_0_13_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput48 i_wb_data[21] VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__clkbuf_2
X_16103_ _06461_ VGND VGND VPWR VPWR _06462_ sky130_fd_sc_hd__clkbuf_4
X_13315_ _03422_ _03423_ _03416_ VGND VGND VPWR VPWR _03425_ sky130_fd_sc_hd__a21o_1
Xinput59 i_wb_data[31] VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__clkbuf_2
X_10527_ _00617_ _00618_ _00619_ VGND VGND VPWR VPWR _00620_ sky130_fd_sc_hd__and3_4
XFILLER_0_122_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17083_ _07525_ _07527_ VGND VGND VPWR VPWR _07528_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14295_ _04495_ _04496_ VGND VGND VPWR VPWR _04497_ sky130_fd_sc_hd__nor2_1
X_16034_ _02985_ _01695_ VGND VGND VPWR VPWR _06387_ sky130_fd_sc_hd__or2_2
X_13246_ _03347_ _03348_ _00747_ _03203_ VGND VGND VPWR VPWR _03350_ sky130_fd_sc_hd__a211o_1
X_10458_ _00545_ _00550_ VGND VGND VPWR VPWR _00551_ sky130_fd_sc_hd__xor2_1
XFILLER_0_149_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10389_ _00468_ _00469_ _00481_ VGND VGND VPWR VPWR _00482_ sky130_fd_sc_hd__a21o_2
X_13177_ _03269_ _03275_ VGND VGND VPWR VPWR _03276_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12128_ _02218_ _02220_ VGND VGND VPWR VPWR _02221_ sky130_fd_sc_hd__nand2_1
X_17985_ _02167_ _02174_ _08424_ _08510_ _03202_ VGND VGND VPWR VPWR _08511_ sky130_fd_sc_hd__o311a_2
X_16936_ _00644_ _06592_ _06551_ VGND VGND VPWR VPWR _07368_ sky130_fd_sc_hd__a21o_1
X_12059_ _02151_ VGND VGND VPWR VPWR _02152_ sky130_fd_sc_hd__inv_2
X_16867_ _07288_ _07291_ VGND VGND VPWR VPWR _07292_ sky130_fd_sc_hd__xor2_2
X_15818_ _03010_ _03012_ _03071_ _03149_ VGND VGND VPWR VPWR _06155_ sky130_fd_sc_hd__and4_1
X_18606_ net279 _09157_ _09161_ _09162_ VGND VGND VPWR VPWR _00024_ sky130_fd_sc_hd__o211a_1
XFILLER_0_149_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16798_ _07038_ _06969_ _07216_ _06527_ VGND VGND VPWR VPWR _07217_ sky130_fd_sc_hd__a22o_1
X_18537_ _09103_ _09104_ _09105_ _09106_ VGND VGND VPWR VPWR _09107_ sky130_fd_sc_hd__or4_2
X_15749_ _06074_ _06080_ VGND VGND VPWR VPWR _06081_ sky130_fd_sc_hd__or2_1
XFILLER_0_90_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18468_ _06412_ _06421_ _09026_ _09033_ VGND VGND VPWR VPWR _09034_ sky130_fd_sc_hd__a31o_1
XFILLER_0_114_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17419_ _07767_ _07768_ _07770_ VGND VGND VPWR VPWR _07894_ sky130_fd_sc_hd__or3_1
X_18399_ _04406_ _07592_ _08957_ VGND VGND VPWR VPWR _08959_ sky130_fd_sc_hd__a21o_1
XFILLER_0_90_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_736 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_479 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_126_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_452 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09606_ _05213_ VGND VGND VPWR VPWR _05224_ sky130_fd_sc_hd__buf_4
XFILLER_0_78_441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09537_ ApproximateM_inst.lob_16.lob1.genblk1\[14\].genblk1.mux.sel VGND VGND VPWR
+ VPWR _04471_ sky130_fd_sc_hd__buf_6
XFILLER_0_149_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09468_ ApproximateM_inst.lob_16.lob2.genblk1\[14\].genblk1.mux.sel VGND VGND VPWR
+ VPWR _03717_ sky130_fd_sc_hd__buf_4
XFILLER_0_109_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_596 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11430_ _01519_ _01522_ VGND VGND VPWR VPWR _01523_ sky130_fd_sc_hd__nor2_1
XFILLER_0_117_771 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_123_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11361_ _01415_ _01438_ _01439_ VGND VGND VPWR VPWR _01454_ sky130_fd_sc_hd__nor3_1
XFILLER_0_104_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10312_ _00184_ _00183_ _03432_ _00205_ VGND VGND VPWR VPWR _00405_ sky130_fd_sc_hd__and4_1
X_13100_ _03178_ _03192_ _02780_ VGND VGND VPWR VPWR _03193_ sky130_fd_sc_hd__mux2_1
X_11292_ _01281_ _01282_ VGND VGND VPWR VPWR _01385_ sky130_fd_sc_hd__or2b_1
X_14080_ _04247_ _04258_ _04260_ VGND VGND VPWR VPWR _04261_ sky130_fd_sc_hd__o21ai_1
X_10243_ _08681_ _09005_ _00333_ _00335_ VGND VGND VPWR VPWR _00336_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_30_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13031_ _02728_ _02965_ _03239_ _03217_ VGND VGND VPWR VPWR _03123_ sky130_fd_sc_hd__or4b_4
X_10174_ _00245_ _00246_ _00265_ VGND VGND VPWR VPWR _00267_ sky130_fd_sc_hd__nand3_2
X_17770_ _08259_ _08166_ _08274_ VGND VGND VPWR VPWR _08276_ sky130_fd_sc_hd__nor3_1
X_14982_ _05146_ _05149_ VGND VGND VPWR VPWR _05247_ sky130_fd_sc_hd__nand2_1
X_16721_ _07122_ _07132_ VGND VGND VPWR VPWR _07133_ sky130_fd_sc_hd__xnor2_1
X_13933_ _04132_ _07962_ _00308_ _04099_ VGND VGND VPWR VPWR _04101_ sky130_fd_sc_hd__a22o_1
XFILLER_0_89_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16652_ _07049_ _07057_ VGND VGND VPWR VPWR _07059_ sky130_fd_sc_hd__xnor2_1
X_13864_ _03861_ _03873_ VGND VGND VPWR VPWR _04026_ sky130_fd_sc_hd__nand2_1
X_15603_ _05920_ _05922_ VGND VGND VPWR VPWR _05923_ sky130_fd_sc_hd__or2_1
X_12815_ _02899_ _02906_ _02905_ VGND VGND VPWR VPWR _02908_ sky130_fd_sc_hd__a21oi_1
X_16583_ _06981_ _06983_ VGND VGND VPWR VPWR _06984_ sky130_fd_sc_hd__or2b_1
X_13795_ _03945_ _03947_ _03948_ VGND VGND VPWR VPWR _03950_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_84_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18322_ _08875_ _08759_ _02893_ VGND VGND VPWR VPWR _08877_ sky130_fd_sc_hd__o21a_1
XTAP_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15534_ _03006_ _04647_ VGND VGND VPWR VPWR _05848_ sky130_fd_sc_hd__nand2_1
X_12746_ _02837_ _02838_ VGND VGND VPWR VPWR _02839_ sky130_fd_sc_hd__and2_1
XFILLER_0_29_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_362 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18253_ _08798_ _08801_ VGND VGND VPWR VPWR _08802_ sky130_fd_sc_hd__nand2_1
X_15465_ _05771_ _05772_ VGND VGND VPWR VPWR _05773_ sky130_fd_sc_hd__and2_1
XFILLER_0_84_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12677_ _02753_ _02761_ VGND VGND VPWR VPWR _02770_ sky130_fd_sc_hd__and2_1
XFILLER_0_154_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17204_ _07658_ _07659_ VGND VGND VPWR VPWR _07660_ sky130_fd_sc_hd__nor2_1
X_14416_ _04626_ _04627_ _04470_ _04488_ VGND VGND VPWR VPWR _04629_ sky130_fd_sc_hd__o211a_1
XFILLER_0_154_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11628_ _01621_ _01640_ _01719_ _01720_ VGND VGND VPWR VPWR _01721_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_108_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18184_ _08725_ _08726_ VGND VGND VPWR VPWR _08727_ sky130_fd_sc_hd__nor2_1
X_15396_ _05549_ _05598_ _05696_ VGND VGND VPWR VPWR _05698_ sky130_fd_sc_hd__and3_1
XFILLER_0_4_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17135_ _07256_ _07568_ _07569_ _07584_ VGND VGND VPWR VPWR _07585_ sky130_fd_sc_hd__a31o_1
X_14347_ _04401_ _04410_ _04553_ VGND VGND VPWR VPWR _04554_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_107_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_590 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11559_ _01649_ _01650_ _01651_ VGND VGND VPWR VPWR _01652_ sky130_fd_sc_hd__and3_1
XFILLER_0_123_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_150_560 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17066_ _07415_ _07423_ VGND VGND VPWR VPWR _07509_ sky130_fd_sc_hd__nor2_1
X_14278_ _04475_ VGND VGND VPWR VPWR _04478_ sky130_fd_sc_hd__inv_2
XFILLER_0_110_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_150_593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16017_ _00716_ VGND VGND VPWR VPWR _06368_ sky130_fd_sc_hd__clkbuf_4
X_13229_ _03317_ _03331_ VGND VGND VPWR VPWR _03332_ sky130_fd_sc_hd__xnor2_2
XTAP_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17968_ _08490_ _08491_ VGND VGND VPWR VPWR _08492_ sky130_fd_sc_hd__nor2_1
X_16919_ _07347_ _07348_ VGND VGND VPWR VPWR _07349_ sky130_fd_sc_hd__and2_4
X_17899_ _08120_ _08219_ _08414_ _08416_ _08325_ VGND VGND VPWR VPWR _08417_ sky130_fd_sc_hd__o311a_1
XFILLER_0_79_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_146_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_733 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_83 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_555 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_114_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_796 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10930_ _00939_ _00938_ _00931_ VGND VGND VPWR VPWR _01023_ sky130_fd_sc_hd__a21o_1
X_10861_ _00925_ _00926_ _00940_ VGND VGND VPWR VPWR _00954_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_79_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_731 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12600_ _02672_ _02673_ _02692_ VGND VGND VPWR VPWR _02693_ sky130_fd_sc_hd__and3_1
XPHY_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13580_ _03696_ _03713_ _03714_ VGND VGND VPWR VPWR _03715_ sky130_fd_sc_hd__or3_2
XPHY_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10792_ _00883_ _00876_ _00880_ VGND VGND VPWR VPWR _00885_ sky130_fd_sc_hd__nor3_1
XFILLER_0_66_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_904 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12531_ _02567_ _02623_ VGND VGND VPWR VPWR _02624_ sky130_fd_sc_hd__xnor2_1
XPHY_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_820 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_137_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15250_ _03009_ _07668_ _01223_ _00461_ VGND VGND VPWR VPWR _05538_ sky130_fd_sc_hd__and4_1
XFILLER_0_136_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12462_ _02545_ _02549_ _02548_ VGND VGND VPWR VPWR _02555_ sky130_fd_sc_hd__a21o_1
XFILLER_0_35_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_136_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14201_ _04390_ _04391_ _04392_ VGND VGND VPWR VPWR _04394_ sky130_fd_sc_hd__o21a_1
XFILLER_0_151_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11413_ _00877_ _07646_ _09354_ _01505_ VGND VGND VPWR VPWR _01506_ sky130_fd_sc_hd__a22o_1
XFILLER_0_152_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15181_ _05353_ _05354_ VGND VGND VPWR VPWR _05463_ sky130_fd_sc_hd__or2_1
XFILLER_0_35_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12393_ _08039_ _00871_ _07548_ _06019_ VGND VGND VPWR VPWR _02486_ sky130_fd_sc_hd__a22o_1
X_14132_ _03005_ _00166_ VGND VGND VPWR VPWR _04319_ sky130_fd_sc_hd__nand2_1
X_11344_ _01416_ _01436_ VGND VGND VPWR VPWR _01437_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_132_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18940_ clknet_4_2_0_clk _00094_ VGND VGND VPWR VPWR cla_inst.in2\[26\] sky130_fd_sc_hd__dfxtp_2
X_14063_ _02976_ _04241_ _03038_ _04243_ VGND VGND VPWR VPWR _04244_ sky130_fd_sc_hd__or4_1
X_11275_ _01337_ _01366_ _01367_ VGND VGND VPWR VPWR _01368_ sky130_fd_sc_hd__or3_1
XFILLER_0_120_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13014_ _01962_ VGND VGND VPWR VPWR _03107_ sky130_fd_sc_hd__clkbuf_8
X_10226_ _06029_ _05649_ _07112_ VGND VGND VPWR VPWR _00319_ sky130_fd_sc_hd__and3_1
X_18871_ clknet_4_14_0_clk net254 VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__dfxtp_1
X_10157_ _00222_ _00224_ VGND VGND VPWR VPWR _00250_ sky130_fd_sc_hd__and2b_1
X_17822_ _08329_ _08330_ _08331_ VGND VGND VPWR VPWR _08334_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_55_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17753_ _08171_ _08181_ VGND VGND VPWR VPWR _08258_ sky130_fd_sc_hd__nand2_1
X_14965_ _05226_ _05227_ VGND VGND VPWR VPWR _05228_ sky130_fd_sc_hd__and2b_1
X_10088_ _00180_ VGND VGND VPWR VPWR _00181_ sky130_fd_sc_hd__buf_6
XFILLER_0_89_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16704_ net147 _07024_ _03790_ VGND VGND VPWR VPWR _07115_ sky130_fd_sc_hd__o21ai_4
X_13916_ _03138_ _03190_ _00494_ VGND VGND VPWR VPWR _04083_ sky130_fd_sc_hd__mux2_1
X_17684_ _08063_ _08149_ _08182_ VGND VGND VPWR VPWR _08183_ sky130_fd_sc_hd__o21ba_1
X_14896_ _05151_ _05152_ VGND VGND VPWR VPWR _05153_ sky130_fd_sc_hd__nor2_1
X_16635_ _06762_ _07038_ _07039_ _06527_ VGND VGND VPWR VPWR _07040_ sky130_fd_sc_hd__a22o_1
X_13847_ _03830_ _03814_ VGND VGND VPWR VPWR _04007_ sky130_fd_sc_hd__or2b_1
XFILLER_0_58_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16566_ _06941_ _06964_ VGND VGND VPWR VPWR _06965_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_146_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13778_ _03772_ _03773_ _03783_ VGND VGND VPWR VPWR _03931_ sky130_fd_sc_hd__nor3_2
XFILLER_0_85_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15517_ _05809_ _05810_ _05827_ VGND VGND VPWR VPWR _05829_ sky130_fd_sc_hd__nor3_1
X_18305_ _08856_ _08857_ VGND VGND VPWR VPWR _08858_ sky130_fd_sc_hd__nor2_1
XFILLER_0_45_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12729_ _02813_ _02821_ VGND VGND VPWR VPWR _02822_ sky130_fd_sc_hd__nor2_1
XFILLER_0_139_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16497_ _06811_ _06889_ _00193_ VGND VGND VPWR VPWR _06890_ sky130_fd_sc_hd__and3b_1
X_18236_ _08781_ _08782_ VGND VGND VPWR VPWR _08783_ sky130_fd_sc_hd__or2_1
XFILLER_0_44_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15448_ _05752_ _05753_ VGND VGND VPWR VPWR _05754_ sky130_fd_sc_hd__nor2_1
XFILLER_0_128_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18167_ _08705_ _08706_ _08707_ VGND VGND VPWR VPWR _08708_ sky130_fd_sc_hd__and3_1
X_15379_ _05678_ VGND VGND VPWR VPWR _05679_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_823 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_130_508 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17118_ _00558_ _07355_ _02347_ VGND VGND VPWR VPWR _07566_ sky130_fd_sc_hd__or3b_1
XFILLER_0_40_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_cap123 _02389_ VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__buf_1
X_18098_ _08617_ _08618_ _08631_ VGND VGND VPWR VPWR _08633_ sky130_fd_sc_hd__a21oi_1
Xmax_cap134 _03587_ VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__buf_1
XFILLER_0_111_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09940_ _08832_ _08843_ _05682_ _07156_ VGND VGND VPWR VPWR _08854_ sky130_fd_sc_hd__and4b_1
X_17049_ _07113_ net145 _07489_ _06542_ VGND VGND VPWR VPWR _07490_ sky130_fd_sc_hd__a22o_1
XFILLER_0_110_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09871_ _08060_ _08082_ _08028_ _07286_ VGND VGND VPWR VPWR _08104_ sky130_fd_sc_hd__o211a_1
XTAP_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_134_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11060_ _01151_ _00176_ _00145_ _04078_ VGND VGND VPWR VPWR _01153_ sky130_fd_sc_hd__a22o_1
X_10011_ _07657_ VGND VGND VPWR VPWR _09354_ sky130_fd_sc_hd__buf_4
X_14750_ _04989_ _04990_ _04991_ VGND VGND VPWR VPWR _04993_ sky130_fd_sc_hd__a21o_1
X_11962_ _01938_ _01939_ _01940_ VGND VGND VPWR VPWR _02055_ sky130_fd_sc_hd__o21ai_1
X_13701_ _03845_ _03846_ VGND VGND VPWR VPWR _03847_ sky130_fd_sc_hd__or2_1
X_10913_ _05235_ _01005_ _00983_ _00982_ VGND VGND VPWR VPWR _01006_ sky130_fd_sc_hd__a31o_1
X_14681_ _04904_ _04905_ _04916_ VGND VGND VPWR VPWR _04918_ sky130_fd_sc_hd__nor3_1
X_11893_ _01895_ _01985_ VGND VGND VPWR VPWR _01986_ sky130_fd_sc_hd__or2_1
XFILLER_0_129_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16420_ _06803_ _06520_ net150 _06805_ sel_op\[0\] VGND VGND VPWR VPWR _06806_ sky130_fd_sc_hd__a2111o_1
X_13632_ _03768_ _03769_ _03770_ VGND VGND VPWR VPWR _03772_ sky130_fd_sc_hd__and3_1
X_10844_ _00934_ _00935_ _00936_ VGND VGND VPWR VPWR _00937_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_67_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_128_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16351_ _03049_ _06618_ _06730_ _06626_ VGND VGND VPWR VPWR _06731_ sky130_fd_sc_hd__o211a_1
X_13563_ _03276_ _03504_ VGND VGND VPWR VPWR _03697_ sky130_fd_sc_hd__or2_1
XFILLER_0_137_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10775_ _00163_ _00214_ VGND VGND VPWR VPWR _00868_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15302_ _05478_ _05553_ _05593_ _05594_ VGND VGND VPWR VPWR _05596_ sky130_fd_sc_hd__a211oi_4
X_12514_ _00514_ _02214_ VGND VGND VPWR VPWR _02607_ sky130_fd_sc_hd__nor2_2
X_16282_ _06655_ VGND VGND VPWR VPWR _06657_ sky130_fd_sc_hd__buf_2
X_13494_ _03606_ _03608_ _03619_ VGND VGND VPWR VPWR _03621_ sky130_fd_sc_hd__or3_4
XFILLER_0_42_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_255 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18021_ _08456_ _08457_ VGND VGND VPWR VPWR _08549_ sky130_fd_sc_hd__nor2_1
X_15233_ _05407_ _05416_ _05520_ VGND VGND VPWR VPWR _05521_ sky130_fd_sc_hd__a21oi_1
X_12445_ _02534_ _02537_ VGND VGND VPWR VPWR _02538_ sky130_fd_sc_hd__or2b_1
XFILLER_0_112_508 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_152_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15164_ _07515_ _00461_ _05856_ _03008_ VGND VGND VPWR VPWR _05445_ sky130_fd_sc_hd__a22oi_1
X_12376_ _02330_ _02467_ _02468_ _02328_ VGND VGND VPWR VPWR _02469_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_23_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14115_ _04297_ _04298_ _04107_ _04266_ VGND VGND VPWR VPWR _04300_ sky130_fd_sc_hd__a211oi_2
X_11327_ _01315_ _01419_ VGND VGND VPWR VPWR _01420_ sky130_fd_sc_hd__xor2_1
XFILLER_0_120_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15095_ _00192_ _08876_ _05368_ VGND VGND VPWR VPWR _05370_ sky130_fd_sc_hd__and3_1
XFILLER_0_22_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14046_ _04222_ _04223_ _04224_ VGND VGND VPWR VPWR _04225_ sky130_fd_sc_hd__or3_4
X_18923_ clknet_4_13_0_clk _00077_ VGND VGND VPWR VPWR ApproximateM_inst.lob_16.lob2.genblk1\[9\].genblk1.mux.sel
+ sky130_fd_sc_hd__dfxtp_1
X_11258_ _01339_ _01340_ _01350_ VGND VGND VPWR VPWR _01351_ sky130_fd_sc_hd__o21a_1
X_10209_ _00288_ _00289_ _00290_ VGND VGND VPWR VPWR _00302_ sky130_fd_sc_hd__a21oi_1
X_18854_ clknet_4_6_0_clk net290 VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__dfxtp_1
X_11189_ _00789_ _00790_ VGND VGND VPWR VPWR _01282_ sky130_fd_sc_hd__xor2_2
X_17805_ _08183_ _08255_ _08313_ VGND VGND VPWR VPWR _08315_ sky130_fd_sc_hd__or3_1
X_18785_ _09297_ VGND VGND VPWR VPWR _00086_ sky130_fd_sc_hd__dlymetal6s2s_1
X_15997_ _05736_ _00194_ VGND VGND VPWR VPWR _06346_ sky130_fd_sc_hd__or2_2
X_14948_ _05116_ _05117_ VGND VGND VPWR VPWR _05209_ sky130_fd_sc_hd__or2_1
X_17736_ _01678_ _06442_ _08239_ VGND VGND VPWR VPWR _08240_ sky130_fd_sc_hd__o21a_1
XFILLER_0_49_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14879_ _05132_ _05133_ VGND VGND VPWR VPWR _05134_ sky130_fd_sc_hd__and2_1
X_17667_ _08162_ _08163_ VGND VGND VPWR VPWR _08164_ sky130_fd_sc_hd__xnor2_1
X_16618_ _07020_ VGND VGND VPWR VPWR _07021_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17598_ _07207_ _07665_ _07650_ _06947_ VGND VGND VPWR VPWR _08089_ sky130_fd_sc_hd__a22o_1
XFILLER_0_92_509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16549_ _06942_ _06943_ _06084_ VGND VGND VPWR VPWR _06946_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_128_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_61 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18219_ _08763_ _06398_ _06399_ _07084_ _08764_ VGND VGND VPWR VPWR _08765_ sky130_fd_sc_hd__a311o_1
XFILLER_0_116_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_122_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_131_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09923_ _08529_ _08648_ _08637_ VGND VGND VPWR VPWR _08670_ sky130_fd_sc_hd__o21a_1
XFILLER_0_1_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09854_ _05812_ _06960_ _07897_ _07908_ VGND VGND VPWR VPWR _07919_ sky130_fd_sc_hd__o211a_2
XTAP_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09785_ _07080_ _07156_ _07134_ _07058_ VGND VGND VPWR VPWR _07167_ sky130_fd_sc_hd__a22o_1
XTAP_2406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_107 net40 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_118 _02099_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_129 _04125_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10560_ _00643_ _00651_ _00652_ VGND VGND VPWR VPWR _00653_ sky130_fd_sc_hd__nand3_2
XFILLER_0_64_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_162 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_134_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10491_ _00580_ _00581_ _00582_ _00537_ VGND VGND VPWR VPWR _00584_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_106_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12230_ _02135_ _02322_ VGND VGND VPWR VPWR _02323_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_134_688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12161_ _02240_ _02253_ VGND VGND VPWR VPWR _02254_ sky130_fd_sc_hd__or2_4
XFILLER_0_31_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11112_ _01126_ _01131_ _01130_ VGND VGND VPWR VPWR _01205_ sky130_fd_sc_hd__a21o_1
X_12092_ _02114_ _02184_ VGND VGND VPWR VPWR _02185_ sky130_fd_sc_hd__nor2_1
X_11043_ _06689_ VGND VGND VPWR VPWR _01136_ sky130_fd_sc_hd__inv_4
X_15920_ net192 _06235_ _06263_ VGND VGND VPWR VPWR _06265_ sky130_fd_sc_hd__a21oi_2
X_15851_ _06131_ _06180_ VGND VGND VPWR VPWR _06190_ sky130_fd_sc_hd__or2_1
Xclkbuf_4_3_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_3_0_clk sky130_fd_sc_hd__clkbuf_8
X_14802_ _05036_ _05037_ _05049_ VGND VGND VPWR VPWR _05051_ sky130_fd_sc_hd__a21o_1
X_15782_ _06113_ _06115_ VGND VGND VPWR VPWR _06117_ sky130_fd_sc_hd__xnor2_1
X_18570_ salida\[7\] _09114_ _09118_ salida\[39\] _09128_ VGND VGND VPWR VPWR _09136_
+ sky130_fd_sc_hd__a221o_1
X_12994_ _03026_ _03086_ _02720_ VGND VGND VPWR VPWR _03087_ sky130_fd_sc_hd__a21o_1
X_17521_ _06750_ _07745_ _08003_ VGND VGND VPWR VPWR _08005_ sky130_fd_sc_hd__a21oi_1
X_14733_ _04838_ _04839_ _04972_ _04974_ VGND VGND VPWR VPWR _04975_ sky130_fd_sc_hd__a211o_1
XFILLER_0_153_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11945_ _02036_ _02037_ VGND VGND VPWR VPWR _02038_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_143_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17452_ _07929_ VGND VGND VPWR VPWR _09392_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14664_ _01317_ VGND VGND VPWR VPWR _04900_ sky130_fd_sc_hd__clkbuf_4
X_11876_ _01933_ _01934_ _01935_ VGND VGND VPWR VPWR _01969_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_67_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16403_ _03912_ _06593_ _06594_ VGND VGND VPWR VPWR _06789_ sky130_fd_sc_hd__a21o_1
X_13615_ _03606_ _03608_ _03619_ VGND VGND VPWR VPWR _03753_ sky130_fd_sc_hd__nor3_1
XFILLER_0_129_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10827_ cla_inst.in2\[16\] ApproximateM_inst.lob_16.lob2.genblk2.mux_final.sel ApproximateM_inst.lob_16.lob1.genblk1\[8\].genblk1.mux.sel
+ ApproximateM_inst.lob_16.lob1.genblk1\[7\].genblk1.mux.sel VGND VGND VPWR VPWR _00920_
+ sky130_fd_sc_hd__and4_1
XFILLER_0_145_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17383_ _07747_ _07748_ _07760_ _07758_ VGND VGND VPWR VPWR _07855_ sky130_fd_sc_hd__a31o_1
X_14595_ _03079_ _02980_ _03533_ VGND VGND VPWR VPWR _04825_ sky130_fd_sc_hd__or3_1
XFILLER_0_94_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16334_ _03161_ _02607_ _03170_ VGND VGND VPWR VPWR _06714_ sky130_fd_sc_hd__or3_1
X_13546_ _00183_ _04657_ _04864_ _00184_ VGND VGND VPWR VPWR _03678_ sky130_fd_sc_hd__a22oi_1
X_10758_ _00831_ _00844_ _00850_ VGND VGND VPWR VPWR _00851_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_14_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16265_ _03152_ _02272_ _03104_ _06467_ _06638_ VGND VGND VPWR VPWR _06639_ sky130_fd_sc_hd__o311a_1
X_13477_ _03600_ _03601_ VGND VGND VPWR VPWR _03602_ sky130_fd_sc_hd__xor2_1
X_10689_ _04001_ _04045_ _00765_ _00781_ VGND VGND VPWR VPWR _00782_ sky130_fd_sc_hd__a31o_1
XFILLER_0_35_480 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15216_ _05459_ _05501_ VGND VGND VPWR VPWR _05502_ sky130_fd_sc_hd__xor2_1
X_18004_ _08484_ _08494_ VGND VGND VPWR VPWR _08531_ sky130_fd_sc_hd__or2b_1
XFILLER_0_113_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12428_ _02515_ _02519_ _02520_ VGND VGND VPWR VPWR _02521_ sky130_fd_sc_hd__nor3_2
XFILLER_0_2_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16196_ _06562_ VGND VGND VPWR VPWR _06563_ sky130_fd_sc_hd__buf_2
XFILLER_0_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15147_ _05398_ _05401_ VGND VGND VPWR VPWR _05426_ sky130_fd_sc_hd__and2b_1
X_12359_ _02443_ _02445_ _02375_ VGND VGND VPWR VPWR _02452_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_77_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15078_ _05231_ _05234_ _05232_ VGND VGND VPWR VPWR _05351_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_120_382 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14029_ _03993_ _04205_ VGND VGND VPWR VPWR _04206_ sky130_fd_sc_hd__xor2_1
X_18906_ clknet_4_10_0_clk _00060_ VGND VGND VPWR VPWR cla_inst.in1\[24\] sky130_fd_sc_hd__dfxtp_2
X_18837_ _09336_ VGND VGND VPWR VPWR _00104_ sky130_fd_sc_hd__clkbuf_1
X_09570_ _03487_ _03542_ _03443_ VGND VGND VPWR VPWR _04831_ sky130_fd_sc_hd__a21bo_1
X_18768_ _04725_ net39 _09276_ VGND VGND VPWR VPWR _09284_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17719_ _08016_ _08018_ _08121_ VGND VGND VPWR VPWR _08221_ sky130_fd_sc_hd__nor3_1
X_18699_ net50 _03052_ _09182_ VGND VGND VPWR VPWR _09230_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_198 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09906_ _08365_ _08376_ _08387_ VGND VGND VPWR VPWR _08485_ sky130_fd_sc_hd__a21o_1
XFILLER_0_10_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09837_ _07722_ VGND VGND VPWR VPWR _07733_ sky130_fd_sc_hd__buf_4
XTAP_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09768_ _06971_ VGND VGND VPWR VPWR _06982_ sky130_fd_sc_hd__buf_4
XTAP_2203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09699_ _06202_ _06213_ _06224_ VGND VGND VPWR VPWR _06234_ sky130_fd_sc_hd__nand3_1
XTAP_2236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer60 _05377_ VGND VGND VPWR VPWR net223 sky130_fd_sc_hd__clkbuf_1
XTAP_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer71 cla_inst.in1\[18\] VGND VGND VPWR VPWR net234 sky130_fd_sc_hd__clkbuf_2
XTAP_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer82 _03772_ VGND VGND VPWR VPWR net329 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11730_ _04493_ ApproximateM_inst.lob_16.lob2.genblk1\[12\].genblk1.mux.sel _00179_
+ _00129_ VGND VGND VPWR VPWR _01823_ sky130_fd_sc_hd__and4_1
XTAP_2269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer93 _00333_ VGND VGND VPWR VPWR net340 sky130_fd_sc_hd__clkbuf_1
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11661_ _01742_ _01753_ VGND VGND VPWR VPWR _01754_ sky130_fd_sc_hd__xor2_1
XFILLER_0_95_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13400_ _03371_ _03372_ _03516_ _03517_ VGND VGND VPWR VPWR _03518_ sky130_fd_sc_hd__o211a_2
X_10612_ _00703_ _00704_ VGND VGND VPWR VPWR _00705_ sky130_fd_sc_hd__nor2_1
XFILLER_0_153_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14380_ _02188_ cla_inst.in1\[30\] _09303_ _04515_ VGND VGND VPWR VPWR _04589_ sky130_fd_sc_hd__a22o_1
X_11592_ _01647_ _01649_ VGND VGND VPWR VPWR _01685_ sky130_fd_sc_hd__nand2_1
XFILLER_0_153_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13331_ _03440_ _00206_ _07526_ _03441_ VGND VGND VPWR VPWR _03442_ sky130_fd_sc_hd__and4b_1
XFILLER_0_51_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10543_ _00474_ _00475_ VGND VGND VPWR VPWR _00636_ sky130_fd_sc_hd__and2_1
X_16050_ _06402_ _06403_ _05721_ VGND VGND VPWR VPWR _06404_ sky130_fd_sc_hd__a21o_1
XFILLER_0_107_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_122_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13262_ _03307_ _03309_ VGND VGND VPWR VPWR _03367_ sky130_fd_sc_hd__or2b_1
XFILLER_0_121_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10474_ _00170_ _04067_ VGND VGND VPWR VPWR _00567_ sky130_fd_sc_hd__nand2_1
XFILLER_0_121_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15001_ _05265_ _05266_ VGND VGND VPWR VPWR _05267_ sky130_fd_sc_hd__nor2_1
X_12213_ _02302_ _02304_ _02305_ VGND VGND VPWR VPWR _02306_ sky130_fd_sc_hd__or3_1
X_13193_ net131 _03266_ _03291_ VGND VGND VPWR VPWR _03294_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_20_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12144_ _02110_ _02109_ VGND VGND VPWR VPWR _02237_ sky130_fd_sc_hd__and2b_1
XFILLER_0_102_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12075_ _01899_ _01904_ VGND VGND VPWR VPWR _02168_ sky130_fd_sc_hd__nor2_1
X_16952_ _07285_ _07295_ VGND VGND VPWR VPWR _07385_ sky130_fd_sc_hd__nand2_1
X_11026_ _01072_ _01074_ _01117_ VGND VGND VPWR VPWR _01119_ sky130_fd_sc_hd__and3_1
X_15903_ _03011_ _03154_ VGND VGND VPWR VPWR _06247_ sky130_fd_sc_hd__and2_1
X_16883_ _07307_ _07309_ VGND VGND VPWR VPWR _07310_ sky130_fd_sc_hd__xor2_1
X_18622_ salida\[28\] _09159_ _09160_ salida\[60\] _09163_ VGND VGND VPWR VPWR _09173_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_2_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15834_ _06171_ _06172_ VGND VGND VPWR VPWR _06173_ sky130_fd_sc_hd__nor2_1
XFILLER_0_87_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18553_ _09124_ VGND VGND VPWR VPWR _09125_ sky130_fd_sc_hd__buf_4
X_15765_ _05966_ _06045_ VGND VGND VPWR VPWR _06098_ sky130_fd_sc_hd__and2b_1
X_12977_ _00121_ _03069_ _03024_ VGND VGND VPWR VPWR _03070_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_99_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17504_ _07985_ _07986_ VGND VGND VPWR VPWR _07987_ sky130_fd_sc_hd__and2_1
XFILLER_0_86_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11928_ _02017_ _02020_ VGND VGND VPWR VPWR _02021_ sky130_fd_sc_hd__and2_1
X_14716_ _03569_ _03582_ _02978_ VGND VGND VPWR VPWR _04957_ sky130_fd_sc_hd__mux2_1
X_15696_ _06004_ VGND VGND VPWR VPWR _06023_ sky130_fd_sc_hd__inv_2
X_18484_ _09047_ _06559_ _09050_ VGND VGND VPWR VPWR _09051_ sky130_fd_sc_hd__or3b_4
XTAP_2770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14647_ _04867_ _04868_ _04879_ VGND VGND VPWR VPWR _04881_ sky130_fd_sc_hd__and3_1
X_17435_ _07802_ _07803_ _07801_ VGND VGND VPWR VPWR _07912_ sky130_fd_sc_hd__a21bo_1
X_11859_ _01950_ _01951_ ApproximateM_inst.lob_16.lob2.genblk1\[5\].genblk1.mux.sel
+ _03399_ VGND VGND VPWR VPWR _01952_ sky130_fd_sc_hd__and4b_1
XFILLER_0_7_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_18 _01115_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_216 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14578_ _04803_ _04804_ _04628_ _04698_ VGND VGND VPWR VPWR _04806_ sky130_fd_sc_hd__a211oi_1
XANTENNA_29 _01115_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17366_ _07834_ _07835_ VGND VGND VPWR VPWR _07836_ sky130_fd_sc_hd__nor2_1
XFILLER_0_103_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13529_ _03656_ _03658_ VGND VGND VPWR VPWR _03659_ sky130_fd_sc_hd__or2_2
X_16317_ _03047_ _07766_ _03150_ VGND VGND VPWR VPWR _06695_ sky130_fd_sc_hd__or3_1
XFILLER_0_55_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_87 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17297_ _07749_ _07760_ VGND VGND VPWR VPWR _07761_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_153_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_772 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_603 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_125_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16248_ _06618_ _06619_ _03152_ VGND VGND VPWR VPWR _06620_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput103 net103 VGND VGND VPWR VPWR o_wb_data[28] sky130_fd_sc_hd__clkbuf_4
Xoutput114 net114 VGND VGND VPWR VPWR o_wb_data[9] sky130_fd_sc_hd__clkbuf_4
X_16179_ _06544_ VGND VGND VPWR VPWR _06545_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_6 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09622_ ApproximateM_inst.lob_16.lob2.genblk1\[10\].genblk1.mux.sel VGND VGND VPWR
+ VPWR _05399_ sky130_fd_sc_hd__buf_4
XFILLER_0_78_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09553_ _04635_ VGND VGND VPWR VPWR _04646_ sky130_fd_sc_hd__buf_6
XFILLER_0_77_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09484_ _03771_ VGND VGND VPWR VPWR _03892_ sky130_fd_sc_hd__buf_6
XFILLER_0_53_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_94 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_109_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_391 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_767 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_131_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_143_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_131_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10190_ _03848_ _03782_ _04569_ _04384_ VGND VGND VPWR VPWR _00283_ sky130_fd_sc_hd__and4_1
X_12900_ _00189_ VGND VGND VPWR VPWR _02993_ sky130_fd_sc_hd__clkbuf_4
X_13880_ _04024_ _04041_ _04042_ VGND VGND VPWR VPWR _04043_ sky130_fd_sc_hd__nor3_1
X_12831_ _00891_ VGND VGND VPWR VPWR _02924_ sky130_fd_sc_hd__inv_2
XTAP_2000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_623 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15550_ _05861_ _05862_ _05757_ VGND VGND VPWR VPWR _05865_ sky130_fd_sc_hd__o21ai_1
XTAP_2044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12762_ _01790_ _01798_ _01799_ VGND VGND VPWR VPWR _02855_ sky130_fd_sc_hd__nor3_1
XTAP_2055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14501_ net179 _04579_ _04573_ VGND VGND VPWR VPWR _04721_ sky130_fd_sc_hd__a21bo_1
XTAP_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11713_ _01784_ _01787_ _01804_ _01805_ VGND VGND VPWR VPWR _01806_ sky130_fd_sc_hd__o211ai_2
X_15481_ _05614_ _05710_ VGND VGND VPWR VPWR _05790_ sky130_fd_sc_hd__nor2_1
XTAP_2099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12693_ _02755_ _02785_ VGND VGND VPWR VPWR _02786_ sky130_fd_sc_hd__nand2_1
XTAP_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14432_ _01139_ VGND VGND VPWR VPWR _04647_ sky130_fd_sc_hd__clkbuf_4
XTAP_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17220_ _02633_ _07676_ _03201_ VGND VGND VPWR VPWR _07677_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_126_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11644_ _01735_ _01736_ VGND VGND VPWR VPWR _01737_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_83_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17151_ _07590_ _07600_ VGND VGND VPWR VPWR _07601_ sky130_fd_sc_hd__xnor2_1
X_14363_ _02986_ _07134_ _04568_ _04570_ VGND VGND VPWR VPWR _04571_ sky130_fd_sc_hd__nand4_2
XFILLER_0_64_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput16 i_wb_addr[22] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__clkbuf_1
X_11575_ _01658_ _01666_ _01667_ VGND VGND VPWR VPWR _01668_ sky130_fd_sc_hd__a21boi_1
Xinput27 i_wb_addr[3] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__clkbuf_4
X_16102_ _02966_ _06459_ VGND VGND VPWR VPWR _06461_ sky130_fd_sc_hd__nor2_1
Xinput38 i_wb_data[12] VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__buf_2
XFILLER_0_24_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13314_ _03416_ _03422_ _03423_ VGND VGND VPWR VPWR _03424_ sky130_fd_sc_hd__nand3_2
XFILLER_0_135_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10526_ _00445_ _00446_ _00438_ VGND VGND VPWR VPWR _00619_ sky130_fd_sc_hd__a21bo_1
Xinput49 i_wb_data[22] VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__clkbuf_2
X_17082_ _07523_ _07524_ VGND VGND VPWR VPWR _07527_ sky130_fd_sc_hd__nand2_1
X_14294_ _00173_ _00175_ _05388_ _05050_ VGND VGND VPWR VPWR _04496_ sky130_fd_sc_hd__and4_1
XFILLER_0_52_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_134_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16033_ _06383_ _06385_ _03588_ VGND VGND VPWR VPWR _06386_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_122_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13245_ _00747_ _03203_ _03347_ _03348_ VGND VGND VPWR VPWR _03349_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_122_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10457_ _00548_ _00549_ VGND VGND VPWR VPWR _00550_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_149_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13176_ _03272_ _03274_ VGND VGND VPWR VPWR _03275_ sky130_fd_sc_hd__or2_1
X_10388_ _00476_ _00480_ VGND VGND VPWR VPWR _00481_ sky130_fd_sc_hd__xnor2_1
X_12127_ _02219_ _02209_ VGND VGND VPWR VPWR _02220_ sky130_fd_sc_hd__xnor2_1
X_17984_ _02167_ _08424_ _02174_ VGND VGND VPWR VPWR _08510_ sky130_fd_sc_hd__o21ai_1
X_12058_ _02148_ _02134_ _02149_ _02150_ VGND VGND VPWR VPWR _02151_ sky130_fd_sc_hd__or4b_4
X_16935_ _03101_ _06436_ _07366_ VGND VGND VPWR VPWR _07367_ sky130_fd_sc_hd__o21a_1
XFILLER_0_74_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11009_ _01098_ _01100_ VGND VGND VPWR VPWR _01102_ sky130_fd_sc_hd__or2b_1
X_16866_ _06562_ _07290_ VGND VGND VPWR VPWR _07291_ sky130_fd_sc_hd__nor2_1
X_18605_ _09125_ VGND VGND VPWR VPWR _09162_ sky130_fd_sc_hd__buf_2
X_15817_ _03012_ _03072_ _03149_ _03010_ VGND VGND VPWR VPWR _06154_ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16797_ _03324_ _06529_ _06814_ _02099_ VGND VGND VPWR VPWR _07216_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_59_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18536_ net9 net12 net11 net15 VGND VGND VPWR VPWR _09106_ sky130_fd_sc_hd__or4_1
X_15748_ net197 _06079_ VGND VGND VPWR VPWR _06080_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18467_ _03036_ _06295_ _09029_ _09032_ VGND VGND VPWR VPWR _09033_ sky130_fd_sc_hd__o211ai_1
X_15679_ _06002_ _06003_ _05957_ _05931_ VGND VGND VPWR VPWR _06005_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_28_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17418_ _07891_ _07892_ VGND VGND VPWR VPWR _07893_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18398_ _04406_ _07592_ _08957_ VGND VGND VPWR VPWR _08958_ sky130_fd_sc_hd__nand3_1
XFILLER_0_28_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17349_ _06421_ _07806_ _07807_ _07817_ VGND VGND VPWR VPWR _07818_ sky130_fd_sc_hd__a31o_1
XFILLER_0_16_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_77 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_83 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09605_ ApproximateM_inst.lob_16.lob2.genblk1\[8\].genblk1.mux.sel VGND VGND VPWR
+ VPWR _05213_ sky130_fd_sc_hd__buf_4
X_09536_ _04449_ VGND VGND VPWR VPWR _04460_ sky130_fd_sc_hd__buf_6
XFILLER_0_78_453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_149_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09467_ _03553_ _03563_ _03695_ VGND VGND VPWR VPWR _03706_ sky130_fd_sc_hd__nand3_1
XFILLER_0_109_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_108_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_512 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11360_ _01362_ _01437_ VGND VGND VPWR VPWR _01453_ sky130_fd_sc_hd__nand2_1
XFILLER_0_132_731 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10311_ _00170_ _00165_ VGND VGND VPWR VPWR _00404_ sky130_fd_sc_hd__nand2_1
X_11291_ _01299_ _01302_ VGND VGND VPWR VPWR _01384_ sky130_fd_sc_hd__and2_1
XFILLER_0_104_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13030_ _02971_ _03122_ VGND VGND VPWR VPWR _09355_ sky130_fd_sc_hd__nand2_1
X_10242_ _00330_ _00331_ _00334_ _00305_ VGND VGND VPWR VPWR _00335_ sky130_fd_sc_hd__o2bb2a_1
X_10173_ _00245_ _00246_ _00265_ VGND VGND VPWR VPWR _00266_ sky130_fd_sc_hd__a21o_1
XFILLER_0_28_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14981_ _05156_ _05155_ VGND VGND VPWR VPWR _05245_ sky130_fd_sc_hd__and2b_1
X_16720_ _07129_ _07131_ VGND VGND VPWR VPWR _07132_ sky130_fd_sc_hd__xnor2_2
X_13932_ _04097_ _04098_ VGND VGND VPWR VPWR _04100_ sky130_fd_sc_hd__xor2_2
XFILLER_0_89_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13863_ _03862_ _03872_ VGND VGND VPWR VPWR _04025_ sky130_fd_sc_hd__or2_1
X_16651_ _07055_ _07056_ VGND VGND VPWR VPWR _07057_ sky130_fd_sc_hd__xnor2_1
X_12814_ _02899_ _02905_ _02906_ VGND VGND VPWR VPWR _02907_ sky130_fd_sc_hd__and3_2
X_15602_ _05918_ _05919_ VGND VGND VPWR VPWR _05922_ sky130_fd_sc_hd__nor2_1
X_13794_ _03945_ _03947_ _03948_ VGND VGND VPWR VPWR _03949_ sky130_fd_sc_hd__nor3b_4
X_16582_ _06934_ _06935_ _06980_ VGND VGND VPWR VPWR _06983_ sky130_fd_sc_hd__or3b_4
XFILLER_0_57_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18321_ _02871_ _02881_ VGND VGND VPWR VPWR _08875_ sky130_fd_sc_hd__nand2_1
X_15533_ _05737_ _05755_ _05844_ VGND VGND VPWR VPWR _05847_ sky130_fd_sc_hd__or3_1
XTAP_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12745_ _02749_ _02748_ VGND VGND VPWR VPWR _02838_ sky130_fd_sc_hd__or2b_1
XTAP_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15464_ _05688_ _05770_ VGND VGND VPWR VPWR _05772_ sky130_fd_sc_hd__or2_1
XTAP_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18252_ _08725_ _08726_ _08728_ _08799_ VGND VGND VPWR VPWR _08801_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_44_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12676_ _02766_ _02767_ VGND VGND VPWR VPWR _02769_ sky130_fd_sc_hd__xor2_1
XFILLER_0_84_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_127_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14415_ _04470_ _04488_ _04626_ _04627_ VGND VGND VPWR VPWR _04628_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_65_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17203_ _06750_ _07650_ _07656_ VGND VGND VPWR VPWR _07659_ sky130_fd_sc_hd__a21oi_1
X_11627_ _01716_ _01717_ _01718_ _01710_ VGND VGND VPWR VPWR _01720_ sky130_fd_sc_hd__a22o_1
X_15395_ _05549_ _05598_ _05696_ VGND VGND VPWR VPWR _05697_ sky130_fd_sc_hd__a21oi_1
X_18183_ _08715_ _08723_ VGND VGND VPWR VPWR _08726_ sky130_fd_sc_hd__nor2_1
XFILLER_0_142_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14346_ _04399_ _04400_ VGND VGND VPWR VPWR _04553_ sky130_fd_sc_hd__nor2_1
XFILLER_0_108_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17134_ _03198_ _04956_ _07572_ _07583_ VGND VGND VPWR VPWR _07584_ sky130_fd_sc_hd__a211o_1
X_11558_ _07352_ _05050_ _01647_ _01648_ VGND VGND VPWR VPWR _01651_ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10509_ _00467_ _00486_ _00487_ _00488_ VGND VGND VPWR VPWR _00602_ sky130_fd_sc_hd__and4_1
XFILLER_0_12_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17065_ _07421_ _07422_ VGND VGND VPWR VPWR _07508_ sky130_fd_sc_hd__nor2_1
X_14277_ _04475_ _00715_ _07526_ _04476_ VGND VGND VPWR VPWR _04477_ sky130_fd_sc_hd__and4b_1
XFILLER_0_111_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11489_ _01529_ _01530_ _01532_ VGND VGND VPWR VPWR _01582_ sky130_fd_sc_hd__a21o_1
XFILLER_0_150_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16016_ _06331_ _06365_ _06366_ VGND VGND VPWR VPWR _06367_ sky130_fd_sc_hd__a21o_1
XFILLER_0_123_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13228_ _03318_ _03330_ VGND VGND VPWR VPWR _03331_ sky130_fd_sc_hd__xor2_2
XFILLER_0_21_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13159_ _03254_ _03255_ _03247_ VGND VGND VPWR VPWR _03257_ sky130_fd_sc_hd__a21o_1
XTAP_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17967_ _08487_ _08488_ _08489_ VGND VGND VPWR VPWR _08491_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_109_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16918_ _07248_ _07252_ _07249_ VGND VGND VPWR VPWR _07348_ sky130_fd_sc_hd__o21ai_2
X_17898_ _08252_ _08324_ VGND VGND VPWR VPWR _08416_ sky130_fd_sc_hd__or2b_1
XFILLER_0_26_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16849_ _00167_ _07179_ _07272_ VGND VGND VPWR VPWR _07273_ sky130_fd_sc_hd__o21a_1
XFILLER_0_149_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18519_ _03913_ _07086_ _08141_ _09087_ VGND VGND VPWR VPWR _09088_ sky130_fd_sc_hd__o31a_1
XFILLER_0_47_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_567 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_114_742 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_98_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10860_ _00948_ _00952_ VGND VGND VPWR VPWR _00953_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_78_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09519_ _04231_ _04253_ _04263_ VGND VGND VPWR VPWR _04274_ sky130_fd_sc_hd__a21bo_1
XPHY_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10791_ _00876_ _00880_ _00883_ VGND VGND VPWR VPWR _00884_ sky130_fd_sc_hd__o21a_1
XFILLER_0_94_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12530_ _02482_ _02532_ VGND VGND VPWR VPWR _02623_ sky130_fd_sc_hd__or2_1
XPHY_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12461_ _02551_ _02553_ VGND VGND VPWR VPWR _02554_ sky130_fd_sc_hd__nand2_1
XFILLER_0_136_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14200_ _04390_ _04391_ _04392_ VGND VGND VPWR VPWR _04393_ sky130_fd_sc_hd__nor3_2
XFILLER_0_62_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11412_ _01504_ VGND VGND VPWR VPWR _01505_ sky130_fd_sc_hd__buf_4
X_15180_ _05362_ _05360_ VGND VGND VPWR VPWR _05462_ sky130_fd_sc_hd__and2b_1
XFILLER_0_50_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12392_ _02422_ _02430_ VGND VGND VPWR VPWR _02485_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_61_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14131_ _04127_ _04141_ _04139_ VGND VGND VPWR VPWR _04317_ sky130_fd_sc_hd__a21o_1
X_11343_ _01434_ _01435_ VGND VGND VPWR VPWR _01436_ sky130_fd_sc_hd__or2_1
XFILLER_0_120_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_132_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14062_ _03533_ _03549_ _03099_ VGND VGND VPWR VPWR _04243_ sky130_fd_sc_hd__mux2_2
X_11274_ _01335_ _01336_ _01079_ _01147_ VGND VGND VPWR VPWR _01367_ sky130_fd_sc_hd__o211a_1
X_13013_ _03103_ _03105_ _03090_ VGND VGND VPWR VPWR _03106_ sky130_fd_sc_hd__mux2_1
X_10225_ _06732_ VGND VGND VPWR VPWR _00318_ sky130_fd_sc_hd__buf_4
X_18870_ clknet_4_13_0_clk net245 VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__dfxtp_1
X_17821_ _08329_ _08330_ _08331_ VGND VGND VPWR VPWR _08332_ sky130_fd_sc_hd__or3_1
X_10156_ _00164_ _00248_ VGND VGND VPWR VPWR _00249_ sky130_fd_sc_hd__nand2_1
X_17752_ _08167_ _08170_ VGND VGND VPWR VPWR _08257_ sky130_fd_sc_hd__nand2_1
X_14964_ _05223_ _05225_ _05119_ VGND VGND VPWR VPWR _05227_ sky130_fd_sc_hd__a21o_1
X_10087_ _00179_ VGND VGND VPWR VPWR _00180_ sky130_fd_sc_hd__buf_4
X_16703_ _07113_ _06655_ _06946_ _07026_ VGND VGND VPWR VPWR _07114_ sky130_fd_sc_hd__and4_1
X_13915_ _04081_ _03185_ _03060_ VGND VGND VPWR VPWR _04082_ sky130_fd_sc_hd__mux2_1
X_17683_ _08171_ _08181_ VGND VGND VPWR VPWR _08182_ sky130_fd_sc_hd__xnor2_1
X_14895_ _05149_ _05150_ _05144_ VGND VGND VPWR VPWR _05152_ sky130_fd_sc_hd__a21oi_1
X_16634_ _07033_ _07034_ _00207_ VGND VGND VPWR VPWR _07039_ sky130_fd_sc_hd__o21a_4
X_13846_ _03857_ _03858_ _03874_ VGND VGND VPWR VPWR _04006_ sky130_fd_sc_hd__a21o_1
XFILLER_0_76_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13777_ _03201_ VGND VGND VPWR VPWR _03930_ sky130_fd_sc_hd__clkbuf_8
X_16565_ _06950_ _06963_ VGND VGND VPWR VPWR _06964_ sky130_fd_sc_hd__xor2_1
X_10989_ ApproximateM_inst.lob_16.lob2.genblk1\[4\].genblk1.mux.sel VGND VGND VPWR
+ VPWR _01082_ sky130_fd_sc_hd__buf_4
X_18304_ _08853_ _08855_ VGND VGND VPWR VPWR _08857_ sky130_fd_sc_hd__nor2_1
X_15516_ _05809_ _05810_ _05827_ VGND VGND VPWR VPWR _05828_ sky130_fd_sc_hd__o21a_1
XFILLER_0_29_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_84_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12728_ _02810_ _02812_ VGND VGND VPWR VPWR _02821_ sky130_fd_sc_hd__and2_1
XFILLER_0_45_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16496_ _06812_ net150 VGND VGND VPWR VPWR _06889_ sky130_fd_sc_hd__nand2_8
XFILLER_0_72_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_84_286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_127_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18235_ _08776_ _08780_ VGND VGND VPWR VPWR _08782_ sky130_fd_sc_hd__and2_1
X_15447_ _05740_ _05662_ _05751_ VGND VGND VPWR VPWR _05753_ sky130_fd_sc_hd__and3_1
X_12659_ _02742_ _02743_ _02735_ VGND VGND VPWR VPWR _02752_ sky130_fd_sc_hd__a21o_1
XFILLER_0_25_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_191 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_108_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18166_ _07332_ _07665_ _08260_ _08625_ VGND VGND VPWR VPWR _08707_ sky130_fd_sc_hd__or4b_2
X_15378_ _07668_ _01139_ _01223_ _03009_ VGND VGND VPWR VPWR _05678_ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17117_ _02347_ _06510_ _02259_ VGND VGND VPWR VPWR _07565_ sky130_fd_sc_hd__a21o_1
XFILLER_0_123_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14329_ _04531_ _04532_ _04492_ VGND VGND VPWR VPWR _04534_ sky130_fd_sc_hd__o21ai_2
Xmax_cap124 _00600_ VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18097_ _08617_ _08618_ _08631_ VGND VGND VPWR VPWR _08632_ sky130_fd_sc_hd__and3_1
XFILLER_0_13_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap135 _03375_ VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__buf_1
XFILLER_0_40_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17048_ _02188_ _06889_ VGND VGND VPWR VPWR _07489_ sky130_fd_sc_hd__and2_2
XFILLER_0_40_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_592 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09870_ _07286_ _08028_ _08082_ _08060_ VGND VGND VPWR VPWR _08093_ sky130_fd_sc_hd__a211o_1
XTAP_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18999_ clknet_4_7_0_clk _09365_ VGND VGND VPWR VPWR salida\[52\] sky130_fd_sc_hd__dfxtp_1
XTAP_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_331 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_134_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_145_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10010_ _09352_ VGND VGND VPWR VPWR _09353_ sky130_fd_sc_hd__buf_4
X_09999_ _07482_ _07908_ _09339_ _09340_ VGND VGND VPWR VPWR _09342_ sky130_fd_sc_hd__a211o_2
X_11961_ _01979_ _01983_ _01982_ VGND VGND VPWR VPWR _02054_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_98_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10912_ _04700_ VGND VGND VPWR VPWR _01005_ sky130_fd_sc_hd__clkbuf_8
X_13700_ _00203_ _05921_ VGND VGND VPWR VPWR _03846_ sky130_fd_sc_hd__nand2_1
X_14680_ _04904_ _04905_ _04916_ VGND VGND VPWR VPWR _04917_ sky130_fd_sc_hd__o21a_1
X_11892_ _01892_ _01894_ _01893_ VGND VGND VPWR VPWR _01985_ sky130_fd_sc_hd__o21a_1
XFILLER_0_98_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13631_ _03595_ _03602_ _03597_ VGND VGND VPWR VPWR _03770_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_79_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10843_ _03345_ net170 _00145_ ApproximateM_inst.lob_16.lob1.genblk1\[2\].genblk1.mux.sel
+ VGND VGND VPWR VPWR _00936_ sky130_fd_sc_hd__nand4_2
XFILLER_0_67_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13562_ _03692_ _03694_ VGND VGND VPWR VPWR _03696_ sky130_fd_sc_hd__xor2_2
X_16350_ _01677_ _06623_ VGND VGND VPWR VPWR _06730_ sky130_fd_sc_hd__or2_1
X_10774_ _00860_ _00866_ VGND VGND VPWR VPWR _00867_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_82_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15301_ _05574_ _05592_ VGND VGND VPWR VPWR _05594_ sky130_fd_sc_hd__and2_1
X_12513_ _02556_ _02594_ _02603_ VGND VGND VPWR VPWR _02606_ sky130_fd_sc_hd__a21oi_1
X_16281_ _06427_ _06651_ VGND VGND VPWR VPWR _06655_ sky130_fd_sc_hd__nor2_2
XFILLER_0_136_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13493_ _03606_ _03608_ _03619_ VGND VGND VPWR VPWR _03620_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_82_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18020_ _08546_ _08547_ VGND VGND VPWR VPWR _08548_ sky130_fd_sc_hd__nor2_1
XFILLER_0_151_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15232_ _05404_ _05406_ VGND VGND VPWR VPWR _05520_ sky130_fd_sc_hd__and2b_1
X_12444_ _02535_ _02536_ VGND VGND VPWR VPWR _02537_ sky130_fd_sc_hd__xor2_2
XFILLER_0_152_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15163_ _03006_ _01678_ VGND VGND VPWR VPWR _05444_ sky130_fd_sc_hd__nand2_1
XFILLER_0_151_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12375_ _02321_ _02325_ _02327_ VGND VGND VPWR VPWR _02468_ sky130_fd_sc_hd__a21o_1
XFILLER_0_50_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14114_ _04107_ _04266_ _04297_ _04298_ VGND VGND VPWR VPWR _04299_ sky130_fd_sc_hd__o211a_2
XFILLER_0_1_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11326_ _00105_ _01418_ VGND VGND VPWR VPWR _01419_ sky130_fd_sc_hd__nor2_2
X_15094_ _00192_ _08876_ _05368_ VGND VGND VPWR VPWR _05369_ sky130_fd_sc_hd__a21oi_1
X_14045_ _04046_ _04048_ VGND VGND VPWR VPWR _04224_ sky130_fd_sc_hd__nor2_1
X_18922_ clknet_4_9_0_clk _00076_ VGND VGND VPWR VPWR ApproximateM_inst.lob_16.lob2.genblk1\[8\].genblk1.mux.sel
+ sky130_fd_sc_hd__dfxtp_2
X_11257_ _01341_ _01349_ VGND VGND VPWR VPWR _01350_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_66_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10208_ _00299_ _00300_ VGND VGND VPWR VPWR _00301_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_66_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18853_ clknet_4_6_0_clk net292 VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__dfxtp_1
X_11188_ net214 _00958_ VGND VGND VPWR VPWR _01281_ sky130_fd_sc_hd__nor2_1
X_17804_ _08183_ _08255_ _08313_ VGND VGND VPWR VPWR _08314_ sky130_fd_sc_hd__o21ai_2
X_10139_ _00142_ _00159_ VGND VGND VPWR VPWR _00232_ sky130_fd_sc_hd__nor2_1
X_18784_ _09273_ _09296_ VGND VGND VPWR VPWR _09297_ sky130_fd_sc_hd__and2_1
X_15996_ _06084_ _00878_ VGND VGND VPWR VPWR _06345_ sky130_fd_sc_hd__or2_2
X_17735_ _06425_ _06443_ VGND VGND VPWR VPWR _08239_ sky130_fd_sc_hd__nor2_1
X_14947_ _05113_ _05114_ VGND VGND VPWR VPWR _05208_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17666_ _07039_ net145 VGND VGND VPWR VPWR _08163_ sky130_fd_sc_hd__nand2_1
X_14878_ _05124_ _05131_ VGND VGND VPWR VPWR _05133_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16617_ _06950_ _06963_ VGND VGND VPWR VPWR _07020_ sky130_fd_sc_hd__nor2_1
X_13829_ _09166_ cla_inst.in2\[29\] _03673_ _00211_ VGND VGND VPWR VPWR _03987_ sky130_fd_sc_hd__and4_1
X_17597_ _07302_ _07303_ _07314_ _07516_ VGND VGND VPWR VPWR _08088_ sky130_fd_sc_hd__or4_1
XFILLER_0_9_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16548_ _06562_ _06571_ _06874_ _06944_ VGND VGND VPWR VPWR _06945_ sky130_fd_sc_hd__or4_4
XFILLER_0_58_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16479_ sel_op\[0\] _06804_ VGND VGND VPWR VPWR _06870_ sky130_fd_sc_hd__or2_1
XFILLER_0_26_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18218_ _08763_ _06399_ _06398_ VGND VGND VPWR VPWR _08764_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_143_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18149_ _06397_ _06790_ _08688_ _03052_ VGND VGND VPWR VPWR _08689_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_124_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_142_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09922_ _08529_ _08637_ _08648_ VGND VGND VPWR VPWR _08659_ sky130_fd_sc_hd__nor3_2
XFILLER_0_40_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09853_ _07886_ _07493_ _07482_ VGND VGND VPWR VPWR _07908_ sky130_fd_sc_hd__nand3b_4
XTAP_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09784_ _07102_ VGND VGND VPWR VPWR _07156_ sky130_fd_sc_hd__buf_4
XFILLER_0_99_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_108 net40 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_119 _02099_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_107_826 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10490_ _00537_ _00580_ _00581_ _00582_ VGND VGND VPWR VPWR _00583_ sky130_fd_sc_hd__or4_4
XFILLER_0_17_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12160_ _02243_ _02251_ _02252_ VGND VGND VPWR VPWR _02253_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_102_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11111_ _01181_ _01201_ _01077_ _01203_ VGND VGND VPWR VPWR _01204_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_102_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12091_ _05747_ _00213_ _02112_ _02113_ VGND VGND VPWR VPWR _02184_ sky130_fd_sc_hd__o2bb2a_1
X_11042_ _01121_ _01133_ VGND VGND VPWR VPWR _01135_ sky130_fd_sc_hd__nand2_1
X_15850_ _04562_ _05623_ _06152_ _03124_ _06189_ VGND VGND VPWR VPWR _09372_ sky130_fd_sc_hd__a221o_1
XFILLER_0_36_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14801_ _05047_ _05048_ VGND VGND VPWR VPWR _05049_ sky130_fd_sc_hd__xnor2_1
X_15781_ _06035_ _06044_ _06114_ VGND VGND VPWR VPWR _06115_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_99_643 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12993_ _00223_ VGND VGND VPWR VPWR _03086_ sky130_fd_sc_hd__clkbuf_4
X_17520_ _06750_ _07745_ _08003_ VGND VGND VPWR VPWR _08004_ sky130_fd_sc_hd__and3_1
X_14732_ _02986_ _08224_ _04970_ _04971_ VGND VGND VPWR VPWR _04974_ sky130_fd_sc_hd__a22oi_2
X_11944_ _01948_ _01947_ VGND VGND VPWR VPWR _02037_ sky130_fd_sc_hd__and2b_1
XFILLER_0_98_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17451_ _07905_ _07909_ _07928_ _06463_ _03108_ VGND VGND VPWR VPWR _07929_ sky130_fd_sc_hd__a32o_2
X_14663_ _04896_ _04898_ VGND VGND VPWR VPWR _04899_ sky130_fd_sc_hd__nor2_2
XFILLER_0_86_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11875_ _01961_ _01965_ _01966_ _01967_ VGND VGND VPWR VPWR _01968_ sky130_fd_sc_hd__or4_4
XFILLER_0_129_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16402_ _06337_ _06335_ _06336_ _06598_ _06786_ VGND VGND VPWR VPWR _06788_ sky130_fd_sc_hd__a311o_1
X_13614_ _03622_ _03623_ _03646_ VGND VGND VPWR VPWR _03752_ sky130_fd_sc_hd__nand3_2
X_10826_ _00912_ _00913_ _00917_ VGND VGND VPWR VPWR _00919_ sky130_fd_sc_hd__a21oi_1
X_17382_ _07851_ _07852_ VGND VGND VPWR VPWR _07854_ sky130_fd_sc_hd__or2_1
XFILLER_0_39_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14594_ _04818_ _04820_ _04823_ VGND VGND VPWR VPWR _04824_ sky130_fd_sc_hd__o21a_1
XFILLER_0_6_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16333_ _01503_ _03083_ _03166_ _03086_ _06477_ _03161_ VGND VGND VPWR VPWR _06713_
+ sky130_fd_sc_hd__mux4_1
X_13545_ _03464_ _03437_ VGND VGND VPWR VPWR _03677_ sky130_fd_sc_hd__and2b_1
X_10757_ _00848_ _00123_ _00849_ VGND VGND VPWR VPWR _00850_ sky130_fd_sc_hd__nor3b_1
XFILLER_0_54_256 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_124_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13476_ _03990_ _05964_ VGND VGND VPWR VPWR _03601_ sky130_fd_sc_hd__nand2_1
X_16264_ _03089_ _06637_ VGND VGND VPWR VPWR _06638_ sky130_fd_sc_hd__or2_1
X_10688_ _03859_ _03793_ _04056_ _03673_ VGND VGND VPWR VPWR _00781_ sky130_fd_sc_hd__and4_1
XFILLER_0_70_738 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_152_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18003_ _08499_ _08500_ VGND VGND VPWR VPWR _08530_ sky130_fd_sc_hd__nand2_1
XFILLER_0_35_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15215_ _05499_ _05500_ VGND VGND VPWR VPWR _05501_ sky130_fd_sc_hd__and2_1
X_12427_ _02448_ _02514_ _02513_ VGND VGND VPWR VPWR _02520_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_106_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16195_ _07657_ _06541_ VGND VGND VPWR VPWR _06562_ sky130_fd_sc_hd__nand2_1
XFILLER_0_112_328 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_140_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15146_ _03035_ _03116_ _03537_ VGND VGND VPWR VPWR _05425_ sky130_fd_sc_hd__mux2_1
X_12358_ _02450_ VGND VGND VPWR VPWR _02451_ sky130_fd_sc_hd__inv_2
X_11309_ _01320_ _01322_ VGND VGND VPWR VPWR _01402_ sky130_fd_sc_hd__or2b_1
X_15077_ _05250_ _05251_ VGND VGND VPWR VPWR _05350_ sky130_fd_sc_hd__or2_1
X_12289_ _02228_ _02351_ _02350_ VGND VGND VPWR VPWR _02382_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_121_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14028_ _04196_ _04204_ VGND VGND VPWR VPWR _04205_ sky130_fd_sc_hd__xnor2_1
X_18905_ clknet_4_10_0_clk _00059_ VGND VGND VPWR VPWR cla_inst.in1\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_120_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18836_ net60 op_code\[3\] _09331_ VGND VGND VPWR VPWR _09336_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18767_ _09283_ VGND VGND VPWR VPWR _00080_ sky130_fd_sc_hd__buf_1
X_15979_ _00908_ _02963_ VGND VGND VPWR VPWR _06326_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17718_ _08120_ _08219_ VGND VGND VPWR VPWR _08220_ sky130_fd_sc_hd__nor2_1
X_18698_ net49 _09190_ _09229_ VGND VGND VPWR VPWR _00058_ sky130_fd_sc_hd__o21a_1
XFILLER_0_77_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17649_ _03120_ _05425_ _08140_ _08144_ VGND VGND VPWR VPWR _08145_ sky130_fd_sc_hd__o211a_1
XFILLER_0_148_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_147_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_724 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_116_623 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_61 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09905_ _08442_ _08463_ VGND VGND VPWR VPWR _08474_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09836_ cla_inst.in1\[28\] VGND VGND VPWR VPWR _07722_ sky130_fd_sc_hd__clkbuf_4
XTAP_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09767_ ApproximateM_inst.lob_16.lob2.genblk1\[2\].genblk1.mux.sel VGND VGND VPWR
+ VPWR _06971_ sky130_fd_sc_hd__buf_4
XTAP_2204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09698_ _03509_ _03804_ _03399_ _03531_ VGND VGND VPWR VPWR _06224_ sky130_fd_sc_hd__a22o_2
XTAP_2226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer50 net212 VGND VGND VPWR VPWR net213 sky130_fd_sc_hd__clkbuf_1
XTAP_2237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer61 _05377_ VGND VGND VPWR VPWR net224 sky130_fd_sc_hd__clkbuf_1
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer72 net234 VGND VGND VPWR VPWR net235 sky130_fd_sc_hd__clkbuf_1
XTAP_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer83 _03595_ VGND VGND VPWR VPWR net330 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer94 _01926_ VGND VGND VPWR VPWR net341 sky130_fd_sc_hd__dlygate4sd1_1
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11660_ _01751_ _01752_ VGND VGND VPWR VPWR _01753_ sky130_fd_sc_hd__nor2_1
XTAP_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10611_ _00173_ _00175_ _04056_ _00563_ VGND VGND VPWR VPWR _00704_ sky130_fd_sc_hd__and4_2
XFILLER_0_138_269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_154_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11591_ _01208_ _01682_ _01683_ VGND VGND VPWR VPWR _01684_ sky130_fd_sc_hd__nand3_2
XFILLER_0_106_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13330_ _09172_ _00218_ _00178_ _09166_ VGND VGND VPWR VPWR _03441_ sky130_fd_sc_hd__a22o_1
X_10542_ _00632_ _00633_ _00450_ _00603_ VGND VGND VPWR VPWR _00635_ sky130_fd_sc_hd__a211o_4
XFILLER_0_92_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13261_ _03352_ _03351_ VGND VGND VPWR VPWR _03365_ sky130_fd_sc_hd__or2b_1
X_10473_ _00564_ _00565_ VGND VGND VPWR VPWR _00566_ sky130_fd_sc_hd__nor2_1
XFILLER_0_106_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15000_ _00189_ _00191_ _07134_ _00309_ VGND VGND VPWR VPWR _05266_ sky130_fd_sc_hd__and4_1
X_12212_ _02151_ _02301_ _02290_ net322 VGND VGND VPWR VPWR _02305_ sky130_fd_sc_hd__a211oi_1
X_13192_ net131 _03266_ _03291_ VGND VGND VPWR VPWR _03293_ sky130_fd_sc_hd__or3_4
XFILLER_0_103_851 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_121_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12143_ _06971_ _03837_ VGND VGND VPWR VPWR _02236_ sky130_fd_sc_hd__nand2_1
XFILLER_0_103_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12074_ _02164_ _02166_ VGND VGND VPWR VPWR _02167_ sky130_fd_sc_hd__and2_1
X_16951_ _07331_ _07338_ VGND VGND VPWR VPWR _07383_ sky130_fd_sc_hd__nand2_1
X_11025_ _01072_ _01074_ _01117_ VGND VGND VPWR VPWR _01118_ sky130_fd_sc_hd__a21oi_1
X_15902_ _05652_ VGND VGND VPWR VPWR _06246_ sky130_fd_sc_hd__buf_2
X_16882_ _07208_ _07211_ _07206_ VGND VGND VPWR VPWR _07309_ sky130_fd_sc_hd__a21bo_1
X_18621_ net267 _09157_ _09171_ _09162_ VGND VGND VPWR VPWR _00031_ sky130_fd_sc_hd__o211a_1
X_15833_ _06112_ _06162_ _06169_ VGND VGND VPWR VPWR _06172_ sky130_fd_sc_hd__nor3_1
XFILLER_0_154_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18552_ net69 VGND VGND VPWR VPWR _09124_ sky130_fd_sc_hd__inv_2
X_15764_ _06095_ _06096_ VGND VGND VPWR VPWR _06097_ sky130_fd_sc_hd__and2_1
XFILLER_0_99_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12976_ _03025_ _03068_ VGND VGND VPWR VPWR _03069_ sky130_fd_sc_hd__and2_1
XFILLER_0_87_635 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17503_ _07868_ _07870_ _07867_ VGND VGND VPWR VPWR _07986_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_59_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14715_ _02975_ _04955_ VGND VGND VPWR VPWR _04956_ sky130_fd_sc_hd__nor2_1
X_11927_ _01952_ _02019_ VGND VGND VPWR VPWR _02020_ sky130_fd_sc_hd__nor2_1
X_18483_ _08978_ _09013_ _09049_ _09012_ _09046_ VGND VGND VPWR VPWR _09050_ sky130_fd_sc_hd__a221o_1
XTAP_2760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15695_ _06017_ _06018_ _06022_ VGND VGND VPWR VPWR _09369_ sky130_fd_sc_hd__o21ai_2
XTAP_2771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_679 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17434_ _03107_ _07355_ _06374_ VGND VGND VPWR VPWR _07911_ sky130_fd_sc_hd__or3b_1
XTAP_2793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14646_ _04867_ _04868_ _04879_ VGND VGND VPWR VPWR _04880_ sky130_fd_sc_hd__a21oi_1
X_11858_ ApproximateM_inst.lob_16.lob2.genblk1\[6\].genblk1.mux.sel ApproximateM_inst.lob_16.lob1.genblk1\[9\].genblk1.mux.sel
+ ApproximateM_inst.lob_16.lob1.genblk1\[8\].genblk1.mux.sel _06008_ VGND VGND VPWR
+ VPWR _01951_ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_19 _01115_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10809_ _00262_ _00901_ VGND VGND VPWR VPWR _00902_ sky130_fd_sc_hd__and2_1
X_17365_ _06764_ _07487_ _07593_ _06653_ VGND VGND VPWR VPWR _07835_ sky130_fd_sc_hd__o22a_1
X_14577_ _04628_ _04698_ _04803_ _04804_ VGND VGND VPWR VPWR _04805_ sky130_fd_sc_hd__o211a_1
X_11789_ _01828_ _01840_ _01836_ _01839_ VGND VGND VPWR VPWR _01882_ sky130_fd_sc_hd__a211o_1
XFILLER_0_138_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16316_ _03199_ _03133_ _06693_ VGND VGND VPWR VPWR _06694_ sky130_fd_sc_hd__a21o_1
X_13528_ _07537_ _00213_ _03655_ _03657_ VGND VGND VPWR VPWR _03658_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_27_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17296_ _07758_ _07759_ VGND VGND VPWR VPWR _07760_ sky130_fd_sc_hd__nor2_1
XFILLER_0_82_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16247_ _03026_ _03052_ _01114_ VGND VGND VPWR VPWR _06619_ sky130_fd_sc_hd__a21o_1
XFILLER_0_140_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_152_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13459_ _03579_ _03581_ _03098_ VGND VGND VPWR VPWR _03582_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput104 net104 VGND VGND VPWR VPWR o_wb_data[29] sky130_fd_sc_hd__clkbuf_4
X_16178_ _06422_ _06459_ VGND VGND VPWR VPWR _06544_ sky130_fd_sc_hd__nor2_1
XFILLER_0_100_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15129_ _05404_ _05406_ VGND VGND VPWR VPWR _05407_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_11_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09621_ _05377_ VGND VGND VPWR VPWR _05388_ sky130_fd_sc_hd__buf_4
XFILLER_0_37_83 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18819_ _09125_ _09323_ VGND VGND VPWR VPWR _09324_ sky130_fd_sc_hd__and2_1
X_09552_ _04493_ VGND VGND VPWR VPWR _04635_ sky130_fd_sc_hd__buf_8
XFILLER_0_78_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09483_ cla_inst.in2\[16\] VGND VGND VPWR VPWR _03881_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_78_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_62 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_512 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_2_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_2_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_104_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09819_ _07526_ VGND VGND VPWR VPWR _07537_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_69_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12830_ _02899_ VGND VGND VPWR VPWR _02923_ sky130_fd_sc_hd__inv_2
XTAP_2001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12761_ _01791_ _01797_ VGND VGND VPWR VPWR _02854_ sky130_fd_sc_hd__nand2_1
XTAP_2056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14500_ _04712_ _04713_ _04718_ VGND VGND VPWR VPWR _04720_ sky130_fd_sc_hd__a21o_1
XTAP_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11712_ _01802_ _01803_ _01776_ _01788_ VGND VGND VPWR VPWR _01805_ sky130_fd_sc_hd__a211o_1
XTAP_2089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15480_ _05786_ _05788_ VGND VGND VPWR VPWR _05789_ sky130_fd_sc_hd__xor2_2
X_12692_ _02783_ _02784_ VGND VGND VPWR VPWR _02785_ sky130_fd_sc_hd__or2_1
XTAP_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14431_ _04643_ _04644_ VGND VGND VPWR VPWR _04645_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_65_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11643_ _01687_ _01688_ _01689_ _01701_ VGND VGND VPWR VPWR _01736_ sky130_fd_sc_hd__a31o_1
XFILLER_0_127_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_139_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17150_ _07598_ _07599_ VGND VGND VPWR VPWR _07600_ sky130_fd_sc_hd__xnor2_2
X_14362_ _03651_ _03662_ _07102_ _05704_ VGND VGND VPWR VPWR _04570_ sky130_fd_sc_hd__nand4_2
X_11574_ _01663_ _01665_ VGND VGND VPWR VPWR _01667_ sky130_fd_sc_hd__or2_1
XFILLER_0_80_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput17 i_wb_addr[23] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__clkbuf_1
Xinput28 i_wb_addr[4] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_91_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16101_ op_code\[2\] op_code\[3\] VGND VGND VPWR VPWR _06459_ sky130_fd_sc_hd__or2_2
Xinput39 i_wb_data[13] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__buf_2
X_13313_ _03419_ _03420_ _03251_ _03252_ VGND VGND VPWR VPWR _03423_ sky130_fd_sc_hd__o211ai_2
X_10525_ _00610_ _00611_ _00616_ VGND VGND VPWR VPWR _00618_ sky130_fd_sc_hd__a21o_1
X_14293_ _00702_ _00443_ _06471_ _00195_ VGND VGND VPWR VPWR _04495_ sky130_fd_sc_hd__a22oi_1
X_17081_ _07523_ _07524_ VGND VGND VPWR VPWR _07525_ sky130_fd_sc_hd__or2_1
X_13244_ _03343_ _03344_ _03346_ VGND VGND VPWR VPWR _03348_ sky130_fd_sc_hd__o21ai_2
X_16032_ _02987_ _01678_ VGND VGND VPWR VPWR _06385_ sky130_fd_sc_hd__or2_1
X_10456_ _00106_ _00206_ VGND VGND VPWR VPWR _00549_ sky130_fd_sc_hd__nand2_1
X_13175_ _00362_ _00878_ _03271_ _03273_ VGND VGND VPWR VPWR _03274_ sky130_fd_sc_hd__a22oi_1
X_10387_ _00477_ _00479_ VGND VGND VPWR VPWR _00480_ sky130_fd_sc_hd__xor2_1
XFILLER_0_103_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12126_ _02181_ _02204_ VGND VGND VPWR VPWR _02219_ sky130_fd_sc_hd__nor2_1
X_17983_ _08447_ _08419_ _08505_ _08508_ VGND VGND VPWR VPWR _08509_ sky130_fd_sc_hd__o31a_1
X_12057_ _02065_ _02147_ _02143_ _02146_ VGND VGND VPWR VPWR _02150_ sky130_fd_sc_hd__a211o_1
X_16934_ _03101_ _06436_ _06424_ VGND VGND VPWR VPWR _07366_ sky130_fd_sc_hd__a21oi_1
X_11008_ _01098_ _01100_ VGND VGND VPWR VPWR _01101_ sky130_fd_sc_hd__xnor2_1
X_16865_ _03324_ _03003_ _06814_ _07289_ VGND VGND VPWR VPWR _07290_ sky130_fd_sc_hd__a211o_2
X_18604_ salida\[20\] _09159_ _09160_ salida\[52\] _09146_ VGND VGND VPWR VPWR _09161_
+ sky130_fd_sc_hd__a221o_1
X_15816_ _03007_ _03067_ VGND VGND VPWR VPWR _06153_ sky130_fd_sc_hd__nand2_1
X_16796_ _07212_ _07214_ VGND VGND VPWR VPWR _07215_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_99_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18535_ net5 net8 net7 net10 VGND VGND VPWR VPWR _09105_ sky130_fd_sc_hd__or4_1
X_15747_ _05795_ _06075_ _06077_ _06078_ VGND VGND VPWR VPWR _06079_ sky130_fd_sc_hd__o211a_1
X_12959_ _01112_ VGND VGND VPWR VPWR _03052_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_59_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18466_ _03913_ _06913_ _08141_ _09031_ _06721_ VGND VGND VPWR VPWR _09032_ sky130_fd_sc_hd__o311a_1
XFILLER_0_8_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15678_ _05957_ _05931_ _06002_ _06003_ VGND VGND VPWR VPWR _06004_ sky130_fd_sc_hd__o211a_1
XTAP_2590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17417_ _07883_ _07890_ VGND VGND VPWR VPWR _07892_ sky130_fd_sc_hd__or2_1
X_14629_ _04852_ _04854_ _04859_ VGND VGND VPWR VPWR _04861_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_90_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18397_ _08955_ _08956_ VGND VGND VPWR VPWR _08957_ sky130_fd_sc_hd__and2_1
XFILLER_0_56_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_362 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17348_ _03198_ _05096_ _06543_ _07809_ _07816_ VGND VGND VPWR VPWR _07817_ sky130_fd_sc_hd__a221o_1
XFILLER_0_114_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_153_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17279_ _02124_ _07592_ VGND VGND VPWR VPWR _07741_ sky130_fd_sc_hd__nand2_4
XFILLER_0_141_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_89 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_592 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19018_ clknet_4_9_0_clk _00003_ VGND VGND VPWR VPWR sel_op\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_139_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09604_ _04733_ _04624_ VGND VGND VPWR VPWR _05203_ sky130_fd_sc_hd__or2b_1
X_09535_ ApproximateM_inst.lob_16.lob1.genblk2.mux_final.sel VGND VGND VPWR VPWR _04449_
+ sky130_fd_sc_hd__buf_6
XFILLER_0_149_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09466_ _03585_ _03640_ _03684_ VGND VGND VPWR VPWR _03695_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_149_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_108_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_354 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10310_ _00203_ _00248_ VGND VGND VPWR VPWR _00403_ sky130_fd_sc_hd__nand2_1
XFILLER_0_132_743 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_771 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_104_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11290_ _01297_ _01298_ VGND VGND VPWR VPWR _01383_ sky130_fd_sc_hd__and2_1
XFILLER_0_120_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10241_ _00303_ _00304_ _08529_ _08659_ VGND VGND VPWR VPWR _00334_ sky130_fd_sc_hd__a211oi_1
X_10172_ _00249_ _00264_ VGND VGND VPWR VPWR _00265_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_100_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14980_ _05009_ _05154_ VGND VGND VPWR VPWR _05244_ sky130_fd_sc_hd__and2b_1
X_13931_ _03933_ _03934_ VGND VGND VPWR VPWR _04098_ sky130_fd_sc_hd__nand2_1
X_16650_ _06749_ _06969_ VGND VGND VPWR VPWR _07056_ sky130_fd_sc_hd__nand2_1
X_13862_ _04021_ _04022_ VGND VGND VPWR VPWR _04024_ sky130_fd_sc_hd__xor2_2
XFILLER_0_88_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15601_ _05918_ _05919_ VGND VGND VPWR VPWR _05920_ sky130_fd_sc_hd__and2_1
X_12813_ _00854_ _02898_ _01465_ _01466_ VGND VGND VPWR VPWR _02906_ sky130_fd_sc_hd__o211ai_1
X_16581_ _06934_ _06935_ _06980_ VGND VGND VPWR VPWR _06981_ sky130_fd_sc_hd__o21ba_1
X_13793_ _03762_ _03767_ _03761_ VGND VGND VPWR VPWR _03948_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_69_465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18320_ _08872_ _08840_ _08841_ VGND VGND VPWR VPWR _08874_ sky130_fd_sc_hd__and3_1
X_15532_ _05737_ _05755_ _05844_ VGND VGND VPWR VPWR _05846_ sky130_fd_sc_hd__o21ai_2
XTAP_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12744_ _02634_ _02668_ VGND VGND VPWR VPWR _02837_ sky130_fd_sc_hd__xnor2_1
XTAP_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18251_ _08730_ _08729_ VGND VGND VPWR VPWR _08799_ sky130_fd_sc_hd__or2b_1
X_15463_ _05688_ _05770_ VGND VGND VPWR VPWR _05771_ sky130_fd_sc_hd__nand2_1
XTAP_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12675_ _02766_ _02767_ VGND VGND VPWR VPWR _02768_ sky130_fd_sc_hd__nor2_1
XFILLER_0_53_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17202_ _06750_ _07650_ _07656_ VGND VGND VPWR VPWR _07658_ sky130_fd_sc_hd__and3_1
XFILLER_0_25_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14414_ _04608_ _04609_ _04625_ VGND VGND VPWR VPWR _04627_ sky130_fd_sc_hd__a21oi_1
X_11626_ _01710_ _01716_ _01717_ _01718_ VGND VGND VPWR VPWR _01719_ sky130_fd_sc_hd__nand4_2
X_18182_ _08715_ _08723_ VGND VGND VPWR VPWR _08725_ sky130_fd_sc_hd__and2_1
X_15394_ _05694_ _05695_ VGND VGND VPWR VPWR _05696_ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17133_ _06462_ _07574_ _07576_ _07582_ VGND VGND VPWR VPWR _07583_ sky130_fd_sc_hd__or4_1
X_14345_ _04550_ _04551_ VGND VGND VPWR VPWR _04552_ sky130_fd_sc_hd__or2_1
XFILLER_0_80_652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11557_ _05682_ _03750_ _01597_ _01596_ _04143_ VGND VGND VPWR VPWR _01650_ sky130_fd_sc_hd__a32o_1
XFILLER_0_52_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10508_ _00291_ _00431_ _00465_ _00466_ VGND VGND VPWR VPWR _00601_ sky130_fd_sc_hd__o211a_1
X_17064_ _07484_ _07506_ VGND VGND VPWR VPWR _07507_ sky130_fd_sc_hd__xor2_1
X_14276_ _07504_ _04012_ _04045_ _00358_ VGND VGND VPWR VPWR _04476_ sky130_fd_sc_hd__a22o_1
X_11488_ _01573_ _01574_ _01580_ VGND VGND VPWR VPWR _01581_ sky130_fd_sc_hd__nand3_2
XFILLER_0_123_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16015_ _02347_ _00558_ VGND VGND VPWR VPWR _06366_ sky130_fd_sc_hd__and2_1
X_10439_ _00529_ _00530_ _00349_ _00531_ VGND VGND VPWR VPWR _00532_ sky130_fd_sc_hd__o211ai_4
X_13227_ _03319_ _03329_ VGND VGND VPWR VPWR _03330_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_100_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13158_ _03247_ _03254_ _03255_ VGND VGND VPWR VPWR _03256_ sky130_fd_sc_hd__nand3_4
XTAP_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12109_ _02140_ _02201_ VGND VGND VPWR VPWR _02202_ sky130_fd_sc_hd__and2_1
X_13089_ _02505_ _02259_ VGND VGND VPWR VPWR _03181_ sky130_fd_sc_hd__nor2_1
X_17966_ _08487_ _08488_ _08489_ VGND VGND VPWR VPWR _08490_ sky130_fd_sc_hd__and3_1
XTAP_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16917_ _07345_ _07346_ VGND VGND VPWR VPWR _07347_ sky130_fd_sc_hd__nor2_1
X_17897_ _08016_ _08121_ _08414_ VGND VGND VPWR VPWR _08415_ sky130_fd_sc_hd__or3_1
XFILLER_0_79_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16848_ _06424_ _06436_ VGND VGND VPWR VPWR _07272_ sky130_fd_sc_hd__nor2_1
XFILLER_0_19_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16779_ _06563_ _07195_ VGND VGND VPWR VPWR _07196_ sky130_fd_sc_hd__nor2_1
X_18518_ _06680_ _09086_ VGND VGND VPWR VPWR _09087_ sky130_fd_sc_hd__nor2_1
XFILLER_0_29_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18449_ _09011_ _09012_ VGND VGND VPWR VPWR _09013_ sky130_fd_sc_hd__and2b_1
XFILLER_0_7_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_141_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_384 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_114_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_538 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_149_640 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09518_ net227 net169 _03421_ _04242_ VGND VGND VPWR VPWR _04263_ sky130_fd_sc_hd__nand4_2
X_10790_ _00882_ _00208_ VGND VGND VPWR VPWR _00883_ sky130_fd_sc_hd__xnor2_1
XPHY_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09449_ _03498_ VGND VGND VPWR VPWR _03509_ sky130_fd_sc_hd__buf_6
XPHY_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12460_ _06971_ _00177_ _02551_ _02552_ VGND VGND VPWR VPWR _02553_ sky130_fd_sc_hd__nand4_2
XFILLER_0_47_693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11411_ _00170_ VGND VGND VPWR VPWR _01504_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_105_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12391_ _02482_ _02483_ VGND VGND VPWR VPWR _02484_ sky130_fd_sc_hd__xor2_1
XFILLER_0_151_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14130_ _04313_ _04314_ _04123_ _04145_ VGND VGND VPWR VPWR _04316_ sky130_fd_sc_hd__a211oi_4
X_11342_ _01421_ _01433_ VGND VGND VPWR VPWR _01435_ sky130_fd_sc_hd__nor2_1
XFILLER_0_104_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_590 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11273_ _01267_ _01365_ VGND VGND VPWR VPWR _01366_ sky130_fd_sc_hd__xnor2_1
X_14061_ _03913_ VGND VGND VPWR VPWR _04241_ sky130_fd_sc_hd__buf_4
XFILLER_0_120_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10224_ _06051_ _07156_ _07134_ _06040_ VGND VGND VPWR VPWR _00317_ sky130_fd_sc_hd__a22o_1
X_13012_ _02373_ _03104_ _03040_ VGND VGND VPWR VPWR _03105_ sky130_fd_sc_hd__o21ai_2
X_17820_ _08231_ _08233_ _08230_ VGND VGND VPWR VPWR _08331_ sky130_fd_sc_hd__a21boi_2
X_10155_ _00247_ VGND VGND VPWR VPWR _00248_ sky130_fd_sc_hd__clkbuf_4
X_17751_ _08185_ _08201_ VGND VGND VPWR VPWR _08255_ sky130_fd_sc_hd__nor2_1
X_14963_ _05119_ _05223_ _05225_ VGND VGND VPWR VPWR _05226_ sky130_fd_sc_hd__and3_1
XFILLER_0_55_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10086_ ApproximateM_inst.lob_16.lob1.genblk1\[4\].genblk1.mux.sel VGND VGND VPWR
+ VPWR _00179_ sky130_fd_sc_hd__buf_4
XFILLER_0_89_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16702_ _06567_ _06570_ _00357_ VGND VGND VPWR VPWR _07113_ sky130_fd_sc_hd__o21a_1
X_13914_ _03177_ VGND VGND VPWR VPWR _04081_ sky130_fd_sc_hd__inv_2
X_17682_ _08172_ _08179_ VGND VGND VPWR VPWR _08181_ sky130_fd_sc_hd__xnor2_1
X_14894_ _05144_ _05149_ _05150_ VGND VGND VPWR VPWR _05151_ sky130_fd_sc_hd__and3_1
X_16633_ _06807_ VGND VGND VPWR VPWR _07038_ sky130_fd_sc_hd__clkbuf_4
X_13845_ _04002_ _04003_ _03811_ _03833_ VGND VGND VPWR VPWR _04005_ sky130_fd_sc_hd__o211a_1
X_16564_ _06959_ _06962_ VGND VGND VPWR VPWR _06963_ sky130_fd_sc_hd__xnor2_1
X_13776_ _03904_ _03905_ _03929_ VGND VGND VPWR VPWR _09380_ sky130_fd_sc_hd__o21ai_2
X_10988_ ApproximateM_inst.lob_16.lob2.genblk1\[3\].genblk1.mux.sel VGND VGND VPWR
+ VPWR _01081_ sky130_fd_sc_hd__buf_4
XFILLER_0_84_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18303_ _08853_ _08855_ VGND VGND VPWR VPWR _08856_ sky130_fd_sc_hd__and2_1
XFILLER_0_128_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15515_ _05825_ _05826_ VGND VGND VPWR VPWR _05827_ sky130_fd_sc_hd__nor2_1
X_12727_ _02803_ _02819_ VGND VGND VPWR VPWR _02820_ sky130_fd_sc_hd__nor2_1
X_16495_ _06867_ _06887_ VGND VGND VPWR VPWR _06888_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_26_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18234_ _08776_ _08780_ VGND VGND VPWR VPWR _08781_ sky130_fd_sc_hd__nor2_1
XFILLER_0_38_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15446_ _05740_ _05662_ _05751_ VGND VGND VPWR VPWR _05752_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_72_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12658_ _02746_ _02750_ VGND VGND VPWR VPWR _02751_ sky130_fd_sc_hd__xor2_1
XFILLER_0_53_630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11609_ _01585_ _01602_ _01700_ _01701_ VGND VGND VPWR VPWR _01702_ sky130_fd_sc_hd__a211oi_2
X_18165_ _07665_ _07708_ _08150_ _07216_ VGND VGND VPWR VPWR _08706_ sky130_fd_sc_hd__a22o_1
X_15377_ _03006_ _04336_ VGND VGND VPWR VPWR _05677_ sky130_fd_sc_hd__nand2_1
XFILLER_0_154_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12589_ _02597_ _02640_ _02639_ VGND VGND VPWR VPWR _02682_ sky130_fd_sc_hd__a21o_1
XFILLER_0_111_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17116_ _07562_ _03930_ _07563_ VGND VGND VPWR VPWR _07564_ sky130_fd_sc_hd__and3_1
X_14328_ _04492_ _04531_ _04532_ VGND VGND VPWR VPWR _04533_ sky130_fd_sc_hd__or3_4
XFILLER_0_4_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18096_ _08629_ _08630_ VGND VGND VPWR VPWR _08631_ sky130_fd_sc_hd__nand2_1
XFILLER_0_80_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_cap125 _01707_ VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__clkbuf_2
Xmax_cap147 _07023_ VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__buf_1
X_17047_ _06563_ _06572_ _07387_ _07487_ VGND VGND VPWR VPWR _07488_ sky130_fd_sc_hd__or4_2
X_14259_ _04445_ _04446_ _04456_ VGND VGND VPWR VPWR _04457_ sky130_fd_sc_hd__o21a_1
XFILLER_0_0_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_96_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18998_ clknet_4_7_0_clk _09364_ VGND VGND VPWR VPWR salida\[51\] sky130_fd_sc_hd__dfxtp_1
XTAP_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17949_ _08353_ _08355_ VGND VGND VPWR VPWR _08471_ sky130_fd_sc_hd__or2_1
XFILLER_0_136_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09998_ _09339_ _09340_ _07482_ _07908_ VGND VGND VPWR VPWR _09341_ sky130_fd_sc_hd__o211a_1
XFILLER_0_98_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11960_ _02027_ _02052_ _01967_ VGND VGND VPWR VPWR _02053_ sky130_fd_sc_hd__o21ai_2
X_10911_ _01000_ _01003_ VGND VGND VPWR VPWR _01004_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_98_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11891_ _01979_ _01982_ _01983_ VGND VGND VPWR VPWR _01984_ sky130_fd_sc_hd__or3_4
X_13630_ _03761_ _03762_ _03767_ VGND VGND VPWR VPWR _03769_ sky130_fd_sc_hd__a21o_1
X_10842_ net169 _00179_ ApproximateM_inst.lob_16.lob1.genblk1\[2\].genblk1.mux.sel
+ net227 VGND VGND VPWR VPWR _00935_ sky130_fd_sc_hd__a22o_1
X_13561_ _00164_ _03693_ VGND VGND VPWR VPWR _03694_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10773_ _00118_ _00865_ VGND VGND VPWR VPWR _00866_ sky130_fd_sc_hd__nor2_1
XFILLER_0_94_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15300_ _05574_ _05592_ VGND VGND VPWR VPWR _05593_ sky130_fd_sc_hd__nor2_1
XFILLER_0_81_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12512_ _02556_ _02594_ _02603_ VGND VGND VPWR VPWR _02605_ sky130_fd_sc_hd__and3_1
X_16280_ _06561_ _06572_ _06579_ _06653_ VGND VGND VPWR VPWR _06654_ sky130_fd_sc_hd__or4_1
X_13492_ _03609_ _03617_ VGND VGND VPWR VPWR _03619_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_19_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_136_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_124_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15231_ _05516_ _05517_ VGND VGND VPWR VPWR _05518_ sky130_fd_sc_hd__or2b_1
X_12443_ _00357_ _02487_ _02486_ VGND VGND VPWR VPWR _02536_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_81_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_679 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15162_ _05432_ _05441_ VGND VGND VPWR VPWR _05443_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_34_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12374_ _02398_ _02465_ _02466_ VGND VGND VPWR VPWR _02467_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_105_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_151_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14113_ _04283_ net133 _04295_ VGND VGND VPWR VPWR _04298_ sky130_fd_sc_hd__or3_1
X_11325_ _01356_ _07646_ _09354_ _01417_ VGND VGND VPWR VPWR _01418_ sky130_fd_sc_hd__a22oi_1
X_15093_ _00189_ _07134_ VGND VGND VPWR VPWR _05368_ sky130_fd_sc_hd__and2_1
X_14044_ net319 _04219_ _04221_ VGND VGND VPWR VPWR _04223_ sky130_fd_sc_hd__o21a_1
X_11256_ _01347_ _01348_ VGND VGND VPWR VPWR _01349_ sky130_fd_sc_hd__nor2_1
X_18921_ clknet_4_13_0_clk _00075_ VGND VGND VPWR VPWR ApproximateM_inst.lob_16.lob2.genblk1\[7\].genblk1.mux.sel
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_120_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10207_ _08615_ _05856_ _08572_ _08561_ VGND VGND VPWR VPWR _00300_ sky130_fd_sc_hd__a31o_1
X_11187_ _00969_ _00971_ _00970_ VGND VGND VPWR VPWR _01280_ sky130_fd_sc_hd__o21ba_1
X_18852_ clknet_4_6_0_clk net286 VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__dfxtp_1
X_17803_ _08294_ _08312_ VGND VGND VPWR VPWR _08313_ sky130_fd_sc_hd__xor2_1
X_10138_ _00162_ _00230_ VGND VGND VPWR VPWR _00231_ sky130_fd_sc_hd__nand2_2
X_18783_ _02987_ net44 _09276_ VGND VGND VPWR VPWR _09296_ sky130_fd_sc_hd__mux2_1
X_15995_ _05747_ _00223_ VGND VGND VPWR VPWR _06344_ sky130_fd_sc_hd__nand2_1
X_17734_ _03588_ _06385_ _06383_ VGND VGND VPWR VPWR _08238_ sky130_fd_sc_hd__a21o_1
X_14946_ _05173_ _05174_ VGND VGND VPWR VPWR _05207_ sky130_fd_sc_hd__or2b_1
X_10069_ _00160_ _00141_ VGND VGND VPWR VPWR _00162_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_89_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17665_ _08160_ _08161_ VGND VGND VPWR VPWR _08162_ sky130_fd_sc_hd__nand2_1
X_14877_ _05124_ _05131_ VGND VGND VPWR VPWR _05132_ sky130_fd_sc_hd__or2_1
X_16616_ _06937_ _07018_ VGND VGND VPWR VPWR _07019_ sky130_fd_sc_hd__or2_1
X_13828_ cla_inst.in2\[31\] _00207_ VGND VGND VPWR VPWR _03986_ sky130_fd_sc_hd__nand2_1
X_17596_ _07038_ _07623_ VGND VGND VPWR VPWR _08087_ sky130_fd_sc_hd__nand2_1
XFILLER_0_106_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16547_ _06942_ _06943_ _06084_ VGND VGND VPWR VPWR _06944_ sky130_fd_sc_hd__a21bo_2
X_13759_ _03909_ _03910_ _02981_ VGND VGND VPWR VPWR _03911_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16478_ _03003_ _03004_ _06523_ VGND VGND VPWR VPWR _06869_ sky130_fd_sc_hd__or3_1
XFILLER_0_143_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18217_ _02994_ _04900_ VGND VGND VPWR VPWR _08763_ sky130_fd_sc_hd__nand2_1
XFILLER_0_122_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15429_ _05685_ _05732_ VGND VGND VPWR VPWR _05733_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_72_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18148_ _02997_ _06593_ _06594_ VGND VGND VPWR VPWR _08688_ sky130_fd_sc_hd__a21o_1
XFILLER_0_13_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_124_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18079_ _06421_ _08597_ _08598_ _08606_ _08612_ VGND VGND VPWR VPWR _08613_ sky130_fd_sc_hd__a311o_1
XFILLER_0_111_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09921_ _08496_ _08507_ _08518_ VGND VGND VPWR VPWR _08648_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_1_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09852_ _07482_ _07493_ _07886_ VGND VGND VPWR VPWR _07897_ sky130_fd_sc_hd__a21bo_1
XTAP_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09783_ _07058_ _07091_ _07123_ _07134_ VGND VGND VPWR VPWR _07145_ sky130_fd_sc_hd__nand4_2
XTAP_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_109 net42 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_755 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_799 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_119_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11110_ _01074_ _01075_ _01202_ _01053_ VGND VGND VPWR VPWR _01203_ sky130_fd_sc_hd__o2bb2a_1
X_12090_ _02177_ _02182_ VGND VGND VPWR VPWR _02183_ sky130_fd_sc_hd__nand2_1
X_11041_ _01121_ _01133_ VGND VGND VPWR VPWR _01134_ sky130_fd_sc_hd__or2_1
X_14800_ _02999_ _04900_ VGND VGND VPWR VPWR _05048_ sky130_fd_sc_hd__nand2_1
X_15780_ _06043_ _06036_ VGND VGND VPWR VPWR _06114_ sky130_fd_sc_hd__and2b_1
XFILLER_0_98_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12992_ _03024_ _03084_ VGND VGND VPWR VPWR _03085_ sky130_fd_sc_hd__nand2_1
XFILLER_0_99_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14731_ _02986_ _07384_ _04970_ _04971_ VGND VGND VPWR VPWR _04972_ sky130_fd_sc_hd__and4_1
X_11943_ _00832_ _04886_ VGND VGND VPWR VPWR _02036_ sky130_fd_sc_hd__nand2_1
XFILLER_0_87_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17450_ _06836_ _07913_ _07915_ _07927_ VGND VGND VPWR VPWR _07928_ sky130_fd_sc_hd__o31a_1
X_14662_ _04885_ _04768_ _04895_ VGND VGND VPWR VPWR _04898_ sky130_fd_sc_hd__and3_1
X_11874_ _01864_ _01964_ VGND VGND VPWR VPWR _01967_ sky130_fd_sc_hd__and2_1
XFILLER_0_79_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16401_ _06337_ _06336_ _06335_ VGND VGND VPWR VPWR _06786_ sky130_fd_sc_hd__a21oi_1
X_13613_ _03649_ _03650_ _03670_ VGND VGND VPWR VPWR _03751_ sky130_fd_sc_hd__nor3_1
X_17381_ _07822_ _07729_ _07850_ VGND VGND VPWR VPWR _07852_ sky130_fd_sc_hd__and3_1
X_10825_ _00912_ _00913_ _00917_ VGND VGND VPWR VPWR _00918_ sky130_fd_sc_hd__and3_1
X_14593_ _03930_ VGND VGND VPWR VPWR _04823_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_94_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16332_ _03916_ _06710_ VGND VGND VPWR VPWR _06712_ sky130_fd_sc_hd__and2_1
X_13544_ _03438_ _03463_ VGND VGND VPWR VPWR _03676_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10756_ _00831_ _00844_ VGND VGND VPWR VPWR _00849_ sky130_fd_sc_hd__xor2_1
XFILLER_0_82_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16263_ _03026_ _03108_ _01963_ VGND VGND VPWR VPWR _06637_ sky130_fd_sc_hd__a21o_1
X_13475_ _03598_ _03599_ VGND VGND VPWR VPWR _03600_ sky130_fd_sc_hd__nand2_1
XFILLER_0_54_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10687_ _04668_ _04679_ _04711_ VGND VGND VPWR VPWR _00780_ sky130_fd_sc_hd__o21ai_1
X_18002_ _08509_ _08511_ _08528_ _06723_ _00813_ VGND VGND VPWR VPWR _09399_ sky130_fd_sc_hd__o32a_1
X_15214_ _05460_ _05384_ _05498_ VGND VGND VPWR VPWR _05500_ sky130_fd_sc_hd__nand3_1
XFILLER_0_124_145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12426_ _02439_ _02518_ VGND VGND VPWR VPWR _02519_ sky130_fd_sc_hd__xnor2_1
X_16194_ net334 VGND VGND VPWR VPWR _06561_ sky130_fd_sc_hd__buf_2
XFILLER_0_106_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15145_ _04823_ _05417_ _05418_ _05424_ VGND VGND VPWR VPWR _09361_ sky130_fd_sc_hd__a31o_1
X_12357_ _02416_ _02448_ net128 _02449_ VGND VGND VPWR VPWR _02450_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_121_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11308_ _01399_ _01400_ VGND VGND VPWR VPWR _01401_ sky130_fd_sc_hd__or2_1
X_15076_ _05258_ _05256_ VGND VGND VPWR VPWR _05349_ sky130_fd_sc_hd__and2b_1
X_12288_ _02378_ _02379_ _02368_ _02376_ VGND VGND VPWR VPWR _02381_ sky130_fd_sc_hd__o211a_1
X_14027_ _04197_ _04203_ VGND VGND VPWR VPWR _04204_ sky130_fd_sc_hd__xnor2_1
X_18904_ clknet_4_10_0_clk _00058_ VGND VGND VPWR VPWR cla_inst.in1\[22\] sky130_fd_sc_hd__dfxtp_4
X_11239_ _01313_ _01314_ _01330_ _01331_ VGND VGND VPWR VPWR _01332_ sky130_fd_sc_hd__a211o_2
X_18835_ _09335_ VGND VGND VPWR VPWR _00103_ sky130_fd_sc_hd__clkbuf_1
X_18766_ _09273_ _09282_ VGND VGND VPWR VPWR _09283_ sky130_fd_sc_hd__and2_1
X_15978_ _06323_ _06324_ _06325_ _03039_ VGND VGND VPWR VPWR _09378_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_117_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17717_ _08014_ _08119_ VGND VGND VPWR VPWR _08219_ sky130_fd_sc_hd__nor2_1
X_14929_ _05065_ _05067_ _05187_ VGND VGND VPWR VPWR _05189_ sky130_fd_sc_hd__nand3_1
XFILLER_0_78_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18697_ _01136_ _09183_ net69 VGND VGND VPWR VPWR _09229_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_78_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17648_ _06630_ _08141_ _08143_ _06720_ VGND VGND VPWR VPWR _08144_ sky130_fd_sc_hd__o211a_1
XFILLER_0_148_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17579_ _07751_ _07394_ _07604_ _07039_ VGND VGND VPWR VPWR _08068_ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_739 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_216 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_116_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_307 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09904_ _03728_ _08452_ VGND VGND VPWR VPWR _08463_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09835_ _07700_ VGND VGND VPWR VPWR _07711_ sky130_fd_sc_hd__clkbuf_4
XTAP_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09766_ _05943_ _06138_ _05812_ _05823_ VGND VGND VPWR VPWR _06960_ sky130_fd_sc_hd__a211oi_2
XTAP_2205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09697_ _03465_ _03914_ VGND VGND VPWR VPWR _06213_ sky130_fd_sc_hd__and2_1
XTAP_2216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer40 _02693_ VGND VGND VPWR VPWR net203 sky130_fd_sc_hd__buf_1
XTAP_2227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer51 _00956_ VGND VGND VPWR VPWR net214 sky130_fd_sc_hd__clkbuf_1
XTAP_2238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer62 _03590_ VGND VGND VPWR VPWR net225 sky130_fd_sc_hd__buf_6
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer73 _03772_ VGND VGND VPWR VPWR net236 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xrebuffer95 _04549_ VGND VGND VPWR VPWR net342 sky130_fd_sc_hd__buf_6
XTAP_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10610_ _00702_ _04154_ _00165_ _00195_ VGND VGND VPWR VPWR _00703_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_64_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11590_ _06982_ _00443_ _01206_ _01207_ VGND VGND VPWR VPWR _01683_ sky130_fd_sc_hd__a22o_1
XFILLER_0_25_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10541_ _00450_ net143 _00632_ _00633_ VGND VGND VPWR VPWR _00634_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_24_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13260_ _03125_ _03133_ _03196_ _03199_ _03364_ VGND VGND VPWR VPWR _09366_ sky130_fd_sc_hd__a221o_1
X_10472_ _00173_ _00183_ _03673_ _00211_ VGND VGND VPWR VPWR _00565_ sky130_fd_sc_hd__and4_1
X_12211_ _02131_ _02303_ VGND VGND VPWR VPWR _02304_ sky130_fd_sc_hd__xor2_1
XFILLER_0_32_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13191_ _03267_ _03290_ VGND VGND VPWR VPWR _03291_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_32_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_863 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12142_ _02211_ _02213_ VGND VGND VPWR VPWR _02235_ sky130_fd_sc_hd__nor2_1
X_12073_ _02165_ _02080_ VGND VGND VPWR VPWR _02166_ sky130_fd_sc_hd__xnor2_2
X_16950_ _07328_ _07329_ VGND VGND VPWR VPWR _07382_ sky130_fd_sc_hd__or2b_1
X_11024_ _01104_ _01116_ VGND VGND VPWR VPWR _01117_ sky130_fd_sc_hd__xnor2_1
X_15901_ _06242_ _06243_ VGND VGND VPWR VPWR _06244_ sky130_fd_sc_hd__and2_1
X_16881_ _07305_ _07306_ VGND VGND VPWR VPWR _07307_ sky130_fd_sc_hd__xnor2_1
X_15832_ _06112_ _06162_ _06169_ VGND VGND VPWR VPWR _06171_ sky130_fd_sc_hd__o21a_1
X_18620_ salida\[27\] _09159_ _09160_ salida\[59\] _09163_ VGND VGND VPWR VPWR _09171_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_99_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15763_ _06088_ _06093_ VGND VGND VPWR VPWR _06096_ sky130_fd_sc_hd__nand2_1
X_18551_ salida\[0\] _09114_ _09118_ salida\[32\] _09121_ VGND VGND VPWR VPWR _09122_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_63_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12975_ _03067_ VGND VGND VPWR VPWR _03068_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_59_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14714_ _03562_ _03577_ _03079_ VGND VGND VPWR VPWR _04955_ sky130_fd_sc_hd__mux2_1
X_17502_ _07982_ _07983_ VGND VGND VPWR VPWR _07985_ sky130_fd_sc_hd__xnor2_1
X_11926_ _06711_ _04067_ _02018_ _01951_ VGND VGND VPWR VPWR _02019_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_87_647 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18482_ _08969_ _09011_ VGND VGND VPWR VPWR _09049_ sky130_fd_sc_hd__or2_1
XTAP_2750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15694_ _03547_ _04249_ _05307_ _06021_ _03039_ VGND VGND VPWR VPWR _06022_ sky130_fd_sc_hd__o32a_1
XTAP_2761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17433_ _06374_ _06511_ _02044_ VGND VGND VPWR VPWR _07910_ sky130_fd_sc_hd__a21oi_1
XTAP_2783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14645_ _04877_ _04878_ VGND VGND VPWR VPWR _04879_ sky130_fd_sc_hd__and2_1
XTAP_2794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11857_ _06008_ ApproximateM_inst.lob_16.lob2.genblk1\[6\].genblk1.mux.sel ApproximateM_inst.lob_16.lob1.genblk1\[9\].genblk1.mux.sel
+ ApproximateM_inst.lob_16.lob1.genblk1\[8\].genblk1.mux.sel VGND VGND VPWR VPWR _01950_
+ sky130_fd_sc_hd__and4_1
XFILLER_0_129_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10808_ _00249_ _00264_ VGND VGND VPWR VPWR _00901_ sky130_fd_sc_hd__or2b_1
X_17364_ _06655_ _06762_ _07489_ _07596_ VGND VGND VPWR VPWR _07834_ sky130_fd_sc_hd__and4_1
X_14576_ _04758_ _04759_ _04801_ _04802_ VGND VGND VPWR VPWR _04804_ sky130_fd_sc_hd__a22o_1
XFILLER_0_82_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11788_ _01540_ _01879_ _01880_ VGND VGND VPWR VPWR _01881_ sky130_fd_sc_hd__nand3_2
XFILLER_0_103_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16315_ _06508_ _06676_ _06677_ _06692_ VGND VGND VPWR VPWR _06693_ sky130_fd_sc_hd__a31o_1
XFILLER_0_138_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13527_ _03654_ VGND VGND VPWR VPWR _03657_ sky130_fd_sc_hd__inv_2
X_10739_ ApproximateM_inst.lob_16.lob2.genblk1\[2\].genblk1.mux.sel VGND VGND VPWR
+ VPWR _00832_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_82_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17295_ _07756_ _07757_ VGND VGND VPWR VPWR _07759_ sky130_fd_sc_hd__and2_1
XFILLER_0_153_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16246_ _03027_ _03044_ _01224_ VGND VGND VPWR VPWR _06618_ sky130_fd_sc_hd__a21o_1
XFILLER_0_153_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13458_ _03090_ _03189_ _03580_ VGND VGND VPWR VPWR _03581_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_70_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_140_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12409_ _01105_ _00514_ _02099_ _00212_ VGND VGND VPWR VPWR _02502_ sky130_fd_sc_hd__or4b_4
XFILLER_0_2_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16177_ _06418_ _06422_ VGND VGND VPWR VPWR _06543_ sky130_fd_sc_hd__nor2_4
X_13389_ _03494_ _03505_ VGND VGND VPWR VPWR _03506_ sky130_fd_sc_hd__xnor2_1
Xoutput105 net105 VGND VGND VPWR VPWR o_wb_data[2] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_88_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15128_ _05405_ _05296_ VGND VGND VPWR VPWR _05406_ sky130_fd_sc_hd__or2_2
XFILLER_0_121_660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15059_ _05223_ _05329_ VGND VGND VPWR VPWR _05330_ sky130_fd_sc_hd__xor2_1
XFILLER_0_49_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09620_ cla_inst.in1\[18\] VGND VGND VPWR VPWR _05377_ sky130_fd_sc_hd__buf_6
X_18818_ _03013_ net56 _09301_ VGND VGND VPWR VPWR _09323_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09551_ _04329_ _04613_ VGND VGND VPWR VPWR _04624_ sky130_fd_sc_hd__xnor2_2
X_18749_ _09245_ _09268_ VGND VGND VPWR VPWR _09269_ sky130_fd_sc_hd__and2_1
XFILLER_0_77_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09482_ _03793_ _03815_ _03837_ _03859_ VGND VGND VPWR VPWR _03870_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_77_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_850 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_148_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_680 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_224 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_135_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_131_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09818_ cla_inst.in2\[28\] VGND VGND VPWR VPWR _07526_ sky130_fd_sc_hd__buf_2
X_09749_ _06732_ VGND VGND VPWR VPWR _06776_ sky130_fd_sc_hd__inv_4
XTAP_2002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12760_ _00591_ _01248_ _01247_ _02852_ VGND VGND VPWR VPWR _02853_ sky130_fd_sc_hd__a31o_2
XTAP_2035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11711_ _01776_ _01788_ _01802_ net210 VGND VGND VPWR VPWR _01804_ sky130_fd_sc_hd__o211ai_2
XTAP_2079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12691_ _07788_ _07570_ VGND VGND VPWR VPWR _02784_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_568 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14430_ _04503_ _04505_ _04502_ VGND VGND VPWR VPWR _04644_ sky130_fd_sc_hd__o21ai_4
XTAP_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11642_ _01733_ _01734_ VGND VGND VPWR VPWR _01735_ sky130_fd_sc_hd__or2_1
XFILLER_0_25_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14361_ _03377_ _07102_ _05693_ _03356_ VGND VGND VPWR VPWR _04568_ sky130_fd_sc_hd__a22o_1
XFILLER_0_119_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11573_ _01663_ _01665_ VGND VGND VPWR VPWR _01666_ sky130_fd_sc_hd__xor2_1
XFILLER_0_135_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_739 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput18 i_wb_addr[24] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__clkbuf_1
X_16100_ _06326_ _04823_ _06327_ _06458_ VGND VGND VPWR VPWR _09418_ sky130_fd_sc_hd__a31o_1
XFILLER_0_92_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13312_ _03251_ _03252_ _03419_ _03420_ VGND VGND VPWR VPWR _03422_ sky130_fd_sc_hd__a211o_2
Xinput29 i_wb_addr[5] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__clkbuf_1
X_10524_ _00610_ _00611_ _00616_ VGND VGND VPWR VPWR _00617_ sky130_fd_sc_hd__nand3_1
X_17080_ _07419_ _07420_ _07416_ VGND VGND VPWR VPWR _07524_ sky130_fd_sc_hd__o21a_1
X_14292_ _04345_ _04344_ VGND VGND VPWR VPWR _04494_ sky130_fd_sc_hd__or2b_1
XFILLER_0_80_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16031_ _06380_ _06381_ _06382_ VGND VGND VPWR VPWR _06383_ sky130_fd_sc_hd__a21bo_1
X_13243_ _03343_ _03344_ _03346_ VGND VGND VPWR VPWR _03347_ sky130_fd_sc_hd__or3_4
XFILLER_0_122_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10455_ _00546_ _00547_ VGND VGND VPWR VPWR _00548_ sky130_fd_sc_hd__nor2_1
XFILLER_0_33_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13174_ _03270_ VGND VGND VPWR VPWR _03273_ sky130_fd_sc_hd__inv_2
X_10386_ _08158_ _00319_ _00478_ VGND VGND VPWR VPWR _00479_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_0_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12125_ _02213_ _02217_ VGND VGND VPWR VPWR _02218_ sky130_fd_sc_hd__nor2_1
X_17982_ _06559_ _08506_ VGND VGND VPWR VPWR _08508_ sky130_fd_sc_hd__nor2_1
XFILLER_0_102_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12056_ _02107_ _02133_ _02122_ _02132_ VGND VGND VPWR VPWR _02149_ sky130_fd_sc_hd__o211a_1
X_16933_ _06361_ _06359_ _06360_ _06598_ _07364_ VGND VGND VPWR VPWR _07365_ sky130_fd_sc_hd__a311oi_1
X_11007_ _01084_ _01099_ VGND VGND VPWR VPWR _01100_ sky130_fd_sc_hd__and2b_1
X_16864_ _05453_ VGND VGND VPWR VPWR _07289_ sky130_fd_sc_hd__inv_2
X_18603_ _09117_ VGND VGND VPWR VPWR _09160_ sky130_fd_sc_hd__clkbuf_4
X_15815_ _03537_ _04560_ _06151_ VGND VGND VPWR VPWR _06152_ sky130_fd_sc_hd__a21o_1
X_16795_ _06766_ _06875_ _07116_ _07213_ VGND VGND VPWR VPWR _07214_ sky130_fd_sc_hd__o31a_1
XFILLER_0_59_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18534_ net29 net31 net30 net33 VGND VGND VPWR VPWR _09104_ sky130_fd_sc_hd__or4_2
X_15746_ _05945_ _06013_ _06014_ VGND VGND VPWR VPWR _06078_ sky130_fd_sc_hd__o21ba_1
X_12958_ _03043_ _03046_ _03050_ VGND VGND VPWR VPWR _03051_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11909_ _04362_ _01031_ _09179_ _04340_ VGND VGND VPWR VPWR _02002_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_90_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15677_ _06000_ _06001_ _05968_ VGND VGND VPWR VPWR _06003_ sky130_fd_sc_hd__a21o_1
X_18465_ _06411_ _06546_ _09030_ _03073_ VGND VGND VPWR VPWR _09031_ sky130_fd_sc_hd__a22oi_1
XTAP_2580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12889_ _01677_ VGND VGND VPWR VPWR _02982_ sky130_fd_sc_hd__clkbuf_4
XTAP_2591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17416_ _07883_ _07890_ VGND VGND VPWR VPWR _07891_ sky130_fd_sc_hd__nand2_1
X_14628_ _04852_ _04854_ _04859_ VGND VGND VPWR VPWR _04860_ sky130_fd_sc_hd__or3_4
XFILLER_0_145_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18396_ _08953_ _08954_ VGND VGND VPWR VPWR _08956_ sky130_fd_sc_hd__or2_1
XTAP_1890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17347_ _06680_ _07812_ _07815_ VGND VGND VPWR VPWR _07816_ sky130_fd_sc_hd__or3_1
X_14559_ _00107_ _05888_ VGND VGND VPWR VPWR _04785_ sky130_fd_sc_hd__nand2_1
XFILLER_0_55_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17278_ _07606_ _07614_ VGND VGND VPWR VPWR _07740_ sky130_fd_sc_hd__and2_1
XFILLER_0_15_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19017_ clknet_4_9_0_clk _00002_ VGND VGND VPWR VPWR sel_op\[2\] sky130_fd_sc_hd__dfxtp_1
X_16229_ _06477_ _03029_ _02784_ _06333_ _06598_ VGND VGND VPWR VPWR _06599_ sky130_fd_sc_hd__a41o_1
XFILLER_0_70_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_468 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_141_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_6 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09603_ _04329_ _04613_ VGND VGND VPWR VPWR _05192_ sky130_fd_sc_hd__or2b_1
XFILLER_0_78_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09534_ _04427_ VGND VGND VPWR VPWR _04438_ sky130_fd_sc_hd__buf_8
XFILLER_0_39_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09465_ _03651_ _03662_ _03673_ _03618_ VGND VGND VPWR VPWR _03684_ sky130_fd_sc_hd__nand4_2
XFILLER_0_78_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_149_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_148_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_117_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_104_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10240_ _00305_ _00330_ _00331_ _00332_ VGND VGND VPWR VPWR _00333_ sky130_fd_sc_hd__and4b_2
XFILLER_0_30_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10171_ _00262_ _00263_ VGND VGND VPWR VPWR _00264_ sky130_fd_sc_hd__and2_1
XFILLER_0_100_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13930_ _04095_ _04096_ VGND VGND VPWR VPWR _04097_ sky130_fd_sc_hd__or2_1
X_13861_ _00163_ _01678_ VGND VGND VPWR VPWR _04022_ sky130_fd_sc_hd__nand2_1
X_15600_ _02998_ _04125_ _05832_ _05833_ VGND VGND VPWR VPWR _05919_ sky130_fd_sc_hd__a31o_1
X_12812_ _02903_ _02904_ VGND VGND VPWR VPWR _02905_ sky130_fd_sc_hd__xor2_1
X_16580_ _06936_ _06979_ VGND VGND VPWR VPWR _06980_ sky130_fd_sc_hd__xnor2_1
X_13792_ _03938_ _03939_ _03944_ VGND VGND VPWR VPWR _03947_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_96_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15531_ _05830_ _05843_ VGND VGND VPWR VPWR _05844_ sky130_fd_sc_hd__xor2_1
XFILLER_0_85_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12743_ _02776_ _02834_ _02835_ VGND VGND VPWR VPWR _02836_ sky130_fd_sc_hd__a21boi_1
XTAP_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18250_ _08796_ _08797_ VGND VGND VPWR VPWR _08798_ sky130_fd_sc_hd__xnor2_1
X_15462_ _05767_ _05768_ VGND VGND VPWR VPWR _05770_ sky130_fd_sc_hd__and2_1
XTAP_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12674_ _02727_ _02730_ VGND VGND VPWR VPWR _02767_ sky130_fd_sc_hd__xnor2_1
XTAP_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17201_ _07654_ _07655_ VGND VGND VPWR VPWR _07656_ sky130_fd_sc_hd__nor2_1
X_14413_ _04608_ _04609_ _04625_ VGND VGND VPWR VPWR _04626_ sky130_fd_sc_hd__and3_1
XFILLER_0_154_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11625_ _01708_ _01709_ _01610_ _01619_ VGND VGND VPWR VPWR _01718_ sky130_fd_sc_hd__a211o_1
X_18181_ _08716_ _08722_ VGND VGND VPWR VPWR _08723_ sky130_fd_sc_hd__xnor2_1
X_15393_ _05692_ _05674_ _05675_ VGND VGND VPWR VPWR _05695_ sky130_fd_sc_hd__nand3_2
XFILLER_0_5_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17132_ _03920_ _07578_ _07580_ _06484_ VGND VGND VPWR VPWR _07582_ sky130_fd_sc_hd__o211a_1
X_14344_ _04546_ _04547_ _04420_ _04397_ VGND VGND VPWR VPWR _04551_ sky130_fd_sc_hd__o211a_1
X_11556_ _06982_ _05050_ _01647_ _01648_ VGND VGND VPWR VPWR _01649_ sky130_fd_sc_hd__nand4_1
XFILLER_0_80_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_664 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10507_ _00537_ _00580_ _00581_ _00582_ VGND VGND VPWR VPWR _00600_ sky130_fd_sc_hd__nor4_1
X_17063_ _07496_ _07505_ VGND VGND VPWR VPWR _07506_ sky130_fd_sc_hd__xnor2_1
X_14275_ _00358_ _09172_ _04864_ _04143_ VGND VGND VPWR VPWR _04475_ sky130_fd_sc_hd__and4_1
X_11487_ _01576_ _01579_ VGND VGND VPWR VPWR _01580_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_21_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16014_ _06363_ _06364_ _01041_ VGND VGND VPWR VPWR _06365_ sky130_fd_sc_hd__a21bo_1
X_13226_ _03320_ _03328_ VGND VGND VPWR VPWR _03329_ sky130_fd_sc_hd__xnor2_2
X_10438_ _00349_ _00350_ _00367_ VGND VGND VPWR VPWR _00531_ sky130_fd_sc_hd__nand3_2
XFILLER_0_20_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_658 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13157_ _03252_ _03253_ _03248_ _03249_ VGND VGND VPWR VPWR _03255_ sky130_fd_sc_hd__a211o_1
XTAP_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10369_ _06460_ _00461_ _00296_ _00295_ VGND VGND VPWR VPWR _00462_ sky130_fd_sc_hd__a31o_1
XFILLER_0_21_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12108_ _02200_ _09354_ _02139_ VGND VGND VPWR VPWR _02201_ sky130_fd_sc_hd__a21o_1
XTAP_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13088_ _02257_ _03179_ _03040_ VGND VGND VPWR VPWR _03180_ sky130_fd_sc_hd__o21ai_1
X_17965_ _07207_ _07623_ _08384_ _08386_ VGND VGND VPWR VPWR _08489_ sky130_fd_sc_hd__a31o_1
X_12039_ _02123_ _02129_ _02130_ _02131_ VGND VGND VPWR VPWR _02132_ sky130_fd_sc_hd__or4_4
X_16916_ _07283_ _07284_ _07344_ VGND VGND VPWR VPWR _07346_ sky130_fd_sc_hd__and3_1
X_17896_ _08218_ _08324_ _08325_ VGND VGND VPWR VPWR _08414_ sky130_fd_sc_hd__nand3_1
X_16847_ _03920_ _07268_ _07270_ _06484_ VGND VGND VPWR VPWR _07271_ sky130_fd_sc_hd__o211a_1
Xclkbuf_4_1_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_1_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_125_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16778_ _07194_ VGND VGND VPWR VPWR _07195_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_149_129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_775 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18517_ _06416_ _06545_ _09085_ _06246_ VGND VGND VPWR VPWR _09086_ sky130_fd_sc_hd__a22o_1
X_15729_ _05989_ _05998_ _06057_ VGND VGND VPWR VPWR _06059_ sky130_fd_sc_hd__nand3_1
XFILLER_0_87_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18448_ _08915_ _08965_ _09010_ VGND VGND VPWR VPWR _09012_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_146_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18379_ _07474_ _08036_ _08937_ _06720_ VGND VGND VPWR VPWR _08938_ sky130_fd_sc_hd__o211a_1
XFILLER_0_28_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09517_ net169 ApproximateM_inst.lob_16.lob1.genblk1\[8\].genblk1.mux.sel _04242_
+ net227 VGND VGND VPWR VPWR _04253_ sky130_fd_sc_hd__a22o_1
XFILLER_0_93_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09448_ cla_inst.in2\[17\] VGND VGND VPWR VPWR _03498_ sky130_fd_sc_hd__buf_6
XPHY_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11410_ _00108_ VGND VGND VPWR VPWR _01503_ sky130_fd_sc_hd__buf_4
XFILLER_0_151_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12390_ _02435_ _02440_ VGND VGND VPWR VPWR _02483_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_151_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11341_ _01421_ _01433_ VGND VGND VPWR VPWR _01434_ sky130_fd_sc_hd__and2_1
XFILLER_0_22_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14060_ _04237_ _04239_ VGND VGND VPWR VPWR _04240_ sky130_fd_sc_hd__or2_1
XFILLER_0_104_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11272_ _01338_ _01364_ VGND VGND VPWR VPWR _01365_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_120_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_550 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13011_ _03028_ _02127_ VGND VGND VPWR VPWR _03104_ sky130_fd_sc_hd__nor2_2
X_10223_ _00314_ _00315_ VGND VGND VPWR VPWR _00316_ sky130_fd_sc_hd__xor2_1
XFILLER_0_120_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10154_ _04067_ VGND VGND VPWR VPWR _00247_ sky130_fd_sc_hd__clkbuf_8
X_17750_ _08215_ _08214_ VGND VGND VPWR VPWR _08254_ sky130_fd_sc_hd__or2b_1
X_14962_ _05208_ _05209_ _05222_ VGND VGND VPWR VPWR _05225_ sky130_fd_sc_hd__nand3_1
X_10085_ _00177_ VGND VGND VPWR VPWR _00178_ sky130_fd_sc_hd__buf_4
X_16701_ _07107_ _07110_ VGND VGND VPWR VPWR _07111_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13913_ _04077_ _04079_ _03081_ VGND VGND VPWR VPWR _04080_ sky130_fd_sc_hd__mux2_1
X_17681_ _08173_ _08178_ VGND VGND VPWR VPWR _08179_ sky130_fd_sc_hd__xnor2_1
X_14893_ _00107_ _01223_ _05145_ _05146_ VGND VGND VPWR VPWR _05150_ sky130_fd_sc_hd__a22o_1
X_13844_ _03811_ _03833_ _04002_ net239 VGND VGND VPWR VPWR _04004_ sky130_fd_sc_hd__a211oi_2
X_16632_ _06560_ _06764_ _06951_ _07035_ VGND VGND VPWR VPWR _07037_ sky130_fd_sc_hd__or4_1
XFILLER_0_69_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13775_ _03123_ _03923_ _03928_ VGND VGND VPWR VPWR _03929_ sky130_fd_sc_hd__or3_2
X_16563_ _06578_ _06961_ VGND VGND VPWR VPWR _06962_ sky130_fd_sc_hd__nor2_1
X_10987_ _07984_ _07973_ cla_inst.in1\[20\] net233 VGND VGND VPWR VPWR _01080_ sky130_fd_sc_hd__nand4_1
X_18302_ _07665_ _07516_ _08150_ _08625_ _08781_ VGND VGND VPWR VPWR _08855_ sky130_fd_sc_hd__a41o_1
XFILLER_0_139_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15514_ _05728_ _05730_ _05824_ VGND VGND VPWR VPWR _05826_ sky130_fd_sc_hd__nor3_1
X_12726_ _02804_ _02813_ _02818_ VGND VGND VPWR VPWR _02819_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_139_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_767 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16494_ _06868_ _06886_ VGND VGND VPWR VPWR _06887_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_127_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15445_ _05749_ _05750_ VGND VGND VPWR VPWR _05751_ sky130_fd_sc_hd__nand2_1
X_18233_ _08777_ _08779_ VGND VGND VPWR VPWR _08780_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_128_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12657_ _02748_ _02749_ VGND VGND VPWR VPWR _02750_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_115_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11608_ _01699_ _01691_ _01690_ VGND VGND VPWR VPWR _01701_ sky130_fd_sc_hd__and3b_1
XFILLER_0_108_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15376_ _05528_ _05531_ VGND VGND VPWR VPWR _05676_ sky130_fd_sc_hd__and2_1
XFILLER_0_108_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18164_ _07751_ _07314_ _08260_ _08625_ VGND VGND VPWR VPWR _08705_ sky130_fd_sc_hd__or4b_1
XFILLER_0_143_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12588_ _02675_ _02679_ _02680_ VGND VGND VPWR VPWR _02681_ sky130_fd_sc_hd__and3_1
XFILLER_0_52_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14327_ _04529_ _04530_ _04511_ VGND VGND VPWR VPWR _04532_ sky130_fd_sc_hd__o21a_1
XFILLER_0_40_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17115_ _02671_ _02842_ VGND VGND VPWR VPWR _07563_ sky130_fd_sc_hd__nand2_1
XFILLER_0_123_530 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11539_ _01625_ _01626_ _01629_ VGND VGND VPWR VPWR _01632_ sky130_fd_sc_hd__a21o_1
X_18095_ _08624_ _08628_ VGND VGND VPWR VPWR _08630_ sky130_fd_sc_hd__nand2_1
Xmax_cap115 _08985_ VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__buf_1
Xmax_cap126 _04670_ VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__buf_1
XFILLER_0_111_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17046_ _07486_ VGND VGND VPWR VPWR _07487_ sky130_fd_sc_hd__clkbuf_4
X_14258_ _04447_ _04455_ VGND VGND VPWR VPWR _04456_ sky130_fd_sc_hd__xnor2_2
Xmax_cap137 _02565_ VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__buf_1
XFILLER_0_150_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13209_ _03307_ _03309_ VGND VGND VPWR VPWR _03310_ sky130_fd_sc_hd__xnor2_2
XTAP_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14189_ _04378_ _04379_ _04161_ _04335_ VGND VGND VPWR VPWR _04381_ sky130_fd_sc_hd__o211a_1
XFILLER_0_29_30 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18997_ clknet_4_3_0_clk _09363_ VGND VGND VPWR VPWR salida\[50\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17948_ _08368_ _08371_ _08369_ VGND VGND VPWR VPWR _08470_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_31_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17879_ _08382_ _08287_ _08393_ VGND VGND VPWR VPWR _08395_ sky130_fd_sc_hd__nor3_1
XFILLER_0_45_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_723 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_152_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_146_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09997_ _09338_ _09337_ _06873_ _06819_ VGND VGND VPWR VPWR _09340_ sky130_fd_sc_hd__o211a_1
XFILLER_0_99_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10910_ _01001_ _01002_ VGND VGND VPWR VPWR _01003_ sky130_fd_sc_hd__and2b_1
X_11890_ _01978_ _01945_ _01976_ VGND VGND VPWR VPWR _01983_ sky130_fd_sc_hd__and3_1
XFILLER_0_98_369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10841_ _03454_ _00129_ VGND VGND VPWR VPWR _00934_ sky130_fd_sc_hd__and2_1
XFILLER_0_39_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13560_ _05921_ VGND VGND VPWR VPWR _03693_ sky130_fd_sc_hd__clkbuf_4
X_10772_ _00863_ _00864_ VGND VGND VPWR VPWR _00865_ sky130_fd_sc_hd__nor2_1
XFILLER_0_54_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12511_ _02556_ _02594_ _02603_ VGND VGND VPWR VPWR _02604_ sky130_fd_sc_hd__nand3_1
X_13491_ _03615_ _03616_ VGND VGND VPWR VPWR _03617_ sky130_fd_sc_hd__and2b_1
XFILLER_0_94_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15230_ _05426_ _05427_ _05515_ VGND VGND VPWR VPWR _05517_ sky130_fd_sc_hd__or3_2
XFILLER_0_19_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12442_ _05747_ _00132_ VGND VGND VPWR VPWR _02535_ sky130_fd_sc_hd__nand2_1
XFILLER_0_125_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_151_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_124_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_152_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15161_ _05439_ _05440_ VGND VGND VPWR VPWR _05441_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_35_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12373_ _02320_ _02312_ VGND VGND VPWR VPWR _02466_ sky130_fd_sc_hd__xnor2_1
X_14112_ _04283_ net133 _04295_ VGND VGND VPWR VPWR _04297_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_50_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_656 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11324_ _09351_ VGND VGND VPWR VPWR _01417_ sky130_fd_sc_hd__clkbuf_4
X_15092_ _05364_ _05365_ VGND VGND VPWR VPWR _05367_ sky130_fd_sc_hd__nor2_1
XFILLER_0_105_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_120_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14043_ _04218_ _04219_ _04221_ VGND VGND VPWR VPWR _04222_ sky130_fd_sc_hd__nor3_1
X_18920_ clknet_4_13_0_clk _00074_ VGND VGND VPWR VPWR ApproximateM_inst.lob_16.lob2.genblk1\[6\].genblk1.mux.sel
+ sky130_fd_sc_hd__dfxtp_2
X_11255_ _01344_ _01345_ _01346_ VGND VGND VPWR VPWR _01348_ sky130_fd_sc_hd__o21ba_1
X_10206_ _00292_ _00298_ VGND VGND VPWR VPWR _00299_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_66_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18851_ clknet_4_6_0_clk net300 VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__dfxtp_1
X_11186_ _01275_ _01276_ _01278_ VGND VGND VPWR VPWR _01279_ sky130_fd_sc_hd__a21oi_4
X_17802_ _08296_ _08310_ VGND VGND VPWR VPWR _08312_ sky130_fd_sc_hd__xnor2_1
X_10137_ _00168_ _00229_ VGND VGND VPWR VPWR _00230_ sky130_fd_sc_hd__xnor2_4
X_18782_ _09294_ VGND VGND VPWR VPWR _00085_ sky130_fd_sc_hd__buf_1
X_15994_ _06084_ _00878_ VGND VGND VPWR VPWR _06343_ sky130_fd_sc_hd__nand2_2
X_17733_ _03588_ _06383_ _06385_ VGND VGND VPWR VPWR _08237_ sky130_fd_sc_hd__nand3_1
X_14945_ _05190_ _05193_ VGND VGND VPWR VPWR _05206_ sky130_fd_sc_hd__or2b_1
X_10068_ _00141_ _00160_ VGND VGND VPWR VPWR _00161_ sky130_fd_sc_hd__or2b_1
X_17664_ _07042_ _07487_ _08056_ VGND VGND VPWR VPWR _08161_ sky130_fd_sc_hd__or3_1
X_14876_ _05128_ _05130_ VGND VGND VPWR VPWR _05131_ sky130_fd_sc_hd__or2_1
XFILLER_0_58_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16615_ _06816_ VGND VGND VPWR VPWR _07018_ sky130_fd_sc_hd__clkbuf_4
X_13827_ _03816_ _03825_ VGND VGND VPWR VPWR _03985_ sky130_fd_sc_hd__and2b_1
X_17595_ _07956_ _07961_ _08085_ VGND VGND VPWR VPWR _08086_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_85_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16546_ _05410_ _06812_ _03003_ _03004_ VGND VGND VPWR VPWR _06943_ sky130_fd_sc_hd__or4_1
X_13758_ _03093_ _03096_ _03050_ VGND VGND VPWR VPWR _03910_ sky130_fd_sc_hd__mux2_1
X_12709_ _02792_ _02793_ VGND VGND VPWR VPWR _02802_ sky130_fd_sc_hd__nor2_1
X_13689_ _03649_ _03751_ _03832_ _03833_ VGND VGND VPWR VPWR _03834_ sky130_fd_sc_hd__o211a_1
XFILLER_0_45_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16477_ _06653_ _06756_ VGND VGND VPWR VPWR _06868_ sky130_fd_sc_hd__nor2_1
XFILLER_0_38_480 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_143_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18216_ _03201_ _08760_ _08761_ VGND VGND VPWR VPWR _08762_ sky130_fd_sc_hd__and3_2
X_15428_ _05730_ _05731_ VGND VGND VPWR VPWR _05732_ sky130_fd_sc_hd__nor2_1
XFILLER_0_60_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_198 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_143_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_86 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_142_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_131_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15359_ _01505_ _00495_ VGND VGND VPWR VPWR _05657_ sky130_fd_sc_hd__nand2_1
X_18147_ _06425_ _06446_ _08686_ VGND VGND VPWR VPWR _08687_ sky130_fd_sc_hd__or3_1
XFILLER_0_40_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18078_ _08609_ _08610_ _08611_ VGND VGND VPWR VPWR _08612_ sky130_fd_sc_hd__a21oi_1
X_09920_ _08605_ _08626_ VGND VGND VPWR VPWR _08637_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_22_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17029_ _03101_ _06436_ _00593_ VGND VGND VPWR VPWR _07469_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09851_ _07690_ _07875_ VGND VGND VPWR VPWR _07886_ sky130_fd_sc_hd__xnor2_2
XTAP_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09782_ _06722_ VGND VGND VPWR VPWR _07134_ sky130_fd_sc_hd__buf_4
XTAP_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11040_ _01126_ _01132_ VGND VGND VPWR VPWR _01133_ sky130_fd_sc_hd__and2_1
XFILLER_0_102_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12991_ _03026_ _03083_ _02783_ VGND VGND VPWR VPWR _03084_ sky130_fd_sc_hd__a21bo_1
X_14730_ _02984_ _01520_ _00498_ _07015_ VGND VGND VPWR VPWR _04971_ sky130_fd_sc_hd__nand4_1
X_11942_ _02032_ _02034_ VGND VGND VPWR VPWR _02035_ sky130_fd_sc_hd__nor2_2
XFILLER_0_98_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14661_ _04885_ _04768_ _04895_ VGND VGND VPWR VPWR _04896_ sky130_fd_sc_hd__a21oi_4
X_11873_ _00846_ _05921_ _01863_ VGND VGND VPWR VPWR _01966_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_39_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16400_ _02807_ _02822_ _03201_ VGND VGND VPWR VPWR _06785_ sky130_fd_sc_hd__o21ai_1
X_13612_ _03039_ _03565_ _03584_ _03121_ _03749_ VGND VGND VPWR VPWR _09379_ sky130_fd_sc_hd__o221ai_2
X_10824_ _00914_ _00915_ _00916_ VGND VGND VPWR VPWR _00917_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_95_851 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17380_ _07822_ _07729_ _07850_ VGND VGND VPWR VPWR _07851_ sky130_fd_sc_hd__a21oi_1
X_14592_ _04818_ _04820_ VGND VGND VPWR VPWR _04822_ sky130_fd_sc_hd__nand2_1
XFILLER_0_109_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13543_ _03671_ _03672_ _03434_ _03586_ VGND VGND VPWR VPWR _03675_ sky130_fd_sc_hd__a211o_1
XFILLER_0_95_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16331_ _06707_ _06709_ _03060_ VGND VGND VPWR VPWR _06710_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10755_ _08191_ _00122_ _00847_ VGND VGND VPWR VPWR _00848_ sky130_fd_sc_hd__a21o_1
XFILLER_0_109_132 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_109_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16262_ _03077_ _06632_ _06634_ VGND VGND VPWR VPWR _06636_ sky130_fd_sc_hd__a21oi_1
X_13474_ _04088_ _03892_ _05617_ _05246_ VGND VGND VPWR VPWR _03599_ sky130_fd_sc_hd__nand4_2
X_10686_ _00762_ _00763_ _00778_ VGND VGND VPWR VPWR _00779_ sky130_fd_sc_hd__nand3_4
XFILLER_0_82_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15213_ _05460_ _05384_ _05498_ VGND VGND VPWR VPWR _05499_ sky130_fd_sc_hd__a21o_1
X_18001_ _07256_ _08515_ _08516_ _08527_ VGND VGND VPWR VPWR _08528_ sky130_fd_sc_hd__a31o_1
XFILLER_0_124_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12425_ _02516_ _02483_ _02517_ VGND VGND VPWR VPWR _02518_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_113_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_850 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16193_ _06522_ _06525_ _01113_ VGND VGND VPWR VPWR _06560_ sky130_fd_sc_hd__a21o_1
XFILLER_0_23_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_152_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15144_ _05307_ _05419_ _05423_ _03039_ VGND VGND VPWR VPWR _05424_ sky130_fd_sc_hd__o22ai_2
X_12356_ _02380_ _02381_ _02382_ _02352_ VGND VGND VPWR VPWR _02449_ sky130_fd_sc_hd__o22a_1
XFILLER_0_105_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11307_ _00843_ _00841_ _00836_ VGND VGND VPWR VPWR _01400_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_121_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15075_ _05132_ _05255_ VGND VGND VPWR VPWR _05348_ sky130_fd_sc_hd__and2b_1
XFILLER_0_77_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12287_ _02368_ _02376_ _02378_ _02379_ VGND VGND VPWR VPWR _02380_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_121_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14026_ _04201_ _04202_ VGND VGND VPWR VPWR _04203_ sky130_fd_sc_hd__xnor2_1
X_18903_ clknet_4_10_0_clk _00057_ VGND VGND VPWR VPWR cla_inst.in1\[21\] sky130_fd_sc_hd__dfxtp_1
X_11238_ net325 _01328_ _01016_ _01014_ VGND VGND VPWR VPWR _01331_ sky130_fd_sc_hd__o211a_1
X_18834_ net57 op_code\[2\] _09331_ VGND VGND VPWR VPWR _09335_ sky130_fd_sc_hd__mux2_1
X_11169_ _01243_ _01260_ VGND VGND VPWR VPWR _01262_ sky130_fd_sc_hd__nor2_1
X_18765_ _02347_ net38 _09276_ VGND VGND VPWR VPWR _09282_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15977_ _05308_ _05306_ _03920_ VGND VGND VPWR VPWR _06325_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17716_ _08216_ _08217_ VGND VGND VPWR VPWR _08218_ sky130_fd_sc_hd__xor2_1
X_14928_ _05065_ _05067_ _05187_ VGND VGND VPWR VPWR _05188_ sky130_fd_sc_hd__a21o_1
X_18696_ net48 _09189_ _09228_ VGND VGND VPWR VPWR _00057_ sky130_fd_sc_hd__o21a_1
XFILLER_0_117_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17647_ _06381_ _06790_ _08142_ _03111_ VGND VGND VPWR VPWR _08143_ sky130_fd_sc_hd__a22oi_1
X_14859_ _05110_ _05111_ VGND VGND VPWR VPWR _05112_ sky130_fd_sc_hd__nor2_1
XFILLER_0_86_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17578_ _02347_ _06891_ _07943_ VGND VGND VPWR VPWR _08067_ sky130_fd_sc_hd__and3_1
XFILLER_0_46_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16529_ _06424_ _06432_ _06924_ VGND VGND VPWR VPWR _06925_ sky130_fd_sc_hd__or3_1
XFILLER_0_133_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09903_ _04580_ VGND VGND VPWR VPWR _08452_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_111_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09834_ ApproximateM_inst.lob_16.lob2.genblk1\[1\].genblk1.mux.sel VGND VGND VPWR
+ VPWR _07700_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_67_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09765_ _05181_ _06181_ _06906_ _06928_ VGND VGND VPWR VPWR _06949_ sky130_fd_sc_hd__a211oi_1
X_09696_ _03356_ _03377_ _03903_ _03410_ VGND VGND VPWR VPWR _06202_ sky130_fd_sc_hd__nand4_2
XFILLER_0_69_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrebuffer30 _01971_ VGND VGND VPWR VPWR net193 sky130_fd_sc_hd__clkbuf_1
XTAP_2217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer41 _01659_ VGND VGND VPWR VPWR net204 sky130_fd_sc_hd__clkbuf_1
XTAP_2228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer52 net342 VGND VGND VPWR VPWR net215 sky130_fd_sc_hd__clkbuf_1
XTAP_2239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer63 net225 VGND VGND VPWR VPWR net226 sky130_fd_sc_hd__clkbuf_1
XTAP_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer74 _02043_ VGND VGND VPWR VPWR net328 sky130_fd_sc_hd__dlygate4sd1_1
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer85 _04432_ VGND VGND VPWR VPWR net332 sky130_fd_sc_hd__dlygate4sd1_1
XTAP_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer96 _06524_ VGND VGND VPWR VPWR net343 sky130_fd_sc_hd__dlygate4sd1_1
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_147_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10540_ _00620_ _00621_ _00631_ VGND VGND VPWR VPWR _00633_ sky130_fd_sc_hd__or3_4
XFILLER_0_134_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10471_ _00175_ _00563_ _00211_ _00173_ VGND VGND VPWR VPWR _00564_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_44_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12210_ _02285_ _02287_ VGND VGND VPWR VPWR _02303_ sky130_fd_sc_hd__nor2_1
X_13190_ _03268_ _03289_ VGND VGND VPWR VPWR _03290_ sky130_fd_sc_hd__xnor2_2
X_12141_ _07363_ _04067_ _02232_ _02233_ VGND VGND VPWR VPWR _02234_ sky130_fd_sc_hd__a31o_1
XFILLER_0_102_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103_875 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12072_ _01990_ _02000_ VGND VGND VPWR VPWR _02165_ sky130_fd_sc_hd__nand2_1
X_11023_ _01110_ _01111_ _01115_ VGND VGND VPWR VPWR _01116_ sky130_fd_sc_hd__or3_1
X_15900_ _06211_ _06241_ VGND VGND VPWR VPWR _06243_ sky130_fd_sc_hd__or2_1
X_16880_ _06874_ _06961_ VGND VGND VPWR VPWR _07306_ sky130_fd_sc_hd__or2_1
X_15831_ _06167_ _06168_ VGND VGND VPWR VPWR _06169_ sky130_fd_sc_hd__and2_1
X_18550_ _09119_ _09120_ _09097_ VGND VGND VPWR VPWR _09121_ sky130_fd_sc_hd__o21ai_1
X_12974_ _09059_ VGND VGND VPWR VPWR _03067_ sky130_fd_sc_hd__buf_2
X_15762_ _06088_ _06093_ VGND VGND VPWR VPWR _06095_ sky130_fd_sc_hd__or2_1
XFILLER_0_87_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17501_ _06875_ _07516_ VGND VGND VPWR VPWR _07983_ sky130_fd_sc_hd__nor2_1
XFILLER_0_151_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14713_ _04946_ _04951_ _03202_ VGND VGND VPWR VPWR _04954_ sky130_fd_sc_hd__o21a_1
X_11925_ net183 VGND VGND VPWR VPWR _02018_ sky130_fd_sc_hd__inv_2
X_18481_ _08969_ _08978_ _09011_ _09012_ _09046_ VGND VGND VPWR VPWR _09047_ sky130_fd_sc_hd__o311a_1
XTAP_2740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15693_ _02974_ _04248_ _06020_ VGND VGND VPWR VPWR _06021_ sky130_fd_sc_hd__o21a_1
XTAP_2751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17432_ _02529_ _07906_ _07907_ VGND VGND VPWR VPWR _07909_ sky130_fd_sc_hd__o21ai_2
X_14644_ _04869_ _04876_ VGND VGND VPWR VPWR _04878_ sky130_fd_sc_hd__nand2_1
X_11856_ _07363_ _00715_ _01947_ _01948_ VGND VGND VPWR VPWR _01949_ sky130_fd_sc_hd__a31o_2
XTAP_2784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10807_ _00893_ _00898_ _00430_ _00899_ VGND VGND VPWR VPWR _00900_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_95_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14575_ _04758_ _04759_ _04801_ _04802_ VGND VGND VPWR VPWR _04803_ sky130_fd_sc_hd__nand4_2
X_17363_ _07707_ _07832_ VGND VGND VPWR VPWR _07833_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_28_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11787_ _01526_ _01539_ VGND VGND VPWR VPWR _01880_ sky130_fd_sc_hd__or2_1
XFILLER_0_27_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16314_ _02810_ _03201_ _06679_ _06691_ VGND VGND VPWR VPWR _06692_ sky130_fd_sc_hd__a31o_1
X_13526_ _03654_ _00212_ _07526_ _03655_ VGND VGND VPWR VPWR _03656_ sky130_fd_sc_hd__and4b_1
X_10738_ _08017_ _00830_ VGND VGND VPWR VPWR _00831_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_103_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_422 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17294_ _07756_ _07757_ VGND VGND VPWR VPWR _07758_ sky130_fd_sc_hd__nor2_1
XFILLER_0_153_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16245_ _06611_ _06616_ _03098_ VGND VGND VPWR VPWR _06617_ sky130_fd_sc_hd__mux2_1
X_13457_ _02982_ _03135_ VGND VGND VPWR VPWR _03580_ sky130_fd_sc_hd__or2_1
X_10669_ _04296_ _04187_ _04285_ VGND VGND VPWR VPWR _00762_ sky130_fd_sc_hd__nand3_2
XFILLER_0_141_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12408_ _02485_ _02499_ VGND VGND VPWR VPWR _02501_ sky130_fd_sc_hd__xor2_1
X_13388_ _03276_ _03504_ VGND VGND VPWR VPWR _03505_ sky130_fd_sc_hd__xor2_1
X_16176_ _07657_ net168 VGND VGND VPWR VPWR _06542_ sky130_fd_sc_hd__and2_2
Xoutput106 net106 VGND VGND VPWR VPWR o_wb_data[30] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_50_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15127_ _05292_ _05294_ VGND VGND VPWR VPWR _05405_ sky130_fd_sc_hd__and2b_1
X_12339_ _02422_ _02430_ _02431_ VGND VGND VPWR VPWR _02432_ sky130_fd_sc_hd__a21oi_1
X_15058_ _05326_ _05328_ VGND VGND VPWR VPWR _05329_ sky130_fd_sc_hd__xnor2_1
X_14009_ _00877_ _05888_ _04182_ VGND VGND VPWR VPWR _04184_ sky130_fd_sc_hd__a21o_1
X_18817_ _09322_ VGND VGND VPWR VPWR _00096_ sky130_fd_sc_hd__clkbuf_1
X_09550_ _04537_ _04602_ VGND VGND VPWR VPWR _04613_ sky130_fd_sc_hd__xor2_2
X_18748_ _03790_ net64 _09251_ VGND VGND VPWR VPWR _09268_ sky130_fd_sc_hd__mux2_1
X_09481_ _03848_ VGND VGND VPWR VPWR _03859_ sky130_fd_sc_hd__clkbuf_4
X_18679_ _02045_ _09190_ _09191_ VGND VGND VPWR VPWR _09217_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_59_862 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_773 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09817_ _07504_ VGND VGND VPWR VPWR _07515_ sky130_fd_sc_hd__clkbuf_4
X_09748_ _05682_ VGND VGND VPWR VPWR _06765_ sky130_fd_sc_hd__inv_6
XTAP_2003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09679_ _06008_ VGND VGND VPWR VPWR _06019_ sky130_fd_sc_hd__clkbuf_4
XTAP_2036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11710_ _01800_ _01801_ _01771_ _01781_ VGND VGND VPWR VPWR _01803_ sky130_fd_sc_hd__a211o_1
XTAP_2058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_607 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12690_ _00120_ _09219_ VGND VGND VPWR VPWR _02783_ sky130_fd_sc_hd__nand2_2
XTAP_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11641_ _01732_ _01731_ _01636_ _01633_ VGND VGND VPWR VPWR _01734_ sky130_fd_sc_hd__o211a_1
XTAP_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14360_ _02984_ _01520_ _07962_ _05964_ VGND VGND VPWR VPWR _04567_ sky130_fd_sc_hd__and4_1
XFILLER_0_64_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11572_ _01645_ _01664_ VGND VGND VPWR VPWR _01665_ sky130_fd_sc_hd__nand2_2
XFILLER_0_91_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13311_ _05834_ _08224_ _03417_ _03418_ VGND VGND VPWR VPWR _03420_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_135_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput19 i_wb_addr[25] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10523_ _00614_ _00615_ VGND VGND VPWR VPWR _00616_ sky130_fd_sc_hd__xor2_1
XFILLER_0_64_386 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14291_ _04317_ _04327_ VGND VGND VPWR VPWR _04492_ sky130_fd_sc_hd__nand2_1
XFILLER_0_150_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_135_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13242_ _00741_ _00743_ VGND VGND VPWR VPWR _03346_ sky130_fd_sc_hd__nor2_1
X_16030_ _02988_ _03111_ VGND VGND VPWR VPWR _06382_ sky130_fd_sc_hd__nand2_1
XFILLER_0_122_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10454_ _00109_ _09349_ _00171_ _00177_ VGND VGND VPWR VPWR _00547_ sky130_fd_sc_hd__and4_1
X_13173_ _03270_ _00172_ _07537_ _03271_ VGND VGND VPWR VPWR _03272_ sky130_fd_sc_hd__and4b_1
X_10385_ _05649_ _07406_ _07112_ _06029_ VGND VGND VPWR VPWR _00478_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12124_ _06765_ _02214_ _02211_ _02216_ VGND VGND VPWR VPWR _02217_ sky130_fd_sc_hd__o22a_1
X_17981_ _08447_ _08419_ _08505_ VGND VGND VPWR VPWR _08506_ sky130_fd_sc_hd__o21a_1
X_12055_ _02143_ _02146_ _02065_ _02147_ VGND VGND VPWR VPWR _02148_ sky130_fd_sc_hd__o211a_1
X_16932_ _06361_ _06360_ _06359_ VGND VGND VPWR VPWR _07364_ sky130_fd_sc_hd__a21oi_1
X_11006_ _00832_ _05617_ _01080_ _01083_ VGND VGND VPWR VPWR _01099_ sky130_fd_sc_hd__a22o_1
XFILLER_0_74_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16863_ net331 _07194_ VGND VGND VPWR VPWR _07288_ sky130_fd_sc_hd__nor2_1
X_18602_ _09113_ VGND VGND VPWR VPWR _09159_ sky130_fd_sc_hd__buf_2
X_15814_ _03537_ _04557_ VGND VGND VPWR VPWR _06151_ sky130_fd_sc_hd__nor2_1
XFILLER_0_99_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16794_ _07114_ VGND VGND VPWR VPWR _07213_ sky130_fd_sc_hd__inv_2
X_18533_ net32 net4 net3 net6 VGND VGND VPWR VPWR _09103_ sky130_fd_sc_hd__or4_1
X_15745_ _05947_ _05950_ _06015_ VGND VGND VPWR VPWR _06077_ sky130_fd_sc_hd__or3_1
X_12957_ _03049_ VGND VGND VPWR VPWR _03050_ sky130_fd_sc_hd__clkbuf_4
X_11908_ _04493_ _04416_ ApproximateM_inst.lob_16.lob1.genblk1\[2\].genblk1.mux.sel
+ ApproximateM_inst.lob_16.lob1.genblk1\[1\].genblk1.mux.sel VGND VGND VPWR VPWR _02001_
+ sky130_fd_sc_hd__and4_1
X_18464_ _03013_ _06593_ _06594_ VGND VGND VPWR VPWR _09030_ sky130_fd_sc_hd__a21o_1
XFILLER_0_47_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15676_ _05968_ _06000_ _06001_ VGND VGND VPWR VPWR _06002_ sky130_fd_sc_hd__nand3_1
XFILLER_0_87_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12888_ _02980_ VGND VGND VPWR VPWR _02981_ sky130_fd_sc_hd__buf_4
XTAP_2581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17415_ _07888_ _07889_ VGND VGND VPWR VPWR _07890_ sky130_fd_sc_hd__xnor2_1
X_14627_ _04858_ VGND VGND VPWR VPWR _04859_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11839_ _01928_ _01931_ VGND VGND VPWR VPWR _01932_ sky130_fd_sc_hd__and2_1
X_18395_ _08953_ _08954_ VGND VGND VPWR VPWR _08955_ sky130_fd_sc_hd__nand2_1
XTAP_1880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17346_ _02972_ _07813_ _07814_ _06484_ VGND VGND VPWR VPWR _07815_ sky130_fd_sc_hd__o211a_1
XFILLER_0_128_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14558_ _04782_ _04783_ VGND VGND VPWR VPWR _04784_ sky130_fd_sc_hd__nor2_1
XFILLER_0_83_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13509_ _03631_ _03419_ _03635_ _03636_ VGND VGND VPWR VPWR _03637_ sky130_fd_sc_hd__o211ai_2
X_17277_ _07488_ _07612_ VGND VGND VPWR VPWR _07739_ sky130_fd_sc_hd__and2b_1
X_14489_ _03651_ _03596_ _07004_ _06722_ VGND VGND VPWR VPWR _04708_ sky130_fd_sc_hd__nand4_2
XFILLER_0_3_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19016_ clknet_4_9_0_clk _00001_ VGND VGND VPWR VPWR sel_op\[1\] sky130_fd_sc_hd__dfxtp_1
X_16228_ _06597_ VGND VGND VPWR VPWR _06598_ sky130_fd_sc_hd__buf_4
XFILLER_0_12_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16159_ ApproximateM_inst.lob_16.lob2.genblk1\[10\].genblk1.mux.sel ApproximateM_inst.lob_16.lob2.genblk1\[9\].genblk1.mux.sel
+ sel_op\[0\] VGND VGND VPWR VPWR _06523_ sky130_fd_sc_hd__or3b_1
XFILLER_0_48_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09602_ _04318_ _04766_ _05159_ _05170_ VGND VGND VPWR VPWR _05181_ sky130_fd_sc_hd__a211o_2
XFILLER_0_79_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09533_ _04416_ VGND VGND VPWR VPWR _04427_ sky130_fd_sc_hd__buf_6
XFILLER_0_64_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09464_ _03476_ VGND VGND VPWR VPWR _03673_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_38_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_148_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_386 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_105_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10170_ _00261_ _00250_ _00251_ VGND VGND VPWR VPWR _00263_ sky130_fd_sc_hd__or3_1
XFILLER_0_100_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13860_ _04018_ _04020_ VGND VGND VPWR VPWR _04021_ sky130_fd_sc_hd__xnor2_2
X_12811_ _01470_ _01472_ _01483_ VGND VGND VPWR VPWR _02904_ sky130_fd_sc_hd__a21o_1
X_13791_ _03938_ _03939_ _03944_ VGND VGND VPWR VPWR _03945_ sky130_fd_sc_hd__and3_2
XFILLER_0_97_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15530_ _05841_ _05842_ VGND VGND VPWR VPWR _05843_ sky130_fd_sc_hd__nor2_1
XTAP_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12742_ _02777_ _02833_ VGND VGND VPWR VPWR _02835_ sky130_fd_sc_hd__nand2_1
XTAP_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_139_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15461_ _05760_ _05766_ VGND VGND VPWR VPWR _05768_ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_832 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12673_ _02764_ _02765_ VGND VGND VPWR VPWR _02766_ sky130_fd_sc_hd__or2b_1
XTAP_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17200_ _07652_ _07531_ _07653_ VGND VGND VPWR VPWR _07655_ sky130_fd_sc_hd__and3_1
XFILLER_0_37_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14412_ _04622_ _04623_ VGND VGND VPWR VPWR _04625_ sky130_fd_sc_hd__and2_1
XTAP_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11624_ _01713_ _01714_ _01715_ VGND VGND VPWR VPWR _01717_ sky130_fd_sc_hd__a21o_1
X_18180_ _08720_ _08721_ VGND VGND VPWR VPWR _08722_ sky130_fd_sc_hd__nor2_1
X_15392_ _05674_ _05675_ _05692_ VGND VGND VPWR VPWR _05694_ sky130_fd_sc_hd__a21o_1
XFILLER_0_65_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17131_ _02973_ _07579_ VGND VGND VPWR VPWR _07580_ sky130_fd_sc_hd__nand2_1
X_11555_ _07254_ _00439_ _04384_ _07232_ VGND VGND VPWR VPWR _01648_ sky130_fd_sc_hd__a22o_1
X_14343_ net342 VGND VGND VPWR VPWR _04550_ sky130_fd_sc_hd__inv_2
XFILLER_0_108_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_107_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10506_ _00418_ _00421_ _00585_ _00586_ VGND VGND VPWR VPWR _00599_ sky130_fd_sc_hd__a211oi_2
X_14274_ _03005_ _00247_ VGND VGND VPWR VPWR _04474_ sky130_fd_sc_hd__nand2_1
XFILLER_0_80_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17062_ _07502_ _07503_ VGND VGND VPWR VPWR _07505_ sky130_fd_sc_hd__or2_1
XFILLER_0_150_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11486_ _01577_ _01578_ VGND VGND VPWR VPWR _01579_ sky130_fd_sc_hd__and2b_1
XFILLER_0_100_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13225_ _03326_ _03327_ VGND VGND VPWR VPWR _03328_ sky130_fd_sc_hd__xnor2_2
X_16013_ _08615_ _00399_ VGND VGND VPWR VPWR _06364_ sky130_fd_sc_hd__or2_1
X_10437_ _00528_ _00527_ _00331_ _00326_ VGND VGND VPWR VPWR _00530_ sky130_fd_sc_hd__o211a_2
XFILLER_0_0_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_122_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13156_ _03248_ _03249_ _03252_ _03253_ VGND VGND VPWR VPWR _03254_ sky130_fd_sc_hd__o211ai_4
XTAP_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10368_ _00460_ VGND VGND VPWR VPWR _00461_ sky130_fd_sc_hd__clkbuf_8
XTAP_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12107_ _02059_ VGND VGND VPWR VPWR _02200_ sky130_fd_sc_hd__clkbuf_8
XTAP_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13087_ _03028_ _02045_ VGND VGND VPWR VPWR _03179_ sky130_fd_sc_hd__nor2_1
X_17964_ _07302_ _07303_ _07741_ _07861_ VGND VGND VPWR VPWR _08488_ sky130_fd_sc_hd__or4_2
X_10299_ _00386_ _00391_ VGND VGND VPWR VPWR _00392_ sky130_fd_sc_hd__xnor2_1
X_12038_ _02126_ _02128_ VGND VGND VPWR VPWR _02131_ sky130_fd_sc_hd__nor2_1
X_16915_ _07283_ _07284_ _07344_ VGND VGND VPWR VPWR _07345_ sky130_fd_sc_hd__a21oi_2
X_17895_ _08320_ _08412_ VGND VGND VPWR VPWR _08413_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_18_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16846_ _02973_ _07269_ VGND VGND VPWR VPWR _07270_ sky130_fd_sc_hd__nand2_1
X_16777_ _00645_ _07105_ VGND VGND VPWR VPWR _07194_ sky130_fd_sc_hd__nand2_4
X_13989_ _04149_ _04150_ _04160_ VGND VGND VPWR VPWR _04162_ sky130_fd_sc_hd__or3_1
XFILLER_0_87_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18516_ _06200_ _06592_ _06551_ VGND VGND VPWR VPWR _09085_ sky130_fd_sc_hd__a21o_1
XFILLER_0_125_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15728_ _05989_ _05998_ _06057_ VGND VGND VPWR VPWR _06058_ sky130_fd_sc_hd__a21o_1
XFILLER_0_88_787 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18447_ _08915_ _08965_ _09010_ VGND VGND VPWR VPWR _09011_ sky130_fd_sc_hd__nor3_1
X_15659_ _05972_ _05982_ VGND VGND VPWR VPWR _05983_ sky130_fd_sc_hd__xor2_1
XFILLER_0_145_303 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_146_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18378_ _06405_ _06790_ _08936_ _03068_ VGND VGND VPWR VPWR _08937_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_44_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_141_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17329_ _03206_ _07795_ VGND VGND VPWR VPWR _07796_ sky130_fd_sc_hd__nor2_1
XFILLER_0_114_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_754 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09516_ ApproximateM_inst.lob_16.lob1.genblk1\[6\].genblk1.mux.sel VGND VGND VPWR
+ VPWR _04242_ sky130_fd_sc_hd__buf_6
XFILLER_0_78_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09447_ _03465_ _03476_ VGND VGND VPWR VPWR _03487_ sky130_fd_sc_hd__and2_1
XPHY_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_117_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_117_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11340_ _01422_ _01432_ VGND VGND VPWR VPWR _01433_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_6_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11271_ _01362_ _01363_ VGND VGND VPWR VPWR _01364_ sky130_fd_sc_hd__nor2_1
XFILLER_0_61_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13010_ _03040_ _03102_ VGND VGND VPWR VPWR _03103_ sky130_fd_sc_hd__nand2_1
X_10222_ _05834_ _05986_ _08778_ _08768_ VGND VGND VPWR VPWR _00315_ sky130_fd_sc_hd__a31o_1
XFILLER_0_30_562 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10153_ _00244_ _00157_ _00232_ VGND VGND VPWR VPWR _00246_ sky130_fd_sc_hd__or3_1
X_14961_ _05208_ _05209_ _05222_ VGND VGND VPWR VPWR _05223_ sky130_fd_sc_hd__a21o_1
X_10084_ _00176_ VGND VGND VPWR VPWR _00177_ sky130_fd_sc_hd__buf_6
X_16700_ _06937_ _06961_ _07109_ _06542_ VGND VGND VPWR VPWR _07110_ sky130_fd_sc_hd__a2bb2o_1
X_13912_ _03062_ _03163_ VGND VGND VPWR VPWR _04079_ sky130_fd_sc_hd__nor2_1
X_17680_ _08176_ _08177_ VGND VGND VPWR VPWR _08178_ sky130_fd_sc_hd__xor2_1
X_14892_ _05147_ VGND VGND VPWR VPWR _05149_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16631_ _07033_ _07034_ _00207_ VGND VGND VPWR VPWR _07035_ sky130_fd_sc_hd__o21ai_4
X_13843_ _03983_ _03984_ _04000_ VGND VGND VPWR VPWR _04003_ sky130_fd_sc_hd__o21a_1
XFILLER_0_69_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_18 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16562_ _06880_ VGND VGND VPWR VPWR _06961_ sky130_fd_sc_hd__buf_2
X_10986_ _01020_ _01021_ _01078_ VGND VGND VPWR VPWR _01079_ sky130_fd_sc_hd__or3_4
X_13774_ _03117_ _03927_ _03036_ VGND VGND VPWR VPWR _03928_ sky130_fd_sc_hd__o21a_1
X_18301_ _08847_ _08852_ VGND VGND VPWR VPWR _08853_ sky130_fd_sc_hd__xnor2_1
X_15513_ _05728_ _05730_ _05824_ VGND VGND VPWR VPWR _05825_ sky130_fd_sc_hd__o21a_1
X_12725_ _02814_ _02817_ VGND VGND VPWR VPWR _02818_ sky130_fd_sc_hd__nor2_1
X_16493_ _06876_ _06885_ VGND VGND VPWR VPWR _06886_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_128_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_139_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18232_ _07314_ _08260_ _08625_ VGND VGND VPWR VPWR _08779_ sky130_fd_sc_hd__or3_1
X_15444_ _03000_ _05652_ _05748_ VGND VGND VPWR VPWR _05750_ sky130_fd_sc_hd__a21o_1
XFILLER_0_37_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12656_ _02694_ _02708_ _02707_ VGND VGND VPWR VPWR _02749_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_37_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11607_ _01690_ _01691_ _01699_ VGND VGND VPWR VPWR _01700_ sky130_fd_sc_hd__a21boi_1
X_18163_ _08701_ _08703_ VGND VGND VPWR VPWR _08704_ sky130_fd_sc_hd__xnor2_1
X_15375_ _05672_ _05673_ _05571_ _05629_ VGND VGND VPWR VPWR _05675_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_5_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12587_ _02638_ _02637_ _02636_ VGND VGND VPWR VPWR _02680_ sky130_fd_sc_hd__a21o_1
XFILLER_0_136_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_142_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17114_ _02671_ _02842_ VGND VGND VPWR VPWR _07562_ sky130_fd_sc_hd__or2_1
X_14326_ _04511_ _04529_ _04530_ VGND VGND VPWR VPWR _04531_ sky130_fd_sc_hd__nor3_2
XFILLER_0_52_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_676 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_135_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11538_ _01547_ _01549_ _01546_ VGND VGND VPWR VPWR _01631_ sky130_fd_sc_hd__a21o_1
X_18094_ _08624_ _08628_ VGND VGND VPWR VPWR _08629_ sky130_fd_sc_hd__or2_1
XFILLER_0_123_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_cap127 _04428_ VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__buf_1
X_17045_ _02188_ _06889_ VGND VGND VPWR VPWR _07486_ sky130_fd_sc_hd__nand2_1
X_14257_ _04448_ _04454_ VGND VGND VPWR VPWR _04455_ sky130_fd_sc_hd__xnor2_2
X_11469_ _01550_ _01561_ VGND VGND VPWR VPWR _01562_ sky130_fd_sc_hd__nor2_1
Xmax_cap138 _01843_ VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_151_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_394 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13208_ _00709_ _00710_ _03308_ VGND VGND VPWR VPWR _03309_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_0_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14188_ _04161_ _04335_ _04378_ _04379_ VGND VGND VPWR VPWR _04380_ sky130_fd_sc_hd__a211oi_2
XTAP_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13139_ _03226_ _03235_ VGND VGND VPWR VPWR _03236_ sky130_fd_sc_hd__xnor2_1
XTAP_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18996_ clknet_4_6_0_clk _09362_ VGND VGND VPWR VPWR salida\[49\] sky130_fd_sc_hd__dfxtp_1
XTAP_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17947_ _08467_ _08468_ VGND VGND VPWR VPWR _08469_ sky130_fd_sc_hd__nor2_1
X_17878_ _08382_ _08287_ _08393_ VGND VGND VPWR VPWR _08394_ sky130_fd_sc_hd__o21a_1
XFILLER_0_24_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16829_ _07157_ _07154_ VGND VGND VPWR VPWR _07251_ sky130_fd_sc_hd__and2b_1
XFILLER_0_45_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_146_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_118_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09996_ _06819_ _06873_ _09337_ _09338_ VGND VGND VPWR VPWR _09339_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_86_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10840_ _00916_ _00915_ _00914_ VGND VGND VPWR VPWR _00933_ sky130_fd_sc_hd__a21o_1
XFILLER_0_39_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10771_ _00105_ _00117_ VGND VGND VPWR VPWR _00864_ sky130_fd_sc_hd__xnor2_1
X_12510_ _02598_ _02601_ _02602_ VGND VGND VPWR VPWR _02603_ sky130_fd_sc_hd__a21bo_1
X_13490_ _03613_ _03614_ _03610_ VGND VGND VPWR VPWR _03616_ sky130_fd_sc_hd__a21o_1
X_12441_ _02533_ _09354_ VGND VGND VPWR VPWR _02534_ sky130_fd_sc_hd__nand2_1
XFILLER_0_124_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_151_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15160_ _05320_ _05324_ VGND VGND VPWR VPWR _05440_ sky130_fd_sc_hd__or2_1
X_12372_ _02462_ _02464_ VGND VGND VPWR VPWR _02465_ sky130_fd_sc_hd__nand2_1
XFILLER_0_50_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14111_ _04286_ _04294_ VGND VGND VPWR VPWR _04295_ sky130_fd_sc_hd__xnor2_2
X_11323_ _01330_ _01332_ VGND VGND VPWR VPWR _01416_ sky130_fd_sc_hd__or2b_1
X_15091_ _05348_ _05349_ _05363_ VGND VGND VPWR VPWR _05365_ sky130_fd_sc_hd__nor3_1
Xclkbuf_4_0_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_0_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_22_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14042_ _04004_ _04050_ VGND VGND VPWR VPWR _04221_ sky130_fd_sc_hd__and2b_1
X_11254_ _01344_ _01345_ _01346_ VGND VGND VPWR VPWR _01347_ sky130_fd_sc_hd__nor3b_2
X_10205_ _00293_ _00297_ VGND VGND VPWR VPWR _00298_ sky130_fd_sc_hd__xnor2_1
X_18850_ clknet_4_6_0_clk net298 VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__dfxtp_1
X_11185_ _00768_ _01277_ VGND VGND VPWR VPWR _01278_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_66_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17801_ _08298_ _08309_ VGND VGND VPWR VPWR _08310_ sky130_fd_sc_hd__xnor2_1
X_10136_ _00227_ _00228_ VGND VGND VPWR VPWR _00229_ sky130_fd_sc_hd__and2b_1
X_18781_ _09273_ _09293_ VGND VGND VPWR VPWR _09294_ sky130_fd_sc_hd__and2_1
X_15993_ _06339_ _06341_ VGND VGND VPWR VPWR _06342_ sky130_fd_sc_hd__or2b_1
X_17732_ _08230_ _08231_ _08233_ VGND VGND VPWR VPWR _08236_ sky130_fd_sc_hd__nand3_1
X_10067_ _00142_ _00159_ VGND VGND VPWR VPWR _00160_ sky130_fd_sc_hd__xor2_2
X_14944_ _03125_ _05096_ _05099_ _03199_ _05205_ VGND VGND VPWR VPWR _09359_ sky130_fd_sc_hd__a221o_1
XFILLER_0_89_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17663_ _07143_ _07487_ _08056_ VGND VGND VPWR VPWR _08160_ sky130_fd_sc_hd__o21ai_1
X_14875_ _07635_ _05888_ _05129_ _05125_ VGND VGND VPWR VPWR _05130_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_15_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16614_ _06940_ _06965_ VGND VGND VPWR VPWR _07017_ sky130_fd_sc_hd__nand2_1
X_13826_ _03786_ _03810_ _03981_ _03982_ VGND VGND VPWR VPWR _03984_ sky130_fd_sc_hd__o211a_1
X_17594_ _07963_ _07955_ VGND VGND VPWR VPWR _08085_ sky130_fd_sc_hd__or2b_1
XFILLER_0_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16545_ _03313_ net150 _06805_ VGND VGND VPWR VPWR _06942_ sky130_fd_sc_hd__or3_1
XFILLER_0_128_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13757_ _03103_ _03105_ _03090_ VGND VGND VPWR VPWR _03909_ sky130_fd_sc_hd__mux2_1
X_10969_ _01060_ _01057_ VGND VGND VPWR VPWR _01062_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_57_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12708_ _02776_ _02778_ _02798_ _02800_ VGND VGND VPWR VPWR _02801_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_72_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16476_ _06572_ _06756_ _06820_ VGND VGND VPWR VPWR _06867_ sky130_fd_sc_hd__or3_2
X_13688_ _03811_ _03812_ _03831_ VGND VGND VPWR VPWR _03833_ sky130_fd_sc_hd__nand3_2
XFILLER_0_122_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18215_ _02871_ _02172_ _02470_ _02851_ VGND VGND VPWR VPWR _08761_ sky130_fd_sc_hd__or4_1
XFILLER_0_128_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15427_ _05728_ _05729_ _05634_ _05636_ VGND VGND VPWR VPWR _05731_ sky130_fd_sc_hd__o211a_1
XFILLER_0_38_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12639_ _02693_ _02696_ _02699_ VGND VGND VPWR VPWR _02732_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_14_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18146_ _04647_ _06445_ _03052_ VGND VGND VPWR VPWR _08686_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_142_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15358_ _05654_ _05655_ VGND VGND VPWR VPWR _05656_ sky130_fd_sc_hd__nor2_1
XFILLER_0_81_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14309_ _04360_ _04366_ VGND VGND VPWR VPWR _04512_ sky130_fd_sc_hd__and2b_1
XFILLER_0_151_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18077_ _08609_ _08610_ _06508_ VGND VGND VPWR VPWR _08611_ sky130_fd_sc_hd__o21ai_1
X_15289_ _05579_ _05580_ VGND VGND VPWR VPWR _05581_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_1_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17028_ _06598_ _07466_ _07467_ VGND VGND VPWR VPWR _07468_ sky130_fd_sc_hd__or3_1
XFILLER_0_0_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09850_ _07831_ _07842_ _07864_ VGND VGND VPWR VPWR _07875_ sky130_fd_sc_hd__and3b_1
XTAP_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09781_ _07112_ VGND VGND VPWR VPWR _07123_ sky130_fd_sc_hd__clkbuf_8
XTAP_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18979_ clknet_4_0_0_clk _09418_ VGND VGND VPWR VPWR salida\[32\] sky130_fd_sc_hd__dfxtp_1
XTAP_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_134_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09979_ _09197_ _09205_ _07526_ _09219_ VGND VGND VPWR VPWR _09226_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_99_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12990_ _01248_ VGND VGND VPWR VPWR _03083_ sky130_fd_sc_hd__clkbuf_4
X_11941_ _02032_ _02033_ ApproximateM_inst.lob_16.lob2.genblk1\[5\].genblk1.mux.sel
+ _03476_ VGND VGND VPWR VPWR _02034_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_98_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14660_ _04893_ _04894_ VGND VGND VPWR VPWR _04895_ sky130_fd_sc_hd__xor2_2
XFILLER_0_98_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11872_ _01864_ _01964_ VGND VGND VPWR VPWR _01965_ sky130_fd_sc_hd__nor2_1
X_13611_ _03747_ _03748_ VGND VGND VPWR VPWR _03749_ sky130_fd_sc_hd__nand2_1
X_10823_ net229 net169 _00772_ _00129_ VGND VGND VPWR VPWR _00916_ sky130_fd_sc_hd__nand4_2
X_14591_ _04819_ _04695_ VGND VGND VPWR VPWR _04820_ sky130_fd_sc_hd__nor2_1
XFILLER_0_95_863 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16330_ _03089_ _02257_ _03181_ _06626_ _06708_ VGND VGND VPWR VPWR _06709_ sky130_fd_sc_hd__o311a_1
X_13542_ _03434_ _03586_ _03671_ _03672_ VGND VGND VPWR VPWR _03674_ sky130_fd_sc_hd__o211ai_2
X_10754_ _00846_ _00322_ _08180_ VGND VGND VPWR VPWR _00847_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_94_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_144 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16261_ _03062_ _06470_ _06633_ _03913_ VGND VGND VPWR VPWR _06634_ sky130_fd_sc_hd__a31o_1
X_13473_ _03782_ _08746_ _06613_ _03881_ VGND VGND VPWR VPWR _03598_ sky130_fd_sc_hd__a22o_1
X_10685_ _00768_ _00776_ _00777_ VGND VGND VPWR VPWR _00778_ sky130_fd_sc_hd__a21o_1
X_18000_ _08520_ _08522_ _08525_ _08526_ VGND VGND VPWR VPWR _08527_ sky130_fd_sc_hd__nand4_1
X_15212_ _05480_ _05496_ VGND VGND VPWR VPWR _05498_ sky130_fd_sc_hd__xnor2_1
X_12424_ _02484_ _02509_ VGND VGND VPWR VPWR _02517_ sky130_fd_sc_hd__or2b_1
X_16192_ _03195_ VGND VGND VPWR VPWR _06559_ sky130_fd_sc_hd__buf_4
XFILLER_0_23_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_124_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15143_ _05420_ _05422_ _03536_ VGND VGND VPWR VPWR _05423_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12355_ _02417_ _02446_ _02447_ VGND VGND VPWR VPWR _02448_ sky130_fd_sc_hd__nand3_2
XFILLER_0_133_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11306_ _00843_ _00836_ _00841_ VGND VGND VPWR VPWR _01399_ sky130_fd_sc_hd__and3_1
X_15074_ _05345_ _05346_ VGND VGND VPWR VPWR _05347_ sky130_fd_sc_hd__xnor2_1
X_12286_ _02264_ _02377_ _02344_ VGND VGND VPWR VPWR _02379_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_121_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14025_ _00106_ _01575_ VGND VGND VPWR VPWR _04202_ sky130_fd_sc_hd__nand2_1
X_11237_ _01014_ _01016_ _01328_ net141 VGND VGND VPWR VPWR _01330_ sky130_fd_sc_hd__a211oi_4
X_18902_ clknet_4_10_0_clk _00056_ VGND VGND VPWR VPWR cla_inst.in1\[20\] sky130_fd_sc_hd__dfxtp_2
X_11168_ _01243_ _01260_ VGND VGND VPWR VPWR _01261_ sky130_fd_sc_hd__and2_1
X_18833_ _09334_ VGND VGND VPWR VPWR _00102_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_93_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10119_ _00211_ VGND VGND VPWR VPWR _00212_ sky130_fd_sc_hd__clkbuf_4
X_18764_ _09281_ VGND VGND VPWR VPWR _00079_ sky130_fd_sc_hd__buf_1
X_11099_ _01187_ _01188_ _01191_ VGND VGND VPWR VPWR _01192_ sky130_fd_sc_hd__nand3_4
X_15976_ _06314_ _06320_ _06322_ _02969_ VGND VGND VPWR VPWR _06324_ sky130_fd_sc_hd__a31o_1
X_17715_ _08111_ _08112_ _08116_ VGND VGND VPWR VPWR _08217_ sky130_fd_sc_hd__a21o_1
X_14927_ _05059_ _05186_ VGND VGND VPWR VPWR _05187_ sky130_fd_sc_hd__xnor2_1
X_18695_ _00813_ _09183_ _09191_ VGND VGND VPWR VPWR _09228_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_78_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17646_ _02988_ _06593_ _06594_ VGND VGND VPWR VPWR _08142_ sky130_fd_sc_hd__a21o_1
X_14858_ _02989_ _04034_ _03455_ _00513_ VGND VGND VPWR VPWR _05111_ sky130_fd_sc_hd__and4_2
X_13809_ _03800_ _03802_ VGND VGND VPWR VPWR _03965_ sky130_fd_sc_hd__and2_1
X_17577_ _07106_ _07332_ _07957_ _07958_ VGND VGND VPWR VPWR _08066_ sky130_fd_sc_hd__o31a_1
X_14789_ _04892_ _04891_ VGND VGND VPWR VPWR _05036_ sky130_fd_sc_hd__or2b_1
X_16528_ _03086_ _06851_ VGND VGND VPWR VPWR _06924_ sky130_fd_sc_hd__nor2_1
XFILLER_0_58_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_128_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16459_ _03920_ _06848_ VGND VGND VPWR VPWR _06849_ sky130_fd_sc_hd__nor2_1
XFILLER_0_128_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_367 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18129_ _08665_ _08666_ VGND VGND VPWR VPWR _08667_ sky130_fd_sc_hd__xnor2_1
X_09902_ _08420_ _08431_ VGND VGND VPWR VPWR _08442_ sky130_fd_sc_hd__nor2_1
XTAP_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09833_ _07624_ _07679_ VGND VGND VPWR VPWR _07690_ sky130_fd_sc_hd__nor2_1
XTAP_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09764_ _05181_ _06181_ _06906_ _06928_ VGND VGND VPWR VPWR _06938_ sky130_fd_sc_hd__a211o_2
X_09695_ _04973_ _05137_ _05148_ VGND VGND VPWR VPWR _06191_ sky130_fd_sc_hd__nand3_1
Xrebuffer20 _01950_ VGND VGND VPWR VPWR net183 sky130_fd_sc_hd__clkbuf_1
XTAP_2207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer31 _00941_ VGND VGND VPWR VPWR net194 sky130_fd_sc_hd__clkbuf_1
XTAP_2218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer42 _07062_ VGND VGND VPWR VPWR net205 sky130_fd_sc_hd__buf_1
XTAP_2229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer53 _06232_ VGND VGND VPWR VPWR net216 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_96_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer64 _03520_ VGND VGND VPWR VPWR net227 sky130_fd_sc_hd__buf_6
XTAP_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_690 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xrebuffer75 _07615_ VGND VGND VPWR VPWR net238 sky130_fd_sc_hd__clkbuf_1
Xrebuffer86 _04432_ VGND VGND VPWR VPWR net333 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_139_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer97 net343 VGND VGND VPWR VPWR net344 sky130_fd_sc_hd__dlygate4sd1_1
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_146_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10470_ _03476_ VGND VGND VPWR VPWR _00563_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_150_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12140_ _07221_ _07243_ _00949_ _03421_ VGND VGND VPWR VPWR _02233_ sky130_fd_sc_hd__and4_1
XFILLER_0_103_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12071_ _02161_ _02163_ VGND VGND VPWR VPWR _02164_ sky130_fd_sc_hd__and2b_1
X_11022_ _00845_ _01112_ _01114_ VGND VGND VPWR VPWR _01115_ sky130_fd_sc_hd__a21oi_4
X_15830_ _06104_ _06108_ _06166_ VGND VGND VPWR VPWR _06168_ sky130_fd_sc_hd__nand3_1
X_15761_ _06091_ _06092_ VGND VGND VPWR VPWR _06093_ sky130_fd_sc_hd__xor2_1
X_12973_ _03050_ _03065_ VGND VGND VPWR VPWR _03066_ sky130_fd_sc_hd__or2_1
X_17500_ _07980_ _07981_ VGND VGND VPWR VPWR _07982_ sky130_fd_sc_hd__nand2_1
X_14712_ _04946_ _04951_ VGND VGND VPWR VPWR _04953_ sky130_fd_sc_hd__nand2_1
X_11924_ _02011_ _02015_ VGND VGND VPWR VPWR _02017_ sky130_fd_sc_hd__xor2_1
X_18480_ _09044_ _09045_ VGND VGND VPWR VPWR _09046_ sky130_fd_sc_hd__nor2_1
XTAP_2730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15692_ _03536_ _03912_ _04243_ VGND VGND VPWR VPWR _06020_ sky130_fd_sc_hd__or3_1
XTAP_2741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17431_ _02529_ _07906_ _04238_ VGND VGND VPWR VPWR _07907_ sky130_fd_sc_hd__a21oi_1
XTAP_2763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14643_ _04869_ _04876_ VGND VGND VPWR VPWR _04877_ sky130_fd_sc_hd__or2_1
XTAP_2774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11855_ ApproximateM_inst.lob_16.lob2.genblk1\[4\].genblk1.mux.sel ApproximateM_inst.lob_16.lob2.genblk1\[3\].genblk1.mux.sel
+ ApproximateM_inst.lob_16.lob1.genblk1\[12\].genblk1.mux.sel _03826_ VGND VGND VPWR
+ VPWR _01948_ sky130_fd_sc_hd__and4_1
XTAP_2785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_362 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10806_ _00427_ _00429_ _00428_ _00270_ VGND VGND VPWR VPWR _00899_ sky130_fd_sc_hd__o211a_1
XFILLER_0_55_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17362_ _07829_ _07830_ VGND VGND VPWR VPWR _07832_ sky130_fd_sc_hd__xnor2_2
X_14574_ _04798_ _04800_ _04667_ net126 VGND VGND VPWR VPWR _04802_ sky130_fd_sc_hd__a211o_1
X_11786_ _01877_ _01878_ VGND VGND VPWR VPWR _01879_ sky130_fd_sc_hd__and2_1
XFILLER_0_94_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16313_ _06680_ _06684_ _06690_ VGND VGND VPWR VPWR _06691_ sky130_fd_sc_hd__or3b_1
XFILLER_0_126_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13525_ cla_inst.in2\[29\] _00205_ _00171_ cla_inst.in2\[30\] VGND VGND VPWR VPWR
+ _03655_ sky130_fd_sc_hd__a22o_1
XFILLER_0_12_34 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10737_ _08104_ _08093_ VGND VGND VPWR VPWR _00830_ sky130_fd_sc_hd__and2b_1
X_17293_ _07630_ _07332_ _07633_ _07631_ VGND VGND VPWR VPWR _07757_ sky130_fd_sc_hd__o31a_1
XFILLER_0_82_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_152_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16244_ _06467_ _06615_ VGND VGND VPWR VPWR _06616_ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13456_ _03180_ _03578_ _03048_ VGND VGND VPWR VPWR _03579_ sky130_fd_sc_hd__mux2_1
X_10668_ _00597_ _00760_ VGND VGND VPWR VPWR _00761_ sky130_fd_sc_hd__nand2_1
XFILLER_0_152_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12407_ _02485_ _02499_ VGND VGND VPWR VPWR _02500_ sky130_fd_sc_hd__or2b_1
XFILLER_0_113_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_752 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16175_ _06531_ _06535_ _06540_ VGND VGND VPWR VPWR _06541_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_140_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10599_ _00507_ _00528_ _00690_ _00691_ VGND VGND VPWR VPWR _00692_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_23_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13387_ _03495_ _03503_ VGND VGND VPWR VPWR _03504_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_51_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput107 net107 VGND VGND VPWR VPWR o_wb_data[31] sky130_fd_sc_hd__clkbuf_4
X_15126_ _05402_ _05403_ VGND VGND VPWR VPWR _05404_ sky130_fd_sc_hd__xor2_2
XFILLER_0_23_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12338_ _02426_ _02429_ VGND VGND VPWR VPWR _02431_ sky130_fd_sc_hd__and2b_1
XFILLER_0_105_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15057_ _05111_ _05221_ _05327_ VGND VGND VPWR VPWR _05328_ sky130_fd_sc_hd__a21bo_1
X_12269_ _07352_ _00563_ VGND VGND VPWR VPWR _02362_ sky130_fd_sc_hd__nand2_1
X_14008_ _00877_ _01678_ _04182_ VGND VGND VPWR VPWR _04183_ sky130_fd_sc_hd__nand3_1
XFILLER_0_37_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18816_ _09298_ _09321_ VGND VGND VPWR VPWR _09322_ sky130_fd_sc_hd__and2_1
X_18747_ _09267_ VGND VGND VPWR VPWR _00074_ sky130_fd_sc_hd__buf_1
X_15959_ _06304_ _06305_ VGND VGND VPWR VPWR _06306_ sky130_fd_sc_hd__or2_1
XFILLER_0_78_616 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09480_ cla_inst.in2\[16\] VGND VGND VPWR VPWR _03848_ sky130_fd_sc_hd__clkbuf_4
X_18678_ net39 _09189_ _09216_ VGND VGND VPWR VPWR _00049_ sky130_fd_sc_hd__o21a_1
XFILLER_0_78_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17629_ _08121_ _08122_ VGND VGND VPWR VPWR _08123_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_59_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_716 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_632 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_143_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09816_ cla_inst.in2\[29\] VGND VGND VPWR VPWR _07504_ sky130_fd_sc_hd__clkbuf_4
X_09747_ _06678_ VGND VGND VPWR VPWR _06754_ sky130_fd_sc_hd__inv_2
XTAP_2004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09678_ ApproximateM_inst.lob_16.lob2.genblk1\[7\].genblk1.mux.sel VGND VGND VPWR
+ VPWR _06008_ sky130_fd_sc_hd__buf_4
XFILLER_0_96_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_619 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11640_ _01633_ _01636_ _01731_ _01732_ VGND VGND VPWR VPWR _01733_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_65_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11571_ _00832_ _00439_ _01643_ _01644_ VGND VGND VPWR VPWR _01664_ sky130_fd_sc_hd__a22o_1
XFILLER_0_64_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13310_ _05224_ _08169_ _03417_ _03418_ VGND VGND VPWR VPWR _03419_ sky130_fd_sc_hd__and4_2
XFILLER_0_91_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10522_ _03728_ _05486_ VGND VGND VPWR VPWR _00615_ sky130_fd_sc_hd__nand2_1
XFILLER_0_134_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14290_ _04376_ VGND VGND VPWR VPWR _04491_ sky130_fd_sc_hd__inv_2
XFILLER_0_64_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_135_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_134_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10453_ _00125_ _00218_ _00178_ _00151_ VGND VGND VPWR VPWR _00546_ sky130_fd_sc_hd__a22oi_1
X_13241_ _03341_ _03342_ _00696_ _03204_ VGND VGND VPWR VPWR _03344_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_150_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10384_ _05736_ _08224_ VGND VGND VPWR VPWR _00477_ sky130_fd_sc_hd__nand2_1
X_13172_ _07504_ _00178_ _00147_ _00358_ VGND VGND VPWR VPWR _03271_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12123_ _06040_ _00194_ _02215_ VGND VGND VPWR VPWR _02216_ sky130_fd_sc_hd__a21oi_2
X_17980_ _08410_ _08504_ VGND VGND VPWR VPWR _08505_ sky130_fd_sc_hd__xor2_1
XFILLER_0_20_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12054_ _02023_ _02063_ _02064_ VGND VGND VPWR VPWR _02147_ sky130_fd_sc_hd__o21ai_1
X_16931_ _07356_ _07357_ _07360_ VGND VGND VPWR VPWR _07362_ sky130_fd_sc_hd__a21o_1
X_11005_ _04580_ _01064_ _01063_ _01066_ VGND VGND VPWR VPWR _01098_ sky130_fd_sc_hd__o2bb2a_1
X_16862_ _07196_ _07197_ VGND VGND VPWR VPWR _07287_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15813_ _04823_ _06140_ _06141_ _06142_ _06150_ VGND VGND VPWR VPWR _09371_ sky130_fd_sc_hd__a32o_1
X_18601_ _09097_ VGND VGND VPWR VPWR _09157_ sky130_fd_sc_hd__buf_2
X_16793_ _07209_ _07211_ VGND VGND VPWR VPWR _07212_ sky130_fd_sc_hd__xor2_1
X_18532_ net14 net17 net16 net19 VGND VGND VPWR VPWR _09102_ sky130_fd_sc_hd__or4_1
X_15744_ _05411_ _05415_ _05792_ _06075_ VGND VGND VPWR VPWR _06076_ sky130_fd_sc_hd__a211o_1
X_12956_ _03048_ VGND VGND VPWR VPWR _03049_ sky130_fd_sc_hd__clkbuf_4
X_18463_ _06425_ _06451_ _09028_ VGND VGND VPWR VPWR _09029_ sky130_fd_sc_hd__or3_1
X_11907_ _01987_ _01989_ _01988_ VGND VGND VPWR VPWR _02000_ sky130_fd_sc_hd__o21ai_1
X_15675_ _05998_ _05999_ _05912_ _05969_ VGND VGND VPWR VPWR _06001_ sky130_fd_sc_hd__a211o_1
XFILLER_0_114_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12887_ _00494_ VGND VGND VPWR VPWR _02980_ sky130_fd_sc_hd__buf_4
XTAP_2571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17414_ _06750_ _07623_ VGND VGND VPWR VPWR _07889_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14626_ _04855_ _04857_ VGND VGND VPWR VPWR _04858_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_74_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11838_ _01851_ _01930_ VGND VGND VPWR VPWR _01931_ sky130_fd_sc_hd__nor2_1
X_18394_ _08848_ _08899_ _08901_ VGND VGND VPWR VPWR _08954_ sky130_fd_sc_hd__o21ai_1
XTAP_1870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17345_ _02978_ _06999_ _02972_ VGND VGND VPWR VPWR _07814_ sky130_fd_sc_hd__o21ai_1
X_14557_ _00148_ _00149_ _06471_ _08452_ VGND VGND VPWR VPWR _04783_ sky130_fd_sc_hd__and4_1
XFILLER_0_16_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11769_ _08452_ VGND VGND VPWR VPWR _01862_ sky130_fd_sc_hd__clkinv_4
XFILLER_0_138_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13508_ _03632_ _03633_ _03634_ VGND VGND VPWR VPWR _03636_ sky130_fd_sc_hd__a21o_1
XFILLER_0_114_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17276_ _07629_ _07736_ _07737_ VGND VGND VPWR VPWR _07738_ sky130_fd_sc_hd__o21ai_1
X_14488_ _03377_ _07004_ cla_inst.in1\[24\] _03356_ VGND VGND VPWR VPWR _04707_ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19015_ clknet_4_9_0_clk _00000_ VGND VGND VPWR VPWR sel_op\[0\] sky130_fd_sc_hd__dfxtp_2
X_16227_ _02965_ _06418_ _06419_ VGND VGND VPWR VPWR _06597_ sky130_fd_sc_hd__a21o_1
X_13439_ _03152_ _03127_ VGND VGND VPWR VPWR _03560_ sky130_fd_sc_hd__or2_1
XFILLER_0_140_223 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16158_ _06518_ _06521_ _03313_ VGND VGND VPWR VPWR _06522_ sky130_fd_sc_hd__a21o_2
XFILLER_0_100_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15109_ _05367_ _05383_ VGND VGND VPWR VPWR _05385_ sky130_fd_sc_hd__or2_1
XFILLER_0_121_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16089_ _04900_ _06446_ VGND VGND VPWR VPWR _06447_ sky130_fd_sc_hd__and2_1
X_09601_ _04973_ _05148_ _05137_ VGND VGND VPWR VPWR _05170_ sky130_fd_sc_hd__a21oi_2
X_09532_ ApproximateM_inst.lob_16.lob2.genblk1\[12\].genblk1.mux.sel VGND VGND VPWR
+ VPWR _04416_ sky130_fd_sc_hd__buf_6
X_09463_ _03366_ VGND VGND VPWR VPWR _03662_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_58_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_579 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_733 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_131_256 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_112_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12810_ _02901_ _02902_ VGND VGND VPWR VPWR _02903_ sky130_fd_sc_hd__nor2_1
X_13790_ _03942_ _03943_ VGND VGND VPWR VPWR _03944_ sky130_fd_sc_hd__xor2_1
XFILLER_0_69_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12741_ _02777_ _02833_ VGND VGND VPWR VPWR _02834_ sky130_fd_sc_hd__xor2_2
XTAP_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15460_ _05760_ _05766_ VGND VGND VPWR VPWR _05767_ sky130_fd_sc_hd__or2_1
XTAP_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12672_ _02759_ _02760_ VGND VGND VPWR VPWR _02765_ sky130_fd_sc_hd__xor2_2
XFILLER_0_38_844 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14411_ _04610_ _04611_ _04621_ VGND VGND VPWR VPWR _04623_ sky130_fd_sc_hd__or3_1
XTAP_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11623_ _01713_ _01714_ _01715_ VGND VGND VPWR VPWR _01716_ sky130_fd_sc_hd__nand3_2
XFILLER_0_37_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15391_ _05690_ _05691_ VGND VGND VPWR VPWR _05692_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_154_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17130_ _02978_ _06843_ VGND VGND VPWR VPWR _07579_ sky130_fd_sc_hd__or2_1
X_14342_ _04420_ _04397_ _04546_ _04547_ VGND VGND VPWR VPWR _04549_ sky130_fd_sc_hd__a211o_4
X_11554_ _07232_ _07254_ _00439_ _04384_ VGND VGND VPWR VPWR _01647_ sky130_fd_sc_hd__nand4_2
XFILLER_0_52_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10505_ _00559_ _00574_ VGND VGND VPWR VPWR _00598_ sky130_fd_sc_hd__or2b_1
X_17061_ _07393_ _07399_ _07501_ VGND VGND VPWR VPWR _07503_ sky130_fd_sc_hd__and3_1
X_14273_ _04301_ _04311_ VGND VGND VPWR VPWR _04473_ sky130_fd_sc_hd__and2_1
X_11485_ _05595_ _04886_ _03815_ _05573_ VGND VGND VPWR VPWR _01578_ sky130_fd_sc_hd__a22o_1
XFILLER_0_69_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16012_ _06359_ _06360_ _06361_ VGND VGND VPWR VPWR _06363_ sky130_fd_sc_hd__a21bo_1
X_13224_ _00107_ _00166_ VGND VGND VPWR VPWR _03327_ sky130_fd_sc_hd__nand2_1
X_10436_ _00326_ _00331_ _00527_ _00528_ VGND VGND VPWR VPWR _00529_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_150_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13155_ _08724_ _08158_ _03250_ _03251_ VGND VGND VPWR VPWR _03253_ sky130_fd_sc_hd__a22o_1
X_10367_ _00459_ VGND VGND VPWR VPWR _00460_ sky130_fd_sc_hd__buf_4
XTAP_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12106_ _02197_ _02183_ _02187_ VGND VGND VPWR VPWR _02199_ sky130_fd_sc_hd__nand3_1
XTAP_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10298_ _00389_ _00390_ VGND VGND VPWR VPWR _00391_ sky130_fd_sc_hd__nor2_1
X_13086_ _03172_ _03177_ _03060_ VGND VGND VPWR VPWR _03178_ sky130_fd_sc_hd__mux2_1
X_17963_ _07207_ _07745_ _07859_ _06947_ VGND VGND VPWR VPWR _08487_ sky130_fd_sc_hd__a22o_1
X_12037_ _00845_ _02124_ _02125_ VGND VGND VPWR VPWR _02130_ sky130_fd_sc_hd__a21oi_2
X_16914_ _07342_ _07343_ VGND VGND VPWR VPWR _07344_ sky130_fd_sc_hd__xor2_1
X_17894_ _08410_ _08411_ VGND VGND VPWR VPWR _08412_ sky130_fd_sc_hd__or2_1
X_16845_ _02978_ _06617_ VGND VGND VPWR VPWR _07269_ sky130_fd_sc_hd__or2_1
X_16776_ _07111_ _07137_ VGND VGND VPWR VPWR _07193_ sky130_fd_sc_hd__or2_1
X_13988_ _04149_ _04150_ _04160_ VGND VGND VPWR VPWR _04161_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_88_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15727_ _06055_ _06056_ VGND VGND VPWR VPWR _06057_ sky130_fd_sc_hd__or2_1
X_18515_ _06246_ _06452_ VGND VGND VPWR VPWR _09084_ sky130_fd_sc_hd__or2_1
X_12939_ _03024_ _03031_ VGND VGND VPWR VPWR _03032_ sky130_fd_sc_hd__nand2_1
XFILLER_0_87_254 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15658_ _05980_ _05981_ VGND VGND VPWR VPWR _05982_ sky130_fd_sc_hd__nor2_1
X_18446_ _09007_ _09009_ VGND VGND VPWR VPWR _09010_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_146_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14609_ _01521_ _07015_ _04837_ _04838_ VGND VGND VPWR VPWR _04839_ sky130_fd_sc_hd__nand4_4
XFILLER_0_145_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18377_ _02992_ _06920_ _06921_ VGND VGND VPWR VPWR _08936_ sky130_fd_sc_hd__a21o_1
XFILLER_0_146_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15589_ _05905_ _05906_ VGND VGND VPWR VPWR _05907_ sky130_fd_sc_hd__nor2_1
XFILLER_0_145_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17328_ _07792_ _07794_ VGND VGND VPWR VPWR _07795_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_154_882 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_114_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17259_ _07607_ _07609_ _07610_ VGND VGND VPWR VPWR _07719_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_114_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09515_ _03454_ _04220_ VGND VGND VPWR VPWR _04231_ sky130_fd_sc_hd__and2_1
XFILLER_0_78_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09446_ ApproximateM_inst.lob_16.lob1.genblk1\[9\].genblk1.mux.sel VGND VGND VPWR
+ VPWR _03476_ sky130_fd_sc_hd__buf_4
XFILLER_0_78_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_162 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_117_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_144_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11270_ _01355_ _01361_ VGND VGND VPWR VPWR _01363_ sky130_fd_sc_hd__and2_1
X_10221_ _00310_ _00313_ VGND VGND VPWR VPWR _00314_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_120_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_574 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10152_ _00157_ _00232_ _00244_ VGND VGND VPWR VPWR _00245_ sky130_fd_sc_hd__o21ai_2
X_14960_ _05111_ _05221_ VGND VGND VPWR VPWR _05222_ sky130_fd_sc_hd__xnor2_1
X_10083_ ApproximateM_inst.lob_16.lob1.genblk1\[5\].genblk1.mux.sel VGND VGND VPWR
+ VPWR _00176_ sky130_fd_sc_hd__buf_4
X_13911_ _03147_ _03159_ _03061_ VGND VGND VPWR VPWR _04077_ sky130_fd_sc_hd__mux2_1
X_14891_ _00106_ _06094_ _05145_ _05146_ VGND VGND VPWR VPWR _05147_ sky130_fd_sc_hd__and4_1
X_16630_ _01005_ _03184_ _06871_ VGND VGND VPWR VPWR _07034_ sky130_fd_sc_hd__a21oi_2
X_13842_ _03983_ _03984_ _04000_ VGND VGND VPWR VPWR _04002_ sky130_fd_sc_hd__nor3_2
X_16561_ _06952_ _06958_ VGND VGND VPWR VPWR _06959_ sky130_fd_sc_hd__xor2_1
X_13773_ _03913_ _03926_ VGND VGND VPWR VPWR _03927_ sky130_fd_sc_hd__or2_2
XFILLER_0_57_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10985_ _01053_ _01077_ VGND VGND VPWR VPWR _01078_ sky130_fd_sc_hd__nor2_1
XFILLER_0_97_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15512_ _05767_ _05822_ VGND VGND VPWR VPWR _05824_ sky130_fd_sc_hd__xnor2_1
X_18300_ _08849_ _08850_ _08851_ VGND VGND VPWR VPWR _08852_ sky130_fd_sc_hd__and3_1
X_12724_ _02791_ _02816_ VGND VGND VPWR VPWR _02817_ sky130_fd_sc_hd__or2_1
XFILLER_0_128_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16492_ _06882_ _06883_ VGND VGND VPWR VPWR _06885_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_57_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18231_ _07650_ _07708_ VGND VGND VPWR VPWR _08777_ sky130_fd_sc_hd__nand2_1
X_15443_ _03000_ _05652_ _05748_ VGND VGND VPWR VPWR _05749_ sky130_fd_sc_hd__nand3_1
XFILLER_0_128_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12655_ _02747_ _02666_ VGND VGND VPWR VPWR _02748_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_72_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11606_ _01694_ _01697_ _01698_ VGND VGND VPWR VPWR _01699_ sky130_fd_sc_hd__or3b_1
X_18162_ _06368_ _07390_ VGND VGND VPWR VPWR _08703_ sky130_fd_sc_hd__nand2_1
XFILLER_0_154_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15374_ _05571_ _05629_ _05672_ _05673_ VGND VGND VPWR VPWR _05674_ sky130_fd_sc_hd__a211o_1
X_12586_ _07591_ _02676_ _02677_ _02678_ VGND VGND VPWR VPWR _02679_ sky130_fd_sc_hd__a22o_1
XFILLER_0_26_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17113_ _07556_ _07557_ _07560_ VGND VGND VPWR VPWR _07561_ sky130_fd_sc_hd__o21a_1
X_14325_ _04369_ _04372_ _04528_ VGND VGND VPWR VPWR _04530_ sky130_fd_sc_hd__and3_1
XFILLER_0_135_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11537_ _01625_ _01626_ _01629_ VGND VGND VPWR VPWR _01630_ sky130_fd_sc_hd__nand3_2
X_18093_ _08625_ _08627_ VGND VGND VPWR VPWR _08628_ sky130_fd_sc_hd__xor2_1
XFILLER_0_151_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_56 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17044_ _06756_ _07318_ VGND VGND VPWR VPWR _07485_ sky130_fd_sc_hd__or2_1
X_14256_ _04452_ _04453_ VGND VGND VPWR VPWR _04454_ sky130_fd_sc_hd__or2_1
X_11468_ _01551_ _01560_ VGND VGND VPWR VPWR _01561_ sky130_fd_sc_hd__xnor2_1
Xmax_cap128 _02383_ VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__buf_2
X_13207_ _00708_ _00707_ VGND VGND VPWR VPWR _03308_ sky130_fd_sc_hd__or2b_1
XFILLER_0_96_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10419_ _00510_ _00511_ VGND VGND VPWR VPWR _00512_ sky130_fd_sc_hd__or2_1
X_14187_ _04376_ _04377_ _04354_ VGND VGND VPWR VPWR _04379_ sky130_fd_sc_hd__a21oi_2
X_11399_ _01415_ _01454_ _01490_ _01491_ VGND VGND VPWR VPWR _01492_ sky130_fd_sc_hd__o211a_2
XTAP_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13138_ _03233_ _03234_ VGND VGND VPWR VPWR _03235_ sky130_fd_sc_hd__and2b_1
XTAP_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18995_ clknet_4_6_0_clk _09361_ VGND VGND VPWR VPWR salida\[48\] sky130_fd_sc_hd__dfxtp_1
XTAP_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13069_ _02983_ VGND VGND VPWR VPWR _03161_ sky130_fd_sc_hd__buf_4
X_17946_ _08359_ net132 _08466_ VGND VGND VPWR VPWR _08468_ sky130_fd_sc_hd__o21a_1
X_17877_ _08391_ _08392_ VGND VGND VPWR VPWR _08393_ sky130_fd_sc_hd__and2_1
X_16828_ _07248_ _07249_ VGND VGND VPWR VPWR _07250_ sky130_fd_sc_hd__or2b_1
XFILLER_0_88_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16759_ _07173_ _06420_ _07174_ VGND VGND VPWR VPWR _07175_ sky130_fd_sc_hd__and3_1
XFILLER_0_76_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_602 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18429_ _06408_ _08991_ VGND VGND VPWR VPWR _08992_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_114_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_80 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09995_ _09152_ _09158_ _09333_ VGND VGND VPWR VPWR _09338_ sky130_fd_sc_hd__nor3_4
XFILLER_0_79_530 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10770_ _00122_ _00862_ VGND VGND VPWR VPWR _00863_ sky130_fd_sc_hd__nand2_1
XFILLER_0_94_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09429_ _03239_ VGND VGND VPWR VPWR _03292_ sky130_fd_sc_hd__inv_2
XFILLER_0_109_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_739 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12440_ _05834_ VGND VGND VPWR VPWR _02533_ sky130_fd_sc_hd__buf_6
XFILLER_0_74_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12371_ _02397_ _02463_ VGND VGND VPWR VPWR _02464_ sky130_fd_sc_hd__nor2_1
XFILLER_0_151_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14110_ _04287_ _04293_ VGND VGND VPWR VPWR _04294_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_50_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11322_ _01312_ _01378_ _01413_ _01414_ VGND VGND VPWR VPWR _01415_ sky130_fd_sc_hd__a211oi_4
X_15090_ _05348_ _05349_ _05363_ VGND VGND VPWR VPWR _05364_ sky130_fd_sc_hd__o21a_1
X_14041_ _04169_ _04170_ _04216_ _04217_ VGND VGND VPWR VPWR _04219_ sky130_fd_sc_hd__o22a_1
X_11253_ _01254_ _01256_ _01255_ VGND VGND VPWR VPWR _01346_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_120_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10204_ _00295_ _00296_ VGND VGND VPWR VPWR _00297_ sky130_fd_sc_hd__and2b_1
X_11184_ _00777_ _00776_ VGND VGND VPWR VPWR _01277_ sky130_fd_sc_hd__and2b_1
X_17800_ _08307_ _08308_ VGND VGND VPWR VPWR _08309_ sky130_fd_sc_hd__nor2_1
X_10135_ _00226_ _00202_ _00209_ VGND VGND VPWR VPWR _00228_ sky130_fd_sc_hd__or3_1
X_18780_ _02988_ net43 _09276_ VGND VGND VPWR VPWR _09293_ sky130_fd_sc_hd__mux2_1
X_15992_ _03790_ _00207_ VGND VGND VPWR VPWR _06341_ sky130_fd_sc_hd__or2_1
X_10066_ _00157_ _00158_ VGND VGND VPWR VPWR _00159_ sky130_fd_sc_hd__or2_1
X_14943_ _05198_ _05202_ _05204_ VGND VGND VPWR VPWR _05205_ sky130_fd_sc_hd__o21a_1
X_17731_ _08230_ _08231_ _08233_ VGND VGND VPWR VPWR _08234_ sky130_fd_sc_hd__a21o_1
X_14874_ _05127_ VGND VGND VPWR VPWR _05129_ sky130_fd_sc_hd__inv_2
XFILLER_0_82_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17662_ _08155_ _08157_ VGND VGND VPWR VPWR _08159_ sky130_fd_sc_hd__xor2_1
X_13825_ _03981_ _03982_ _03786_ net189 VGND VGND VPWR VPWR _03983_ sky130_fd_sc_hd__a211oi_2
X_16613_ _03169_ _06464_ _06987_ _07016_ VGND VGND VPWR VPWR _09414_ sky130_fd_sc_hd__o2bb2a_2
X_17593_ _07979_ _07989_ _07987_ VGND VGND VPWR VPWR _08084_ sky130_fd_sc_hd__a21o_1
X_16544_ _06876_ _06885_ VGND VGND VPWR VPWR _06941_ sky130_fd_sc_hd__nand2_1
XFILLER_0_85_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13756_ _03906_ _03907_ _02980_ VGND VGND VPWR VPWR _03908_ sky130_fd_sc_hd__mux2_1
X_10968_ _01057_ _01060_ VGND VGND VPWR VPWR _01061_ sky130_fd_sc_hd__and2b_1
XFILLER_0_128_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12707_ _02762_ _02799_ VGND VGND VPWR VPWR _02800_ sky130_fd_sc_hd__xor2_2
X_16475_ _06828_ _06831_ VGND VGND VPWR VPWR _06866_ sky130_fd_sc_hd__and2b_1
X_13687_ _03811_ _03812_ _03831_ VGND VGND VPWR VPWR _03832_ sky130_fd_sc_hd__a21o_1
XFILLER_0_57_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10899_ _06008_ VGND VGND VPWR VPWR _00992_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_127_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15426_ _05634_ _05636_ _05728_ _05729_ VGND VGND VPWR VPWR _05730_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_66_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18214_ _08759_ _02871_ VGND VGND VPWR VPWR _08760_ sky130_fd_sc_hd__or2b_1
XFILLER_0_5_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12638_ _02727_ _02730_ VGND VGND VPWR VPWR _02731_ sky130_fd_sc_hd__nand2_1
XFILLER_0_122_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_603 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15357_ _00190_ _00192_ _07744_ _08224_ VGND VGND VPWR VPWR _05655_ sky130_fd_sc_hd__and4_1
X_18145_ _06598_ _08683_ _08684_ VGND VGND VPWR VPWR _08685_ sky130_fd_sc_hd__or3_1
X_12569_ _02654_ _02660_ _02661_ VGND VGND VPWR VPWR _02662_ sky130_fd_sc_hd__and3_1
XFILLER_0_108_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14308_ _04509_ _04510_ VGND VGND VPWR VPWR _04511_ sky130_fd_sc_hd__xor2_4
XFILLER_0_103_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18076_ _08513_ _08514_ _08512_ VGND VGND VPWR VPWR _08610_ sky130_fd_sc_hd__a21boi_2
X_15288_ _01505_ _00339_ VGND VGND VPWR VPWR _05580_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17027_ _01041_ _06364_ _06363_ VGND VGND VPWR VPWR _07467_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_22_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14239_ net201 _04433_ _04270_ _04271_ VGND VGND VPWR VPWR _04435_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_150_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09780_ _07102_ VGND VGND VPWR VPWR _07112_ sky130_fd_sc_hd__buf_6
XTAP_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18978_ clknet_4_3_0_clk _09410_ VGND VGND VPWR VPWR salida\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17929_ _08378_ _08379_ VGND VGND VPWR VPWR _08449_ sky130_fd_sc_hd__and2_1
XTAP_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_146_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09978_ _09212_ VGND VGND VPWR VPWR _09219_ sky130_fd_sc_hd__buf_4
X_11940_ _05638_ _03421_ _03607_ _00992_ VGND VGND VPWR VPWR _02033_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_98_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11871_ _07711_ _01962_ _01963_ VGND VGND VPWR VPWR _01964_ sky130_fd_sc_hd__and3_2
X_13610_ _03741_ _03746_ _02969_ VGND VGND VPWR VPWR _03748_ sky130_fd_sc_hd__a21oi_1
X_10822_ net169 _00772_ _00129_ net227 VGND VGND VPWR VPWR _00915_ sky130_fd_sc_hd__a22o_1
X_14590_ _04688_ _04689_ VGND VGND VPWR VPWR _04819_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13541_ _03649_ _03650_ _03670_ VGND VGND VPWR VPWR _03672_ sky130_fd_sc_hd__or3_4
XFILLER_0_95_875 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10753_ _00845_ VGND VGND VPWR VPWR _00846_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_27_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16260_ _01746_ _01503_ _03083_ _03166_ _06477_ _03161_ VGND VGND VPWR VPWR _06633_
+ sky130_fd_sc_hd__mux4_1
X_13472_ _03593_ _03594_ _03591_ _03592_ VGND VGND VPWR VPWR _03597_ sky130_fd_sc_hd__o211ai_2
X_10684_ _00771_ _00775_ _00769_ _00770_ VGND VGND VPWR VPWR _00777_ sky130_fd_sc_hd__o211a_1
X_15211_ _05494_ _05495_ VGND VGND VPWR VPWR _05496_ sky130_fd_sc_hd__xor2_2
XFILLER_0_124_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12423_ _02482_ VGND VGND VPWR VPWR _02516_ sky130_fd_sc_hd__inv_2
X_16191_ _03029_ _06464_ _06465_ _06557_ VGND VGND VPWR VPWR _09386_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_23_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15142_ _04254_ _04258_ _02780_ VGND VGND VPWR VPWR _05422_ sky130_fd_sc_hd__mux2_1
X_12354_ _02443_ _02444_ _02433_ _02441_ VGND VGND VPWR VPWR _02447_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_23_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_121_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11305_ _00846_ _00119_ _00121_ VGND VGND VPWR VPWR _01398_ sky130_fd_sc_hd__a21oi_2
X_15073_ _05227_ _05239_ _05226_ VGND VGND VPWR VPWR _05346_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_50_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12285_ _02264_ _02344_ _02377_ VGND VGND VPWR VPWR _02378_ sky130_fd_sc_hd__and3_1
XFILLER_0_121_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14024_ _04199_ _04200_ VGND VGND VPWR VPWR _04201_ sky130_fd_sc_hd__nor2_1
X_18901_ clknet_4_12_0_clk _00055_ VGND VGND VPWR VPWR cla_inst.in1\[19\] sky130_fd_sc_hd__dfxtp_2
X_11236_ _01315_ _01327_ _01316_ _01318_ VGND VGND VPWR VPWR _01329_ sky130_fd_sc_hd__nor4_1
X_18832_ net46 _03217_ _09331_ VGND VGND VPWR VPWR _09334_ sky130_fd_sc_hd__mux2_1
X_11167_ _01253_ _01259_ VGND VGND VPWR VPWR _01260_ sky130_fd_sc_hd__xnor2_1
X_10118_ _00210_ VGND VGND VPWR VPWR _00211_ sky130_fd_sc_hd__clkbuf_8
X_18763_ _09273_ _09280_ VGND VGND VPWR VPWR _09281_ sky130_fd_sc_hd__and2_1
X_11098_ _01189_ _01190_ VGND VGND VPWR VPWR _01191_ sky130_fd_sc_hd__xnor2_4
X_15975_ _06314_ _06320_ _06322_ VGND VGND VPWR VPWR _06323_ sky130_fd_sc_hd__a21oi_1
X_17714_ _08214_ _08215_ VGND VGND VPWR VPWR _08216_ sky130_fd_sc_hd__xnor2_1
X_14926_ _05184_ _05185_ VGND VGND VPWR VPWR _05186_ sky130_fd_sc_hd__xnor2_1
X_10049_ _00124_ _00137_ VGND VGND VPWR VPWR _00142_ sky130_fd_sc_hd__nand2_2
X_18694_ net47 _09189_ _09227_ VGND VGND VPWR VPWR _00056_ sky130_fd_sc_hd__o21a_1
XFILLER_0_117_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17645_ _08036_ VGND VGND VPWR VPWR _08141_ sky130_fd_sc_hd__clkbuf_4
X_14857_ _04034_ _03456_ _00665_ _02989_ VGND VGND VPWR VPWR _05110_ sky130_fd_sc_hd__a22oi_4
X_13808_ _03961_ _03962_ net236 _03931_ VGND VGND VPWR VPWR _03964_ sky130_fd_sc_hd__a211o_4
X_17576_ _08063_ _08064_ VGND VGND VPWR VPWR _08065_ sky130_fd_sc_hd__or2b_1
X_14788_ _05016_ _04917_ _05033_ VGND VGND VPWR VPWR _05035_ sky130_fd_sc_hd__nor3_1
XFILLER_0_19_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13739_ net121 _03885_ _03887_ VGND VGND VPWR VPWR _03889_ sky130_fd_sc_hd__o21a_1
XFILLER_0_73_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16527_ _06346_ _06790_ _06922_ _03086_ VGND VGND VPWR VPWR _06923_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16458_ _06469_ _06476_ _06498_ _06473_ _03079_ _03077_ VGND VGND VPWR VPWR _06848_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_5_302 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_143_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15409_ _05614_ _05618_ _05612_ VGND VGND VPWR VPWR _05712_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_6_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16389_ _06664_ _06772_ _06654_ VGND VGND VPWR VPWR _06773_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18128_ _08577_ _08580_ _08576_ VGND VGND VPWR VPWR _08666_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_112_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18059_ _06559_ _08590_ VGND VGND VPWR VPWR _08591_ sky130_fd_sc_hd__or2_1
XFILLER_0_41_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09901_ _03859_ _04121_ _04460_ _04482_ VGND VGND VPWR VPWR _08431_ sky130_fd_sc_hd__and4_1
XFILLER_0_6_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09832_ _07635_ _07646_ _07657_ _07668_ VGND VGND VPWR VPWR _07679_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_67_62 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09763_ _06863_ _06873_ _06917_ _06548_ VGND VGND VPWR VPWR _06928_ sky130_fd_sc_hd__o2bb2a_1
XTAP_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09694_ _05181_ _06149_ _06159_ _06170_ VGND VGND VPWR VPWR _06181_ sky130_fd_sc_hd__nand4_4
Xrebuffer10 _04094_ VGND VGND VPWR VPWR net173 sky130_fd_sc_hd__clkbuf_1
Xrebuffer21 _00305_ VGND VGND VPWR VPWR net184 sky130_fd_sc_hd__dlygate4sd1_1
XTAP_2208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer32 net194 VGND VGND VPWR VPWR net195 sky130_fd_sc_hd__buf_1
XTAP_2219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer43 _00772_ VGND VGND VPWR VPWR net206 sky130_fd_sc_hd__clkbuf_2
Xrebuffer54 _04681_ VGND VGND VPWR VPWR net217 sky130_fd_sc_hd__buf_1
XFILLER_0_95_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer65 net227 VGND VGND VPWR VPWR net228 sky130_fd_sc_hd__clkbuf_1
XTAP_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer76 _04003_ VGND VGND VPWR VPWR net239 sky130_fd_sc_hd__clkbuf_1
XTAP_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer87 _06560_ VGND VGND VPWR VPWR net334 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_146_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_355 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_146_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_889 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_452 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12070_ _02053_ _02162_ VGND VGND VPWR VPWR _02163_ sky130_fd_sc_hd__xnor2_1
X_11021_ _01113_ _06776_ VGND VGND VPWR VPWR _01114_ sky130_fd_sc_hd__nor2_4
XFILLER_0_99_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15760_ _03015_ _03072_ VGND VGND VPWR VPWR _06092_ sky130_fd_sc_hd__nand2_1
X_12972_ _09263_ _03064_ _03024_ VGND VGND VPWR VPWR _03065_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_99_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14711_ _04410_ _04947_ _04950_ VGND VGND VPWR VPWR _04951_ sky130_fd_sc_hd__a21o_1
X_11923_ _02011_ _02015_ VGND VGND VPWR VPWR _02016_ sky130_fd_sc_hd__and2_1
X_15691_ _06015_ _06016_ _04823_ VGND VGND VPWR VPWR _06018_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_99_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14642_ _04872_ _04874_ VGND VGND VPWR VPWR _04876_ sky130_fd_sc_hd__or2_1
X_17430_ _02589_ _02844_ _02587_ VGND VGND VPWR VPWR _07906_ sky130_fd_sc_hd__o21ba_1
XTAP_2764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11854_ ApproximateM_inst.lob_16.lob2.genblk1\[3\].genblk1.mux.sel ApproximateM_inst.lob_16.lob1.genblk1\[12\].genblk1.mux.sel
+ _03826_ ApproximateM_inst.lob_16.lob2.genblk1\[4\].genblk1.mux.sel VGND VGND VPWR
+ VPWR _01947_ sky130_fd_sc_hd__a22o_1
XFILLER_0_67_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10805_ _00893_ _00895_ _00897_ VGND VGND VPWR VPWR _00898_ sky130_fd_sc_hd__nand3_2
X_14573_ _04667_ net126 _04798_ _04800_ VGND VGND VPWR VPWR _04801_ sky130_fd_sc_hd__o211ai_4
X_17361_ net331 _07706_ VGND VGND VPWR VPWR _07830_ sky130_fd_sc_hd__nor2_1
XFILLER_0_67_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11785_ _01508_ _01513_ VGND VGND VPWR VPWR _01878_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_28_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13524_ cla_inst.in2\[30\] cla_inst.in2\[29\] _00205_ _00171_ VGND VGND VPWR VPWR
+ _03654_ sky130_fd_sc_hd__and4_1
X_16312_ _06687_ _06597_ _06688_ VGND VGND VPWR VPWR _06690_ sky130_fd_sc_hd__or3_1
X_10736_ _00827_ _00828_ VGND VGND VPWR VPWR _00829_ sky130_fd_sc_hd__nand2_1
X_17292_ _07753_ _07754_ VGND VGND VPWR VPWR _07756_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_55_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16243_ _06612_ _06614_ _02982_ VGND VGND VPWR VPWR _06615_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13455_ _03187_ VGND VGND VPWR VPWR _03578_ sky130_fd_sc_hd__inv_2
X_10667_ _00594_ _00596_ VGND VGND VPWR VPWR _00760_ sky130_fd_sc_hd__nand2_1
XFILLER_0_125_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12406_ _02491_ _02498_ VGND VGND VPWR VPWR _02499_ sky130_fd_sc_hd__or2b_1
XFILLER_0_35_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16174_ _06536_ _06538_ _06539_ _03313_ _06520_ VGND VGND VPWR VPWR _06540_ sky130_fd_sc_hd__a2111o_1
X_13386_ _03496_ _03502_ VGND VGND VPWR VPWR _03503_ sky130_fd_sc_hd__xor2_1
XFILLER_0_3_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10598_ _00688_ _00689_ _00482_ _00487_ VGND VGND VPWR VPWR _00691_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_2_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15125_ _03368_ _03067_ _05278_ _05276_ VGND VGND VPWR VPWR _05403_ sky130_fd_sc_hd__a31o_1
Xoutput108 net108 VGND VGND VPWR VPWR o_wb_data[3] sky130_fd_sc_hd__clkbuf_4
X_12337_ _02426_ _02429_ VGND VGND VPWR VPWR _02430_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_51_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15056_ _05219_ _05220_ VGND VGND VPWR VPWR _05327_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12268_ _02357_ _02360_ VGND VGND VPWR VPWR _02361_ sky130_fd_sc_hd__nor2_1
X_14007_ _04180_ _04181_ VGND VGND VPWR VPWR _04182_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_120_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11219_ net220 _01020_ _01310_ _01311_ VGND VGND VPWR VPWR _01312_ sky130_fd_sc_hd__o211ai_4
X_12199_ _02288_ _02289_ _02203_ VGND VGND VPWR VPWR _02292_ sky130_fd_sc_hd__a21oi_1
Xoutput90 net90 VGND VGND VPWR VPWR o_wb_data[16] sky130_fd_sc_hd__clkbuf_4
X_18815_ _03016_ net55 _09301_ VGND VGND VPWR VPWR _09321_ sky130_fd_sc_hd__mux2_1
X_18746_ _09245_ _09266_ VGND VGND VPWR VPWR _09267_ sky130_fd_sc_hd__and2_1
X_15958_ _06272_ _06280_ _06278_ VGND VGND VPWR VPWR _06305_ sky130_fd_sc_hd__o21ai_1
X_14909_ _05165_ _05166_ VGND VGND VPWR VPWR _05167_ sky130_fd_sc_hd__xnor2_1
X_18677_ _02127_ _09190_ _09191_ VGND VGND VPWR VPWR _09216_ sky130_fd_sc_hd__a21oi_1
X_15889_ _06183_ _06225_ VGND VGND VPWR VPWR _06231_ sky130_fd_sc_hd__or2_1
X_17628_ _08016_ _08018_ _08014_ VGND VGND VPWR VPWR _08122_ sky130_fd_sc_hd__o21ba_1
X_17559_ _06655_ _07825_ VGND VGND VPWR VPWR _08046_ sky130_fd_sc_hd__nand2_1
XFILLER_0_129_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09815_ _07472_ _07210_ _07319_ VGND VGND VPWR VPWR _07493_ sky130_fd_sc_hd__nand3_2
X_09746_ _06678_ _06700_ _06711_ _06732_ VGND VGND VPWR VPWR _06743_ sky130_fd_sc_hd__and4b_1
XTAP_2005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09677_ _05747_ _05986_ VGND VGND VPWR VPWR _05997_ sky130_fd_sc_hd__nand2_2
XTAP_2016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11570_ _04056_ net204 _01660_ _01662_ VGND VGND VPWR VPWR _01663_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_119_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10521_ _00443_ _00612_ _00613_ VGND VGND VPWR VPWR _00614_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_52_539 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13240_ _00696_ _03204_ _03341_ _03342_ VGND VGND VPWR VPWR _03343_ sky130_fd_sc_hd__o211a_1
XFILLER_0_150_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10452_ _07526_ _00132_ _00360_ _00359_ _07570_ VGND VGND VPWR VPWR _00545_ sky130_fd_sc_hd__a32o_1
XFILLER_0_33_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13171_ _09166_ _09172_ _00178_ _00181_ VGND VGND VPWR VPWR _03270_ sky130_fd_sc_hd__and4_1
X_10383_ _00474_ _00475_ VGND VGND VPWR VPWR _00476_ sky130_fd_sc_hd__xor2_1
XFILLER_0_0_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12122_ _06051_ _00172_ VGND VGND VPWR VPWR _02215_ sky130_fd_sc_hd__and2_1
XFILLER_0_103_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12053_ _02144_ _02145_ VGND VGND VPWR VPWR _02146_ sky130_fd_sc_hd__and2_1
X_16930_ _07356_ _07357_ _07360_ VGND VGND VPWR VPWR _07361_ sky130_fd_sc_hd__nand3_1
X_11004_ _01094_ _01096_ VGND VGND VPWR VPWR _01097_ sky130_fd_sc_hd__nand2_2
X_16861_ _06937_ _07130_ VGND VGND VPWR VPWR _07285_ sky130_fd_sc_hd__nor2_1
X_18600_ net265 _09140_ _09156_ _09144_ VGND VGND VPWR VPWR _00023_ sky130_fd_sc_hd__o211a_1
X_15812_ _03121_ _06148_ VGND VGND VPWR VPWR _06150_ sky130_fd_sc_hd__nand2_1
X_16792_ _07018_ _06875_ VGND VGND VPWR VPWR _07211_ sky130_fd_sc_hd__nor2_1
X_18531_ net18 net21 net20 net22 VGND VGND VPWR VPWR _09100_ sky130_fd_sc_hd__or4b_1
X_15743_ _05948_ _05875_ _05947_ _06015_ VGND VGND VPWR VPWR _06075_ sky130_fd_sc_hd__or4_1
X_12955_ _03047_ VGND VGND VPWR VPWR _03048_ sky130_fd_sc_hd__clkbuf_4
X_11906_ _01997_ _01998_ VGND VGND VPWR VPWR _01999_ sky130_fd_sc_hd__or2_1
X_18462_ _06408_ _06449_ _03073_ VGND VGND VPWR VPWR _09028_ sky130_fd_sc_hd__a21oi_1
X_15674_ _05912_ _05969_ _05998_ _05999_ VGND VGND VPWR VPWR _06000_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_87_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12886_ _02978_ VGND VGND VPWR VPWR _02979_ sky130_fd_sc_hd__clkbuf_4
XTAP_2550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17413_ _07885_ _07887_ VGND VGND VPWR VPWR _07888_ sky130_fd_sc_hd__nor2_1
XFILLER_0_56_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14625_ _04725_ _03455_ _04856_ VGND VGND VPWR VPWR _04857_ sky130_fd_sc_hd__and3_1
X_11837_ _06711_ _04045_ _01929_ _01850_ VGND VGND VPWR VPWR _01930_ sky130_fd_sc_hd__a22oi_1
X_18393_ _08950_ _08952_ VGND VGND VPWR VPWR _08953_ sky130_fd_sc_hd__xor2_1
XTAP_2594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14556_ _03321_ _06471_ _04591_ _03322_ VGND VGND VPWR VPWR _04782_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_23_78 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17344_ _06696_ _06701_ _06703_ _06707_ _03061_ _03079_ VGND VGND VPWR VPWR _07813_
+ sky130_fd_sc_hd__mux4_1
X_11768_ _01859_ _01860_ VGND VGND VPWR VPWR _01861_ sky130_fd_sc_hd__nand2_1
XFILLER_0_138_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13507_ _03632_ _03633_ _03634_ VGND VGND VPWR VPWR _03635_ sky130_fd_sc_hd__nand3_1
XFILLER_0_15_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10719_ _08060_ VGND VGND VPWR VPWR _00812_ sky130_fd_sc_hd__inv_2
X_14487_ _01521_ _07962_ _04568_ _04570_ VGND VGND VPWR VPWR _04706_ sky130_fd_sc_hd__and4_1
XFILLER_0_70_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17275_ _07637_ _07638_ VGND VGND VPWR VPWR _07737_ sky130_fd_sc_hd__or2_1
X_11699_ _01764_ _01765_ _01767_ VGND VGND VPWR VPWR _01792_ sky130_fd_sc_hd__nor3b_1
XFILLER_0_130_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19014_ clknet_4_3_0_clk _00104_ VGND VGND VPWR VPWR op_code\[3\] sky130_fd_sc_hd__dfxtp_4
XFILLER_0_113_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13438_ _03532_ _03559_ VGND VGND VPWR VPWR _09377_ sky130_fd_sc_hd__nand2_1
X_16226_ _02784_ _06333_ _03030_ VGND VGND VPWR VPWR _06596_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_125_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xrebuffer1 _00694_ VGND VGND VPWR VPWR net164 sky130_fd_sc_hd__buf_1
XFILLER_0_70_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16157_ _03281_ _06519_ _06520_ VGND VGND VPWR VPWR _06521_ sky130_fd_sc_hd__a21o_1
XFILLER_0_140_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13369_ _03482_ _03483_ VGND VGND VPWR VPWR _03484_ sky130_fd_sc_hd__nand2_1
XFILLER_0_51_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15108_ _05367_ _05383_ VGND VGND VPWR VPWR _05384_ sky130_fd_sc_hd__nand2_1
X_16088_ _03052_ _04647_ _06445_ VGND VGND VPWR VPWR _06446_ sky130_fd_sc_hd__and3_1
X_15039_ _02976_ _03039_ _05306_ _05307_ _05308_ VGND VGND VPWR VPWR _05309_ sky130_fd_sc_hd__o32a_1
XFILLER_0_139_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09600_ _04973_ _05137_ _05148_ VGND VGND VPWR VPWR _05159_ sky130_fd_sc_hd__and3_1
XFILLER_0_64_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09531_ _04351_ _04373_ _04384_ _04395_ VGND VGND VPWR VPWR _04406_ sky130_fd_sc_hd__and4_4
X_18729_ _09253_ VGND VGND VPWR VPWR _00068_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09462_ _03531_ VGND VGND VPWR VPWR _03651_ sky130_fd_sc_hd__buf_8
XFILLER_0_19_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_514 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_132_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_666 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09729_ _05006_ _05104_ VGND VGND VPWR VPWR _06558_ sky130_fd_sc_hd__or2b_1
XFILLER_0_69_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12740_ _02801_ _02831_ _02832_ VGND VGND VPWR VPWR _02833_ sky130_fd_sc_hd__a21o_1
XTAP_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12671_ _08865_ _01357_ VGND VGND VPWR VPWR _02764_ sky130_fd_sc_hd__nand2_1
XTAP_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14410_ _04610_ _04611_ _04621_ VGND VGND VPWR VPWR _04622_ sky130_fd_sc_hd__o21ai_1
XTAP_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_856 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11622_ _01625_ _01630_ VGND VGND VPWR VPWR _01715_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15390_ _05536_ _05547_ _05534_ VGND VGND VPWR VPWR _05691_ sky130_fd_sc_hd__a21oi_2
XTAP_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_108_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14341_ _04544_ _04545_ _04350_ _04422_ VGND VGND VPWR VPWR _04547_ sky130_fd_sc_hd__o211a_1
X_11553_ _01643_ _01645_ VGND VGND VPWR VPWR _01646_ sky130_fd_sc_hd__nand2_2
XFILLER_0_53_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10504_ _00594_ _00596_ VGND VGND VPWR VPWR _00597_ sky130_fd_sc_hd__or2_1
X_17060_ _07393_ _07399_ _07501_ VGND VGND VPWR VPWR _07502_ sky130_fd_sc_hd__a21oi_1
X_14272_ _04468_ _04469_ _04299_ _04428_ VGND VGND VPWR VPWR _04472_ sky130_fd_sc_hd__a211o_2
XFILLER_0_123_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11484_ _05573_ _05595_ _04886_ _03815_ VGND VGND VPWR VPWR _01577_ sky130_fd_sc_hd__and4_1
XFILLER_0_150_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16011_ _00644_ _00248_ VGND VGND VPWR VPWR _06361_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13223_ _03323_ _03325_ VGND VGND VPWR VPWR _03326_ sky130_fd_sc_hd__nor2_1
X_10435_ _00507_ _00508_ _00526_ VGND VGND VPWR VPWR _00528_ sky130_fd_sc_hd__nor3_4
XFILLER_0_111_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13154_ _08724_ _08158_ _03250_ _03251_ VGND VGND VPWR VPWR _03252_ sky130_fd_sc_hd__nand4_4
X_10366_ _06613_ VGND VGND VPWR VPWR _00459_ sky130_fd_sc_hd__clkbuf_8
XTAP_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12105_ _02183_ _02187_ _02197_ VGND VGND VPWR VPWR _02198_ sky130_fd_sc_hd__a21o_1
XTAP_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13085_ _03174_ _03176_ _03047_ VGND VGND VPWR VPWR _03177_ sky130_fd_sc_hd__mux2_1
X_17962_ _08367_ _08375_ _08373_ VGND VGND VPWR VPWR _08486_ sky130_fd_sc_hd__a21o_1
X_10297_ cla_inst.in2\[25\] _00172_ _00387_ _00388_ VGND VGND VPWR VPWR _00390_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_20_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12036_ _02126_ _02128_ VGND VGND VPWR VPWR _02129_ sky130_fd_sc_hd__and2_1
X_16913_ _07233_ _07234_ _07237_ VGND VGND VPWR VPWR _07343_ sky130_fd_sc_hd__a21o_1
X_17893_ _08314_ _08347_ _08408_ VGND VGND VPWR VPWR _08411_ sky130_fd_sc_hd__and3_1
X_16844_ _03912_ _06629_ _07267_ VGND VGND VPWR VPWR _07268_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_18_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16775_ _07152_ _07153_ VGND VGND VPWR VPWR _07192_ sky130_fd_sc_hd__and2b_1
X_13987_ _04158_ _04159_ VGND VGND VPWR VPWR _04160_ sky130_fd_sc_hd__and2_1
XFILLER_0_87_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18514_ _06248_ _06414_ _09076_ VGND VGND VPWR VPWR _09083_ sky130_fd_sc_hd__or3b_1
X_15726_ _05917_ _06054_ VGND VGND VPWR VPWR _06056_ sky130_fd_sc_hd__nor2_1
X_12938_ _03027_ _01746_ _03030_ VGND VGND VPWR VPWR _03031_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_75_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18445_ _08961_ _09008_ VGND VGND VPWR VPWR _09009_ sky130_fd_sc_hd__nor2_1
XFILLER_0_34_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15657_ _05978_ _05979_ _05973_ VGND VGND VPWR VPWR _05981_ sky130_fd_sc_hd__a21oi_1
XTAP_2380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12869_ _02958_ _02960_ _02961_ VGND VGND VPWR VPWR _02962_ sky130_fd_sc_hd__a21oi_2
XTAP_2391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14608_ _03651_ _03596_ cla_inst.in1\[27\] _07112_ VGND VGND VPWR VPWR _04838_ sky130_fd_sc_hd__nand4_4
X_18376_ _03068_ _06448_ VGND VGND VPWR VPWR _08935_ sky130_fd_sc_hd__nor2_1
XFILLER_0_141_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15588_ _05903_ _05904_ _05815_ _05817_ VGND VGND VPWR VPWR _05906_ sky130_fd_sc_hd__o211a_1
XTAP_1690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_145_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17327_ _07671_ _07558_ _07670_ _07793_ VGND VGND VPWR VPWR _07794_ sky130_fd_sc_hd__o31a_4
X_14539_ _01504_ _06094_ VGND VGND VPWR VPWR _04763_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17258_ _07705_ _07717_ VGND VGND VPWR VPWR _07718_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_113_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16209_ _06574_ _06576_ _03324_ VGND VGND VPWR VPWR _06577_ sky130_fd_sc_hd__a21o_1
X_17189_ _07619_ _07642_ VGND VGND VPWR VPWR _07643_ sky130_fd_sc_hd__xor2_1
XFILLER_0_11_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09514_ ApproximateM_inst.lob_16.lob1.genblk1\[7\].genblk1.mux.sel VGND VGND VPWR
+ VPWR _04220_ sky130_fd_sc_hd__buf_6
XFILLER_0_149_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09445_ _03454_ VGND VGND VPWR VPWR _03465_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_91_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_620 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_667 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_144_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_596 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_870 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10220_ _00311_ _00312_ VGND VGND VPWR VPWR _00313_ sky130_fd_sc_hd__and2b_1
XFILLER_0_30_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10151_ _00233_ _00243_ VGND VGND VPWR VPWR _00244_ sky130_fd_sc_hd__xor2_1
XFILLER_0_100_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10082_ _00174_ VGND VGND VPWR VPWR _00175_ sky130_fd_sc_hd__clkbuf_4
X_13910_ _02978_ _04075_ VGND VGND VPWR VPWR _04076_ sky130_fd_sc_hd__nor2_1
X_14890_ _00148_ _00149_ _00459_ _05845_ VGND VGND VPWR VPWR _05146_ sky130_fd_sc_hd__nand4_2
XFILLER_0_89_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13841_ _03985_ _03999_ VGND VGND VPWR VPWR _04000_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_97_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16560_ _06522_ _06525_ _06957_ _00515_ VGND VGND VPWR VPWR _06958_ sky130_fd_sc_hd__a211o_1
X_13772_ _03033_ _03924_ _03099_ VGND VGND VPWR VPWR _03926_ sky130_fd_sc_hd__mux2_1
X_10984_ _01053_ _01074_ _01075_ _01076_ VGND VGND VPWR VPWR _01077_ sky130_fd_sc_hd__and4b_1
XFILLER_0_85_704 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15511_ _05811_ _05821_ VGND VGND VPWR VPWR _05822_ sky130_fd_sc_hd__xor2_1
XFILLER_0_139_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12723_ _02789_ _02815_ VGND VGND VPWR VPWR _02816_ sky130_fd_sc_hd__nor2_1
XFILLER_0_139_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16491_ _06578_ _06816_ VGND VGND VPWR VPWR _06883_ sky130_fd_sc_hd__nor2_1
XFILLER_0_84_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18230_ _08774_ _08775_ VGND VGND VPWR VPWR _08776_ sky130_fd_sc_hd__nand2_1
X_15442_ _05745_ _05746_ VGND VGND VPWR VPWR _05748_ sky130_fd_sc_hd__xnor2_1
X_12654_ _02611_ _02654_ VGND VGND VPWR VPWR _02747_ sky130_fd_sc_hd__or2_1
XFILLER_0_154_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11605_ _07853_ _01695_ _01696_ _01673_ VGND VGND VPWR VPWR _01698_ sky130_fd_sc_hd__a31o_2
XFILLER_0_26_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18161_ _08699_ _08700_ VGND VGND VPWR VPWR _08701_ sky130_fd_sc_hd__and2b_1
XFILLER_0_143_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15373_ _05651_ _05670_ VGND VGND VPWR VPWR _05673_ sky130_fd_sc_hd__and2_1
X_12585_ _07243_ ApproximateM_inst.lob_16.lob1.genblk1\[1\].genblk1.mux.sel ApproximateM_inst.lob_16.lob1.mux.sel
+ _07221_ VGND VGND VPWR VPWR _02678_ sky130_fd_sc_hd__a22o_1
XFILLER_0_136_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17112_ _06559_ _07558_ VGND VGND VPWR VPWR _07560_ sky130_fd_sc_hd__nor2_1
X_14324_ _04369_ _04372_ _04528_ VGND VGND VPWR VPWR _04529_ sky130_fd_sc_hd__a21oi_2
X_11536_ _01627_ _01628_ VGND VGND VPWR VPWR _01629_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_53_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18092_ _07332_ _08260_ _08459_ VGND VGND VPWR VPWR _08627_ sky130_fd_sc_hd__or3_1
XFILLER_0_135_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_151_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14255_ _06460_ _00502_ _04450_ _04451_ VGND VGND VPWR VPWR _04453_ sky130_fd_sc_hd__o2bb2a_1
X_17043_ _07392_ _07404_ VGND VGND VPWR VPWR _07484_ sky130_fd_sc_hd__or2b_1
XFILLER_0_150_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap118 _05863_ VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__buf_1
X_11467_ _01556_ _01559_ VGND VGND VPWR VPWR _01560_ sky130_fd_sc_hd__xor2_1
XFILLER_0_1_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap129 _02293_ VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__buf_1
XFILLER_0_111_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13206_ _03305_ _03306_ VGND VGND VPWR VPWR _03307_ sky130_fd_sc_hd__nand2_1
XFILLER_0_110_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10418_ cla_inst.in2\[31\] _07700_ _00509_ _07559_ VGND VGND VPWR VPWR _00511_ sky130_fd_sc_hd__and4_1
XFILLER_0_110_216 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14186_ _04354_ _04376_ _04377_ VGND VGND VPWR VPWR _04378_ sky130_fd_sc_hd__and3_2
X_11398_ _01468_ _01489_ _01488_ VGND VGND VPWR VPWR _01491_ sky130_fd_sc_hd__a21o_1
XTAP_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13137_ _03231_ _03232_ _03227_ VGND VGND VPWR VPWR _03234_ sky130_fd_sc_hd__a21o_1
XTAP_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10349_ _03793_ _00440_ _00441_ VGND VGND VPWR VPWR _00442_ sky130_fd_sc_hd__a21bo_1
X_18994_ clknet_4_0_0_clk _09360_ VGND VGND VPWR VPWR salida\[47\] sky130_fd_sc_hd__dfxtp_1
XTAP_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13068_ _03159_ VGND VGND VPWR VPWR _03160_ sky130_fd_sc_hd__inv_2
X_17945_ _08359_ net132 _08466_ VGND VGND VPWR VPWR _08467_ sky130_fd_sc_hd__nor3_1
X_12019_ _05562_ _05584_ _04220_ _04242_ VGND VGND VPWR VPWR _02112_ sky130_fd_sc_hd__and4_1
X_17876_ _08389_ _08390_ VGND VGND VPWR VPWR _08392_ sky130_fd_sc_hd__or2_1
XFILLER_0_136_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16827_ _07191_ _07192_ _07247_ VGND VGND VPWR VPWR _07249_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_45_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_520 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16758_ _07172_ _06355_ _06354_ VGND VGND VPWR VPWR _07174_ sky130_fd_sc_hd__a21o_1
X_15709_ _01417_ _00665_ VGND VGND VPWR VPWR _06037_ sky130_fd_sc_hd__and2_1
XFILLER_0_76_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16689_ _07096_ _07097_ _07098_ VGND VGND VPWR VPWR _07099_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_146_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18428_ _03016_ _06592_ _06551_ VGND VGND VPWR VPWR _08991_ sky130_fd_sc_hd__a21o_1
XFILLER_0_119_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_89 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18359_ _08862_ _08894_ _08914_ VGND VGND VPWR VPWR _08916_ sky130_fd_sc_hd__or3_1
XFILLER_0_145_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_840 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09994_ _09152_ _09158_ _09333_ VGND VGND VPWR VPWR _09337_ sky130_fd_sc_hd__o21a_2
XFILLER_0_79_542 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_149_452 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09428_ sel_op\[1\] VGND VGND VPWR VPWR _03281_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_94_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_125_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12370_ _02311_ _02396_ _02392_ _02395_ VGND VGND VPWR VPWR _02463_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_22_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11321_ _01394_ _01395_ _01412_ VGND VGND VPWR VPWR _01414_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_132_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_120_503 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_132_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14040_ _04169_ _04170_ _04216_ _04217_ VGND VGND VPWR VPWR _04218_ sky130_fd_sc_hd__nor4_2
XFILLER_0_133_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11252_ _00169_ _00131_ _01342_ _01343_ VGND VGND VPWR VPWR _01345_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_132_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10203_ _00294_ _05322_ _05333_ _04504_ VGND VGND VPWR VPWR _00296_ sky130_fd_sc_hd__a22o_1
X_11183_ _00965_ _00961_ VGND VGND VPWR VPWR _01276_ sky130_fd_sc_hd__or2b_4
XFILLER_0_101_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10134_ _00202_ _00209_ _00226_ VGND VGND VPWR VPWR _00227_ sky130_fd_sc_hd__o21a_1
X_15991_ _03790_ _00207_ VGND VGND VPWR VPWR _06339_ sky130_fd_sc_hd__and2_1
X_17730_ _08025_ _08026_ _08132_ _08232_ VGND VGND VPWR VPWR _08233_ sky130_fd_sc_hd__a31o_1
X_10065_ _08202_ _00143_ _00156_ VGND VGND VPWR VPWR _00158_ sky130_fd_sc_hd__nor3_1
X_14942_ _05198_ _05202_ _04238_ VGND VGND VPWR VPWR _05204_ sky130_fd_sc_hd__a21oi_1
X_17661_ _08156_ _08051_ _08048_ VGND VGND VPWR VPWR _08157_ sky130_fd_sc_hd__a21o_1
X_14873_ _05125_ _05888_ _07635_ _05127_ VGND VGND VPWR VPWR _05128_ sky130_fd_sc_hd__and4b_1
X_16612_ _06992_ _06994_ _07011_ _07014_ VGND VGND VPWR VPWR _07016_ sky130_fd_sc_hd__a211o_1
X_13824_ _03963_ _03964_ _03980_ VGND VGND VPWR VPWR _03982_ sky130_fd_sc_hd__nand3_2
X_17592_ _08079_ _08081_ VGND VGND VPWR VPWR _08083_ sky130_fd_sc_hd__xor2_1
XFILLER_0_106_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16543_ _06937_ _06766_ VGND VGND VPWR VPWR _06940_ sky130_fd_sc_hd__nor2_1
X_10967_ _01058_ _01059_ VGND VGND VPWR VPWR _01060_ sky130_fd_sc_hd__xnor2_4
X_13755_ _03110_ _03113_ _03090_ VGND VGND VPWR VPWR _03907_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12706_ _02774_ _02773_ VGND VGND VPWR VPWR _02799_ sky130_fd_sc_hd__and2b_1
X_16474_ _03166_ _06464_ _06865_ VGND VGND VPWR VPWR _09412_ sky130_fd_sc_hd__a21oi_2
X_13686_ _03814_ _03830_ VGND VGND VPWR VPWR _03831_ sky130_fd_sc_hd__xnor2_1
X_10898_ _05682_ _05388_ VGND VGND VPWR VPWR _00991_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18213_ _02172_ _02470_ _02851_ VGND VGND VPWR VPWR _08759_ sky130_fd_sc_hd__nor3_1
X_15425_ _05720_ _05727_ VGND VGND VPWR VPWR _05729_ sky130_fd_sc_hd__nor2_1
XFILLER_0_116_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12637_ _02600_ _02729_ VGND VGND VPWR VPWR _02730_ sky130_fd_sc_hd__nor2_1
XFILLER_0_31_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18144_ _08682_ _06397_ _06396_ VGND VGND VPWR VPWR _08684_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_5_539 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15356_ _02996_ _00339_ _09059_ _02993_ VGND VGND VPWR VPWR _05654_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_53_453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12568_ _02534_ _02537_ VGND VGND VPWR VPWR _02661_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_108_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14307_ _01873_ _03044_ VGND VGND VPWR VPWR _04510_ sky130_fd_sc_hd__nand2_2
X_11519_ _04690_ _03673_ _01172_ _01173_ VGND VGND VPWR VPWR _01612_ sky130_fd_sc_hd__a22o_1
XFILLER_0_151_650 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18075_ _08607_ _08608_ VGND VGND VPWR VPWR _08609_ sky130_fd_sc_hd__nand2_1
X_15287_ _05577_ _05578_ VGND VGND VPWR VPWR _05579_ sky130_fd_sc_hd__nor2_1
X_12499_ _02582_ _02591_ VGND VGND VPWR VPWR _02592_ sky130_fd_sc_hd__or2_1
XFILLER_0_111_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17026_ _01041_ _06363_ _06364_ VGND VGND VPWR VPWR _07466_ sky130_fd_sc_hd__and3_1
X_14238_ _04270_ _04271_ net200 _04433_ VGND VGND VPWR VPWR _04434_ sky130_fd_sc_hd__a211o_1
XFILLER_0_21_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14169_ _00115_ _02124_ _04201_ _04200_ VGND VGND VPWR VPWR _04359_ sky130_fd_sc_hd__a31o_1
XTAP_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18977_ clknet_4_6_0_clk _09409_ VGND VGND VPWR VPWR salida\[30\] sky130_fd_sc_hd__dfxtp_1
XTAP_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17928_ _08405_ _08407_ VGND VGND VPWR VPWR _08448_ sky130_fd_sc_hd__and2b_1
XTAP_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17859_ _08269_ _08271_ _08372_ VGND VGND VPWR VPWR _08373_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_89_884 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_146_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_228 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_388 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_126_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_503 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_114_385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_130_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09977_ ApproximateM_inst.lob_16.lob1.genblk1\[2\].genblk1.mux.sel VGND VGND VPWR
+ VPWR _09212_ sky130_fd_sc_hd__buf_4
XFILLER_0_98_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11870_ _00515_ _01862_ VGND VGND VPWR VPWR _01963_ sky130_fd_sc_hd__nor2_2
XFILLER_0_86_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10821_ cla_inst.in2\[18\] _00179_ VGND VGND VPWR VPWR _00914_ sky130_fd_sc_hd__and2_1
X_13540_ _03649_ _03650_ _03670_ VGND VGND VPWR VPWR _03671_ sky130_fd_sc_hd__o21ai_2
X_10752_ _07711_ VGND VGND VPWR VPWR _00845_ sky130_fd_sc_hd__buf_4
XFILLER_0_95_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13471_ _03591_ _03592_ _03593_ _03594_ VGND VGND VPWR VPWR _03595_ sky130_fd_sc_hd__a211o_1
X_10683_ _00769_ _00770_ _00771_ _00775_ VGND VGND VPWR VPWR _00776_ sky130_fd_sc_hd__a211o_1
XFILLER_0_152_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15210_ _01873_ _03071_ VGND VGND VPWR VPWR _05495_ sky130_fd_sc_hd__nand2_1
X_12422_ _02448_ _02513_ _02514_ VGND VGND VPWR VPWR _02515_ sky130_fd_sc_hd__and3_1
X_16190_ _06481_ _06484_ _06506_ _06556_ VGND VGND VPWR VPWR _06557_ sky130_fd_sc_hd__a31o_1
XFILLER_0_35_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15141_ _02977_ _02980_ _03560_ VGND VGND VPWR VPWR _05420_ sky130_fd_sc_hd__or3_1
X_12353_ _02445_ VGND VGND VPWR VPWR _02446_ sky130_fd_sc_hd__inv_2
XFILLER_0_140_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11304_ _00122_ _00862_ VGND VGND VPWR VPWR _01397_ sky130_fd_sc_hd__nor2_1
XFILLER_0_120_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15072_ _05342_ _05343_ VGND VGND VPWR VPWR _05345_ sky130_fd_sc_hd__nand2_1
X_12284_ _02261_ _02262_ _02263_ _02256_ VGND VGND VPWR VPWR _02377_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_22_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14023_ cla_inst.in2\[27\] _09349_ _04657_ _04864_ VGND VGND VPWR VPWR _04200_ sky130_fd_sc_hd__and4_1
X_18900_ clknet_4_10_0_clk _00054_ VGND VGND VPWR VPWR cla_inst.in1\[18\] sky130_fd_sc_hd__dfxtp_2
X_11235_ _01315_ _01316_ _01318_ _01327_ VGND VGND VPWR VPWR _01328_ sky130_fd_sc_hd__o31a_1
XFILLER_0_121_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18831_ _09332_ VGND VGND VPWR VPWR _00101_ sky130_fd_sc_hd__clkbuf_1
X_11166_ _01241_ _01258_ VGND VGND VPWR VPWR _01259_ sky130_fd_sc_hd__xor2_1
XFILLER_0_101_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10117_ ApproximateM_inst.lob_16.lob1.genblk1\[8\].genblk1.mux.sel VGND VGND VPWR
+ VPWR _00210_ sky130_fd_sc_hd__buf_4
X_18762_ _08615_ net37 _09276_ VGND VGND VPWR VPWR _09280_ sky130_fd_sc_hd__mux2_1
X_11097_ _01123_ _01122_ VGND VGND VPWR VPWR _01190_ sky130_fd_sc_hd__and2b_1
X_15974_ _06271_ _06307_ _06321_ VGND VGND VPWR VPWR _06322_ sky130_fd_sc_hd__and3_1
X_17713_ _07978_ _08105_ _08108_ VGND VGND VPWR VPWR _08215_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_26_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14925_ _05014_ _05063_ VGND VGND VPWR VPWR _05185_ sky130_fd_sc_hd__nand2_1
X_10048_ _00118_ _00139_ _00140_ VGND VGND VPWR VPWR _00141_ sky130_fd_sc_hd__a21oi_2
X_18693_ _01692_ _09183_ _09191_ VGND VGND VPWR VPWR _09227_ sky130_fd_sc_hd__a21oi_1
Xhold90 _00009_ VGND VGND VPWR VPWR net253 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_117_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17644_ _06425_ _06442_ _08139_ VGND VGND VPWR VPWR _08140_ sky130_fd_sc_hd__or3_1
X_14856_ _05106_ _05108_ VGND VGND VPWR VPWR _05109_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_77_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13807_ net236 _03931_ _03961_ _03962_ VGND VGND VPWR VPWR _03963_ sky130_fd_sc_hd__o211ai_4
X_17575_ _08043_ _08044_ _08062_ VGND VGND VPWR VPWR _08064_ sky130_fd_sc_hd__or3b_1
X_14787_ _05016_ _04917_ _05033_ VGND VGND VPWR VPWR _05034_ sky130_fd_sc_hd__o21a_1
X_11999_ _02014_ _02091_ VGND VGND VPWR VPWR _02092_ sky130_fd_sc_hd__or2_1
XFILLER_0_42_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16526_ _03036_ _06920_ _06921_ VGND VGND VPWR VPWR _06922_ sky130_fd_sc_hd__a21o_1
X_13738_ net121 _03885_ _03887_ VGND VGND VPWR VPWR _03888_ sky130_fd_sc_hd__nor3_1
XFILLER_0_133_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16457_ _06843_ _06846_ _03080_ VGND VGND VPWR VPWR _06847_ sky130_fd_sc_hd__mux2_1
X_13669_ _03809_ net326 _03622_ _03752_ VGND VGND VPWR VPWR _03812_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_6_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15408_ _05710_ VGND VGND VPWR VPWR _05711_ sky130_fd_sc_hd__inv_2
XFILLER_0_116_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16388_ _06572_ _06664_ VGND VGND VPWR VPWR _06772_ sky130_fd_sc_hd__nor2_1
XFILLER_0_41_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18127_ _08662_ _08664_ VGND VGND VPWR VPWR _08665_ sky130_fd_sc_hd__xnor2_1
X_15339_ _09353_ _07025_ _05633_ _05634_ VGND VGND VPWR VPWR _05635_ sky130_fd_sc_hd__and4_1
XFILLER_0_13_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18058_ _08586_ _08589_ VGND VGND VPWR VPWR _08590_ sky130_fd_sc_hd__nor2_1
XFILLER_0_151_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_112_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09900_ _03793_ _04460_ _08409_ _03859_ VGND VGND VPWR VPWR _08420_ sky130_fd_sc_hd__a22oi_2
X_17009_ _07379_ _07380_ _07445_ _07446_ VGND VGND VPWR VPWR _07447_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_111_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09831_ _07515_ VGND VGND VPWR VPWR _07668_ sky130_fd_sc_hd__clkbuf_4
XTAP_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09762_ _06526_ _06537_ _04973_ _06191_ VGND VGND VPWR VPWR _06917_ sky130_fd_sc_hd__o211a_1
XTAP_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09693_ _05159_ _05170_ _04318_ _04766_ VGND VGND VPWR VPWR _06170_ sky130_fd_sc_hd__o211ai_4
Xrebuffer11 net173 VGND VGND VPWR VPWR net174 sky130_fd_sc_hd__clkbuf_1
Xrebuffer22 _00772_ VGND VGND VPWR VPWR net185 sky130_fd_sc_hd__buf_1
XTAP_2209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer33 _04741_ VGND VGND VPWR VPWR net196 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrebuffer44 net206 VGND VGND VPWR VPWR net207 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_96_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrebuffer55 _04152_ VGND VGND VPWR VPWR net218 sky130_fd_sc_hd__buf_1
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer66 net227 VGND VGND VPWR VPWR net229 sky130_fd_sc_hd__clkbuf_1
XTAP_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer77 _03376_ VGND VGND VPWR VPWR net240 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer88 _04458_ VGND VGND VPWR VPWR net335 sky130_fd_sc_hd__dlygate4sd1_1
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_504 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_147_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_367 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_130_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_114_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_664 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11020_ _00514_ VGND VGND VPWR VPWR _01113_ sky130_fd_sc_hd__clkbuf_8
X_12971_ _03028_ _00516_ VGND VGND VPWR VPWR _03064_ sky130_fd_sc_hd__nor2_1
X_14710_ _04817_ _04948_ _04949_ VGND VGND VPWR VPWR _04950_ sky130_fd_sc_hd__nand3_4
X_11922_ _02012_ _02014_ VGND VGND VPWR VPWR _02015_ sky130_fd_sc_hd__or2_1
XTAP_2710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15690_ _06015_ _06016_ VGND VGND VPWR VPWR _06017_ sky130_fd_sc_hd__and2_1
XTAP_2721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14641_ _03014_ _05921_ _04873_ _04870_ VGND VGND VPWR VPWR _04874_ sky130_fd_sc_hd__o2bb2a_1
XTAP_2754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11853_ _01848_ _01856_ VGND VGND VPWR VPWR _01946_ sky130_fd_sc_hd__xnor2_1
XTAP_2765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10804_ _00896_ VGND VGND VPWR VPWR _00897_ sky130_fd_sc_hd__inv_2
X_17360_ _07824_ _07826_ _07827_ _07828_ VGND VGND VPWR VPWR _07829_ sky130_fd_sc_hd__o22a_1
XTAP_2798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14572_ _04796_ _04797_ _04622_ VGND VGND VPWR VPWR _04800_ sky130_fd_sc_hd__o21ai_2
X_11784_ _01825_ _01824_ VGND VGND VPWR VPWR _01877_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_95_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16311_ _06685_ _06332_ _06686_ VGND VGND VPWR VPWR _06688_ sky130_fd_sc_hd__a21oi_1
X_13523_ _03005_ _00223_ VGND VGND VPWR VPWR _03653_ sky130_fd_sc_hd__nand2_1
X_10735_ _00826_ _00825_ _00818_ _00801_ VGND VGND VPWR VPWR _00828_ sky130_fd_sc_hd__o211ai_1
X_17291_ _06875_ _07318_ VGND VGND VPWR VPWR _07754_ sky130_fd_sc_hd__or2_1
XFILLER_0_137_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16242_ _07810_ _03069_ VGND VGND VPWR VPWR _06614_ sky130_fd_sc_hd__or2_1
XFILLER_0_42_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10666_ _00757_ _00758_ VGND VGND VPWR VPWR _00759_ sky130_fd_sc_hd__nor2_2
X_13454_ _03575_ _03576_ _03098_ VGND VGND VPWR VPWR _03577_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12405_ _02491_ _02496_ _02497_ VGND VGND VPWR VPWR _02498_ sky130_fd_sc_hd__or3_1
X_13385_ _03500_ _03501_ VGND VGND VPWR VPWR _03502_ sky130_fd_sc_hd__xnor2_1
X_16173_ _04449_ _04471_ _03281_ VGND VGND VPWR VPWR _06539_ sky130_fd_sc_hd__o21a_1
X_10597_ _00482_ _00487_ _00688_ _00689_ VGND VGND VPWR VPWR _00690_ sky130_fd_sc_hd__a211o_2
XFILLER_0_152_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15124_ _05398_ _05401_ VGND VGND VPWR VPWR _05402_ sky130_fd_sc_hd__xor2_2
XFILLER_0_50_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput109 net109 VGND VGND VPWR VPWR o_wb_data[4] sky130_fd_sc_hd__clkbuf_4
X_12336_ _02427_ _02428_ VGND VGND VPWR VPWR _02429_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_50_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15055_ _05324_ _05325_ VGND VGND VPWR VPWR _05326_ sky130_fd_sc_hd__nor2_1
X_12267_ _02357_ _02358_ _02359_ VGND VGND VPWR VPWR _02360_ sky130_fd_sc_hd__and3b_1
XFILLER_0_120_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11218_ _01290_ _01309_ _01308_ VGND VGND VPWR VPWR _01311_ sky130_fd_sc_hd__o21ai_2
X_14006_ _04008_ _04011_ _04009_ VGND VGND VPWR VPWR _04181_ sky130_fd_sc_hd__o21ba_1
X_12198_ _02285_ _02286_ _02268_ _02275_ VGND VGND VPWR VPWR _02291_ sky130_fd_sc_hd__o211a_1
Xoutput80 net80 VGND VGND VPWR VPWR leds[8] sky130_fd_sc_hd__buf_2
Xoutput91 net91 VGND VGND VPWR VPWR o_wb_data[17] sky130_fd_sc_hd__clkbuf_4
X_18814_ _09320_ VGND VGND VPWR VPWR _00095_ sky130_fd_sc_hd__clkbuf_1
X_11149_ _00169_ _09188_ _07591_ _00175_ VGND VGND VPWR VPWR _01242_ sky130_fd_sc_hd__a22o_1
XFILLER_0_37_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18745_ _02728_ net63 _09251_ VGND VGND VPWR VPWR _09266_ sky130_fd_sc_hd__mux2_1
X_15957_ _06274_ _06302_ _06303_ VGND VGND VPWR VPWR _06304_ sky130_fd_sc_hd__o21ba_1
X_14908_ _01504_ _01317_ VGND VGND VPWR VPWR _05166_ sky130_fd_sc_hd__nand2_1
X_18676_ net38 _09189_ _09215_ VGND VGND VPWR VPWR _00048_ sky130_fd_sc_hd__o21a_1
X_15888_ _06227_ _06228_ _06230_ VGND VGND VPWR VPWR _09373_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_144_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17627_ _08119_ _08120_ VGND VGND VPWR VPWR _08121_ sky130_fd_sc_hd__or2_1
X_14839_ _03538_ _04241_ _03918_ VGND VGND VPWR VPWR _05091_ sky130_fd_sc_hd__and3_1
X_17558_ _06755_ _07741_ VGND VGND VPWR VPWR _08045_ sky130_fd_sc_hd__or2_1
XFILLER_0_74_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16509_ _06902_ VGND VGND VPWR VPWR _06903_ sky130_fd_sc_hd__inv_2
X_17489_ _07968_ _07969_ VGND VGND VPWR VPWR _07970_ sky130_fd_sc_hd__nand2_1
XFILLER_0_144_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_116_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09814_ _07210_ _07319_ _07472_ VGND VGND VPWR VPWR _07482_ sky130_fd_sc_hd__a21o_2
X_09745_ _06722_ VGND VGND VPWR VPWR _06732_ sky130_fd_sc_hd__buf_4
XTAP_2006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09676_ _05975_ VGND VGND VPWR VPWR _05986_ sky130_fd_sc_hd__buf_4
XTAP_2017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_684 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_119_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10520_ _03892_ _05333_ _05039_ _03881_ VGND VGND VPWR VPWR _00613_ sky130_fd_sc_hd__a22o_1
XFILLER_0_64_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10451_ _00388_ _00389_ VGND VGND VPWR VPWR _00544_ sky130_fd_sc_hd__or2_1
XFILLER_0_91_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13170_ _03005_ _01248_ VGND VGND VPWR VPWR _03269_ sky130_fd_sc_hd__nand2_1
X_10382_ _08724_ _00309_ _00312_ _00311_ VGND VGND VPWR VPWR _00475_ sky130_fd_sc_hd__a31o_1
XFILLER_0_20_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12121_ _03607_ VGND VGND VPWR VPWR _02214_ sky130_fd_sc_hd__inv_2
XFILLER_0_102_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12052_ _02104_ _02103_ VGND VGND VPWR VPWR _02145_ sky130_fd_sc_hd__xnor2_1
X_11003_ _07352_ _00459_ _01094_ _01095_ VGND VGND VPWR VPWR _01096_ sky130_fd_sc_hd__nand4_2
X_16860_ _07245_ _07246_ VGND VGND VPWR VPWR _07284_ sky130_fd_sc_hd__nand2_1
X_15811_ _02974_ _06144_ _06147_ VGND VGND VPWR VPWR _06148_ sky130_fd_sc_hd__a21o_1
X_16791_ _07206_ _07208_ VGND VGND VPWR VPWR _07209_ sky130_fd_sc_hd__nand2_1
X_18530_ net26 net25 net23 VGND VGND VPWR VPWR _09099_ sky130_fd_sc_hd__or3b_2
X_15742_ _06071_ _06072_ VGND VGND VPWR VPWR _06074_ sky130_fd_sc_hd__and2_1
X_12954_ _01106_ VGND VGND VPWR VPWR _03047_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_59_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18461_ _06328_ _06411_ _06410_ _06024_ VGND VGND VPWR VPWR _09026_ sky130_fd_sc_hd__a211o_1
X_11905_ _01810_ _01903_ VGND VGND VPWR VPWR _01998_ sky130_fd_sc_hd__xnor2_4
X_15673_ _05991_ _05996_ VGND VGND VPWR VPWR _05999_ sky130_fd_sc_hd__nand2_1
XTAP_2540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12885_ _02977_ VGND VGND VPWR VPWR _02978_ sky130_fd_sc_hd__clkbuf_4
XTAP_2562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17412_ _07742_ _07747_ _07884_ VGND VGND VPWR VPWR _07887_ sky130_fd_sc_hd__and3_1
X_14624_ _02188_ _00502_ VGND VGND VPWR VPWR _04856_ sky130_fd_sc_hd__nand2_1
XTAP_2573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_504 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11836_ net182 VGND VGND VPWR VPWR _01929_ sky130_fd_sc_hd__inv_2
X_18392_ _03107_ _07596_ VGND VGND VPWR VPWR _08952_ sky130_fd_sc_hd__nand2_1
XTAP_2584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17343_ _06371_ _06545_ _07811_ _03311_ VGND VGND VPWR VPWR _07812_ sky130_fd_sc_hd__a22o_1
X_14555_ _04614_ _04616_ VGND VGND VPWR VPWR _04781_ sky130_fd_sc_hd__nor2_1
XTAP_1883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11767_ net175 net180 VGND VGND VPWR VPWR _01860_ sky130_fd_sc_hd__nand2_1
XTAP_1894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13506_ _05213_ cla_inst.in1\[28\] VGND VGND VPWR VPWR _03634_ sky130_fd_sc_hd__and2_2
X_10718_ _00805_ _00809_ VGND VGND VPWR VPWR _00811_ sky130_fd_sc_hd__xor2_1
X_17274_ _07637_ _07638_ VGND VGND VPWR VPWR _07736_ sky130_fd_sc_hd__and2_1
X_14486_ _02984_ _01520_ _07112_ _00308_ VGND VGND VPWR VPWR _04705_ sky130_fd_sc_hd__and4_1
XFILLER_0_153_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11698_ _01221_ _01693_ _01774_ VGND VGND VPWR VPWR _01791_ sky130_fd_sc_hd__nor3_1
XFILLER_0_70_326 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19013_ clknet_4_3_0_clk _00103_ VGND VGND VPWR VPWR op_code\[2\] sky130_fd_sc_hd__dfxtp_4
X_16225_ _03161_ _06593_ _06594_ VGND VGND VPWR VPWR _06595_ sky130_fd_sc_hd__a21o_1
X_13437_ _02976_ _03038_ _03534_ _03558_ _03121_ VGND VGND VPWR VPWR _03559_ sky130_fd_sc_hd__o32a_1
XFILLER_0_130_47 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10649_ _00739_ _00740_ _00529_ _00699_ VGND VGND VPWR VPWR _00742_ sky130_fd_sc_hd__a211oi_2
Xrebuffer2 _00662_ VGND VGND VPWR VPWR net165 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16156_ sel_op\[3\] _03281_ sel_op\[2\] VGND VGND VPWR VPWR _06520_ sky130_fd_sc_hd__o21bai_4
XFILLER_0_51_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13368_ _03480_ _03481_ VGND VGND VPWR VPWR _03483_ sky130_fd_sc_hd__nand2_1
X_15107_ _05381_ _05382_ VGND VGND VPWR VPWR _05383_ sky130_fd_sc_hd__and2_1
X_12319_ _02410_ _02405_ _02409_ VGND VGND VPWR VPWR _02412_ sky130_fd_sc_hd__and3_1
X_16087_ _03044_ _06444_ VGND VGND VPWR VPWR _06445_ sky130_fd_sc_hd__and2_1
X_13299_ _03393_ _03394_ _03405_ VGND VGND VPWR VPWR _03407_ sky130_fd_sc_hd__or3_2
X_15038_ _04246_ _04249_ _04247_ VGND VGND VPWR VPWR _05308_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16989_ _07409_ _07424_ VGND VGND VPWR VPWR _07425_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_79_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09530_ ApproximateM_inst.lob_16.lob1.genblk1\[14\].genblk1.mux.sel VGND VGND VPWR
+ VPWR _04395_ sky130_fd_sc_hd__buf_6
XFILLER_0_64_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18728_ _09245_ _09252_ VGND VGND VPWR VPWR _09253_ sky130_fd_sc_hd__and2_1
X_09461_ _03596_ _03476_ _03618_ _03629_ VGND VGND VPWR VPWR _03640_ sky130_fd_sc_hd__a22o_1
XFILLER_0_64_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18659_ _09202_ VGND VGND VPWR VPWR _00042_ sky130_fd_sc_hd__buf_1
XFILLER_0_94_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_526 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_136_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_304 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_140_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09728_ _04973_ _06191_ _06526_ _06537_ VGND VGND VPWR VPWR _06548_ sky130_fd_sc_hd__a211oi_2
X_09659_ _05551_ _05791_ VGND VGND VPWR VPWR _05802_ sky130_fd_sc_hd__xnor2_2
XTAP_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12670_ _02733_ _02738_ _02737_ VGND VGND VPWR VPWR _02763_ sky130_fd_sc_hd__a21o_1
XTAP_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11621_ _01192_ _01712_ _01711_ VGND VGND VPWR VPWR _01714_ sky130_fd_sc_hd__a21o_1
XFILLER_0_148_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14340_ _04350_ _04422_ _04544_ _04545_ VGND VGND VPWR VPWR _04546_ sky130_fd_sc_hd__a211oi_2
X_11552_ _06971_ _04580_ _01643_ _01644_ VGND VGND VPWR VPWR _01645_ sky130_fd_sc_hd__nand4_2
XFILLER_0_107_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10503_ _00589_ _00595_ VGND VGND VPWR VPWR _00596_ sky130_fd_sc_hd__or2_2
X_14271_ _04299_ net127 _04468_ _04469_ VGND VGND VPWR VPWR _04470_ sky130_fd_sc_hd__o211ai_4
X_11483_ _05736_ _01575_ VGND VGND VPWR VPWR _01576_ sky130_fd_sc_hd__nand2_1
XFILLER_0_61_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16010_ _00644_ _00248_ VGND VGND VPWR VPWR _06360_ sky130_fd_sc_hd__or2_1
X_10434_ _00507_ _00508_ _00526_ VGND VGND VPWR VPWR _00527_ sky130_fd_sc_hd__o21a_1
X_13222_ _00148_ _09350_ _00212_ _00206_ VGND VGND VPWR VPWR _03325_ sky130_fd_sc_hd__and4_1
XFILLER_0_150_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_735 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10365_ _00456_ _00457_ VGND VGND VPWR VPWR _00458_ sky130_fd_sc_hd__and2b_1
X_13153_ _05453_ _00645_ _07156_ _06732_ VGND VGND VPWR VPWR _03251_ sky130_fd_sc_hd__nand4_4
XTAP_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12104_ _02195_ _02196_ VGND VGND VPWR VPWR _02197_ sky130_fd_sc_hd__nand2_1
X_13084_ _02563_ _03175_ _03022_ VGND VGND VPWR VPWR _03176_ sky130_fd_sc_hd__o21ai_1
X_17961_ _08482_ _08483_ VGND VGND VPWR VPWR _08484_ sky130_fd_sc_hd__nand2_1
XTAP_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10296_ _00387_ _00388_ cla_inst.in2\[25\] _00172_ VGND VGND VPWR VPWR _00389_ sky130_fd_sc_hd__and4bb_1
X_12035_ _01106_ _00515_ _02045_ _02127_ VGND VGND VPWR VPWR _02128_ sky130_fd_sc_hd__or4_4
X_16912_ _07339_ _07340_ VGND VGND VPWR VPWR _07342_ sky130_fd_sc_hd__xnor2_1
X_17892_ _08314_ _08347_ _08408_ VGND VGND VPWR VPWR _08410_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_18_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16843_ _02979_ _06642_ VGND VGND VPWR VPWR _07267_ sky130_fd_sc_hd__nor2_1
XFILLER_0_88_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16774_ _07149_ _07151_ VGND VGND VPWR VPWR _07191_ sky130_fd_sc_hd__and2_1
X_13986_ _04155_ _04157_ _04151_ VGND VGND VPWR VPWR _04159_ sky130_fd_sc_hd__o21ai_1
X_18513_ _06248_ _06414_ _09076_ VGND VGND VPWR VPWR _09082_ sky130_fd_sc_hd__o21bai_1
X_15725_ _05917_ _06054_ VGND VGND VPWR VPWR _06055_ sky130_fd_sc_hd__and2_1
XFILLER_0_88_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12937_ _03028_ _03029_ VGND VGND VPWR VPWR _03030_ sky130_fd_sc_hd__nand2_1
XFILLER_0_34_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18444_ _08912_ _08965_ VGND VGND VPWR VPWR _09008_ sky130_fd_sc_hd__nor2_1
X_15656_ _05973_ _05978_ _05979_ VGND VGND VPWR VPWR _05980_ sky130_fd_sc_hd__and3_1
XFILLER_0_75_418 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12868_ _02949_ _02955_ _02954_ VGND VGND VPWR VPWR _02961_ sky130_fd_sc_hd__a21bo_1
XTAP_2381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14607_ _03377_ cla_inst.in1\[27\] _07102_ _03356_ VGND VGND VPWR VPWR _04837_ sky130_fd_sc_hd__a22o_1
X_18375_ _08932_ _08933_ VGND VGND VPWR VPWR _08934_ sky130_fd_sc_hd__xnor2_4
X_11819_ _06460_ _00147_ _01911_ _01909_ VGND VGND VPWR VPWR _01912_ sky130_fd_sc_hd__a31o_1
X_15587_ _05815_ _05817_ _05903_ _05904_ VGND VGND VPWR VPWR _05905_ sky130_fd_sc_hd__a211oi_2
XTAP_1680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12799_ _02884_ _02886_ VGND VGND VPWR VPWR _02892_ sky130_fd_sc_hd__or2_2
X_17326_ _07669_ VGND VGND VPWR VPWR _07793_ sky130_fd_sc_hd__inv_2
X_14538_ _04760_ _04761_ VGND VGND VPWR VPWR _04762_ sky130_fd_sc_hd__nor2_1
XFILLER_0_141_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17257_ _07710_ _07716_ VGND VGND VPWR VPWR _07717_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_153_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14469_ net177 _04684_ _04685_ VGND VGND VPWR VPWR _04687_ sky130_fd_sc_hd__o21ai_1
X_16208_ _03281_ _06575_ _06520_ VGND VGND VPWR VPWR _06576_ sky130_fd_sc_hd__a21o_1
XFILLER_0_113_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17188_ _07620_ _07641_ VGND VGND VPWR VPWR _07642_ sky130_fd_sc_hd__xor2_1
XFILLER_0_59_20 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_595 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16139_ _06499_ _06500_ _03152_ VGND VGND VPWR VPWR _06501_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_122_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09513_ _03684_ _03640_ _03585_ VGND VGND VPWR VPWR _04209_ sky130_fd_sc_hd__a21o_1
XFILLER_0_149_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09444_ cla_inst.in2\[18\] VGND VGND VPWR VPWR _03454_ sky130_fd_sc_hd__buf_6
XPHY_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_531 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_679 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_104_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_882 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10150_ _00234_ _00242_ VGND VGND VPWR VPWR _00243_ sky130_fd_sc_hd__xnor2_1
X_10081_ cla_inst.in2\[23\] VGND VGND VPWR VPWR _00174_ sky130_fd_sc_hd__buf_2
X_13840_ _03997_ _03998_ VGND VGND VPWR VPWR _03999_ sky130_fd_sc_hd__nor2_1
X_13771_ _03085_ _03088_ _03050_ VGND VGND VPWR VPWR _03924_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10983_ _01051_ _01052_ _01039_ _01050_ VGND VGND VPWR VPWR _01076_ sky130_fd_sc_hd__a211o_1
XFILLER_0_97_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15510_ _05819_ _05820_ VGND VGND VPWR VPWR _05821_ sky130_fd_sc_hd__nor2_1
XFILLER_0_85_716 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12722_ _02759_ _02790_ VGND VGND VPWR VPWR _02815_ sky130_fd_sc_hd__and2_1
XFILLER_0_139_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16490_ _06877_ _06881_ VGND VGND VPWR VPWR _06882_ sky130_fd_sc_hd__xor2_1
XFILLER_0_78_790 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15441_ _05654_ _05657_ _05655_ VGND VGND VPWR VPWR _05746_ sky130_fd_sc_hd__o21ba_1
X_12653_ _02710_ _02745_ VGND VGND VPWR VPWR _02746_ sky130_fd_sc_hd__or2_1
X_11604_ _00845_ _01695_ _01696_ VGND VGND VPWR VPWR _01697_ sky130_fd_sc_hd__a21oi_2
X_18160_ _06366_ _07592_ _07650_ _07596_ VGND VGND VPWR VPWR _08700_ sky130_fd_sc_hd__a22o_1
X_15372_ _05651_ _05670_ VGND VGND VPWR VPWR _05672_ sky130_fd_sc_hd__nor2_1
XFILLER_0_53_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12584_ ApproximateM_inst.lob_16.lob2.genblk1\[2\].genblk1.mux.sel _01031_ VGND VGND
+ VPWR VPWR _02677_ sky130_fd_sc_hd__and2_2
XFILLER_0_26_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_154_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17111_ _07345_ _07349_ _07447_ _07448_ _07556_ VGND VGND VPWR VPWR _07558_ sky130_fd_sc_hd__o311a_4
XFILLER_0_142_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14323_ _04525_ _04527_ VGND VGND VPWR VPWR _04528_ sky130_fd_sc_hd__nand2_1
X_11535_ _01212_ _01211_ VGND VGND VPWR VPWR _01628_ sky130_fd_sc_hd__and2b_1
X_18091_ _07318_ _07706_ VGND VGND VPWR VPWR _08625_ sky130_fd_sc_hd__nor2_2
XFILLER_0_151_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17042_ _07285_ _07295_ _07405_ VGND VGND VPWR VPWR _07483_ sky130_fd_sc_hd__and3_1
X_14254_ _04450_ _04451_ _04558_ _00502_ VGND VGND VPWR VPWR _04452_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_151_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11466_ _01557_ _01558_ VGND VGND VPWR VPWR _01559_ sky130_fd_sc_hd__xor2_1
XFILLER_0_34_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13205_ _01745_ _00716_ _03304_ VGND VGND VPWR VPWR _03306_ sky130_fd_sc_hd__a21o_1
XFILLER_0_111_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10417_ _07788_ _00509_ _07570_ cla_inst.in2\[31\] VGND VGND VPWR VPWR _00510_ sky130_fd_sc_hd__a22oi_1
X_14185_ _04355_ _04356_ _04375_ VGND VGND VPWR VPWR _04377_ sky130_fd_sc_hd__nand3_1
X_11397_ _01468_ _01488_ _01489_ VGND VGND VPWR VPWR _01490_ sky130_fd_sc_hd__nand3_2
XFILLER_0_110_228 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13136_ _03227_ _03231_ _03232_ VGND VGND VPWR VPWR _03233_ sky130_fd_sc_hd__and3_1
XTAP_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10348_ _03892_ _05028_ _00439_ _03881_ VGND VGND VPWR VPWR _00441_ sky130_fd_sc_hd__a22o_1
XTAP_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18993_ clknet_4_6_0_clk _09359_ VGND VGND VPWR VPWR salida\[46\] sky130_fd_sc_hd__dfxtp_1
XTAP_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10279_ _00370_ _00371_ _09152_ _09338_ VGND VGND VPWR VPWR _00372_ sky130_fd_sc_hd__a211o_1
XTAP_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13067_ _03090_ _03151_ _03158_ VGND VGND VPWR VPWR _03159_ sky130_fd_sc_hd__o21ai_2
X_17944_ _08464_ _08465_ VGND VGND VPWR VPWR _08466_ sky130_fd_sc_hd__and2_1
X_12018_ _07363_ _04045_ _02109_ _02110_ VGND VGND VPWR VPWR _02111_ sky130_fd_sc_hd__a31o_1
X_17875_ _08389_ _08390_ VGND VGND VPWR VPWR _08391_ sky130_fd_sc_hd__nand2_1
XFILLER_0_45_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16826_ _07191_ _07192_ _07247_ VGND VGND VPWR VPWR _07248_ sky130_fd_sc_hd__nor3_1
X_16757_ _07172_ _06354_ _06355_ VGND VGND VPWR VPWR _07173_ sky130_fd_sc_hd__nand3_1
X_13969_ _04128_ _04129_ _04138_ VGND VGND VPWR VPWR _04140_ sky130_fd_sc_hd__and3_1
XFILLER_0_76_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15708_ _03015_ _03067_ _05960_ _05959_ VGND VGND VPWR VPWR _06036_ sky130_fd_sc_hd__a31o_1
X_16688_ _07096_ _07097_ _06836_ VGND VGND VPWR VPWR _07098_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15639_ _05959_ _03067_ _03015_ _05960_ VGND VGND VPWR VPWR _05961_ sky130_fd_sc_hd__and4b_1
X_18427_ _06408_ _06449_ _08989_ VGND VGND VPWR VPWR _08990_ sky130_fd_sc_hd__o21ai_1
X_18358_ _08862_ _08894_ _08914_ VGND VGND VPWR VPWR _08915_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_84_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_22 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17309_ _07773_ VGND VGND VPWR VPWR _07774_ sky130_fd_sc_hd__inv_2
XFILLER_0_127_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18289_ _08736_ _08739_ _08809_ VGND VGND VPWR VPWR _08840_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_43_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_852 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09993_ _09240_ _09326_ VGND VGND VPWR VPWR _09333_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_50_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09427_ sel_op\[3\] _03206_ _03260_ _03239_ VGND VGND VPWR VPWR _00003_ sky130_fd_sc_hd__a22o_1
XFILLER_0_137_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_771 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_443 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_117_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_117_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11320_ _01394_ _01395_ _01412_ VGND VGND VPWR VPWR _01413_ sky130_fd_sc_hd__nor3b_4
XFILLER_0_105_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11251_ _00169_ _00130_ _01342_ _01343_ VGND VGND VPWR VPWR _01344_ sky130_fd_sc_hd__and4_1
XFILLER_0_120_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10202_ _04504_ _00294_ _08049_ _05377_ VGND VGND VPWR VPWR _00295_ sky130_fd_sc_hd__and4_1
X_11182_ _00964_ _00963_ VGND VGND VPWR VPWR _01275_ sky130_fd_sc_hd__or2b_1
XFILLER_0_101_762 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10133_ _00215_ _00225_ VGND VGND VPWR VPWR _00226_ sky130_fd_sc_hd__xnor2_1
X_15990_ _06335_ _06336_ _06337_ VGND VGND VPWR VPWR _06338_ sky130_fd_sc_hd__a21bo_1
X_10064_ _08202_ _00143_ _00156_ VGND VGND VPWR VPWR _00157_ sky130_fd_sc_hd__o21a_1
X_14941_ _04951_ _05200_ _05201_ VGND VGND VPWR VPWR _05202_ sky130_fd_sc_hd__a21boi_1
X_17660_ _08045_ _08046_ VGND VGND VPWR VPWR _08156_ sky130_fd_sc_hd__nand2_1
X_14872_ _00678_ _06471_ _08452_ _00679_ VGND VGND VPWR VPWR _05127_ sky130_fd_sc_hd__a22o_1
X_16611_ _02828_ _07012_ _03930_ _07013_ VGND VGND VPWR VPWR _07014_ sky130_fd_sc_hd__o211a_1
X_13823_ _03963_ _03964_ _03980_ VGND VGND VPWR VPWR _03981_ sky130_fd_sc_hd__a21o_1
X_17591_ _07954_ _07964_ _08080_ VGND VGND VPWR VPWR _08081_ sky130_fd_sc_hd__a21o_1
X_16542_ _06653_ _06937_ _06886_ VGND VGND VPWR VPWR _06939_ sky130_fd_sc_hd__nor3_1
X_13754_ _03043_ _03046_ _03090_ VGND VGND VPWR VPWR _03906_ sky130_fd_sc_hd__mux2_1
X_10966_ _00987_ _00986_ VGND VGND VPWR VPWR _01059_ sky130_fd_sc_hd__and2b_1
XFILLER_0_57_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12705_ _02795_ _02797_ VGND VGND VPWR VPWR _02798_ sky130_fd_sc_hd__and2b_1
X_16473_ _06833_ _06835_ _06864_ VGND VGND VPWR VPWR _06865_ sky130_fd_sc_hd__o21a_1
X_13685_ _03828_ _03829_ VGND VGND VPWR VPWR _03830_ sky130_fd_sc_hd__nand2_1
X_10897_ _00985_ _00988_ VGND VGND VPWR VPWR _00990_ sky130_fd_sc_hd__xor2_1
X_18212_ _04900_ _06446_ VGND VGND VPWR VPWR _08758_ sky130_fd_sc_hd__nor2_1
X_15424_ _05720_ _05727_ VGND VGND VPWR VPWR _05728_ sky130_fd_sc_hd__and2_1
XFILLER_0_66_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12636_ _08865_ _01746_ _01357_ _02728_ VGND VGND VPWR VPWR _02729_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_65_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18143_ _08682_ _06396_ _06397_ VGND VGND VPWR VPWR _08683_ sky130_fd_sc_hd__and3_1
X_15355_ _05582_ _05581_ VGND VGND VPWR VPWR _05653_ sky130_fd_sc_hd__or2b_1
XFILLER_0_142_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12567_ _02613_ _02653_ _02643_ _02652_ VGND VGND VPWR VPWR _02660_ sky130_fd_sc_hd__a211o_1
XFILLER_0_109_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14306_ _04507_ _04508_ VGND VGND VPWR VPWR _04509_ sky130_fd_sc_hd__nor2_2
XFILLER_0_81_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11518_ _01552_ _01554_ _01553_ VGND VGND VPWR VPWR _01611_ sky130_fd_sc_hd__a21bo_1
X_18074_ _04647_ _08428_ _02998_ VGND VGND VPWR VPWR _08608_ sky130_fd_sc_hd__or3b_1
XFILLER_0_25_189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15286_ _02993_ _02996_ _09059_ _00322_ VGND VGND VPWR VPWR _05578_ sky130_fd_sc_hd__and4_1
XFILLER_0_40_115 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12498_ _02580_ _02581_ _02574_ VGND VGND VPWR VPWR _02591_ sky130_fd_sc_hd__o21a_1
XFILLER_0_151_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_151_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17025_ _07462_ _07463_ _07464_ VGND VGND VPWR VPWR _07465_ sky130_fd_sc_hd__a21o_1
X_14237_ _02986_ _00309_ _04430_ _04431_ VGND VGND VPWR VPWR _04433_ sky130_fd_sc_hd__a22oi_4
X_11449_ _04427_ _03607_ _00217_ _04504_ VGND VGND VPWR VPWR _01542_ sky130_fd_sc_hd__a22o_1
X_14168_ _04196_ _04204_ VGND VGND VPWR VPWR _04358_ sky130_fd_sc_hd__and2_1
XTAP_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13119_ _03210_ _03211_ _03212_ VGND VGND VPWR VPWR _03214_ sky130_fd_sc_hd__a21o_1
XTAP_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14099_ _04276_ _04281_ VGND VGND VPWR VPWR _04282_ sky130_fd_sc_hd__xnor2_1
X_18976_ clknet_4_7_0_clk _09407_ VGND VGND VPWR VPWR salida\[29\] sky130_fd_sc_hd__dfxtp_1
XTAP_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17927_ _08320_ _08412_ VGND VGND VPWR VPWR _08447_ sky130_fd_sc_hd__nor2_1
XTAP_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17858_ _08370_ _08371_ VGND VGND VPWR VPWR _08372_ sky130_fd_sc_hd__xor2_1
XFILLER_0_22_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16809_ _07193_ _07228_ VGND VGND VPWR VPWR _07229_ sky130_fd_sc_hd__or2_1
X_17789_ _08179_ _08172_ VGND VGND VPWR VPWR _08297_ sky130_fd_sc_hd__and2b_1
XFILLER_0_88_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_127_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_114_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09976_ _09172_ _07559_ _07602_ _09166_ VGND VGND VPWR VPWR _09205_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_99_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10820_ _03454_ _00909_ _00910_ _00911_ VGND VGND VPWR VPWR _00913_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10751_ _00836_ _00841_ _00843_ VGND VGND VPWR VPWR _00844_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_94_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13470_ _03574_ _05039_ _03376_ _03378_ VGND VGND VPWR VPWR _03594_ sky130_fd_sc_hd__and4_1
XFILLER_0_94_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10682_ _00771_ _00773_ _03454_ _00774_ VGND VGND VPWR VPWR _00775_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_137_467 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12421_ _02446_ _02447_ _02417_ VGND VGND VPWR VPWR _02514_ sky130_fd_sc_hd__a21o_1
XFILLER_0_124_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15140_ _04259_ _04262_ _03081_ VGND VGND VPWR VPWR _05419_ sky130_fd_sc_hd__mux2_1
X_12352_ _02433_ _02441_ _02443_ _02444_ VGND VGND VPWR VPWR _02445_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_133_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11303_ _00863_ VGND VGND VPWR VPWR _01396_ sky130_fd_sc_hd__inv_2
X_15071_ _05330_ _05341_ VGND VGND VPWR VPWR _05343_ sky130_fd_sc_hd__or2_1
X_12283_ _02369_ _02372_ _02374_ _02375_ VGND VGND VPWR VPWR _02376_ sky130_fd_sc_hd__or4_4
X_14022_ _00125_ _03750_ _04864_ _00151_ VGND VGND VPWR VPWR _04199_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_31_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11234_ _01324_ _01326_ VGND VGND VPWR VPWR _01327_ sky130_fd_sc_hd__xor2_1
XFILLER_0_120_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18830_ net35 _03239_ _09331_ VGND VGND VPWR VPWR _09332_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11165_ _01254_ _01257_ VGND VGND VPWR VPWR _01258_ sky130_fd_sc_hd__xnor2_1
X_10116_ _00204_ _00207_ _00208_ VGND VGND VPWR VPWR _00209_ sky130_fd_sc_hd__and3_1
X_11096_ _06711_ _04591_ VGND VGND VPWR VPWR _01189_ sky130_fd_sc_hd__nand2_2
X_18761_ _09278_ VGND VGND VPWR VPWR _00078_ sky130_fd_sc_hd__clkbuf_1
X_15973_ _06282_ _06308_ VGND VGND VPWR VPWR _06321_ sky130_fd_sc_hd__nand2_1
X_17712_ _08211_ _08212_ VGND VGND VPWR VPWR _08214_ sky130_fd_sc_hd__xnor2_1
X_14924_ _05139_ _05183_ VGND VGND VPWR VPWR _05184_ sky130_fd_sc_hd__xnor2_1
X_10047_ _00123_ _00138_ VGND VGND VPWR VPWR _00140_ sky130_fd_sc_hd__and2_1
XFILLER_0_117_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18692_ _09225_ VGND VGND VPWR VPWR _00055_ sky130_fd_sc_hd__buf_1
XFILLER_0_89_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold91 ApproximateM_inst.lob_16.lob1.genblk1\[1\].genblk1.mux.sel VGND VGND VPWR
+ VPWR net254 sky130_fd_sc_hd__buf_1
XFILLER_0_26_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14855_ _05107_ _04972_ VGND VGND VPWR VPWR _05108_ sky130_fd_sc_hd__nor2_2
X_17643_ _03693_ _06441_ _03111_ VGND VGND VPWR VPWR _08139_ sky130_fd_sc_hd__a21oi_1
X_13806_ _03949_ _03950_ _03960_ VGND VGND VPWR VPWR _03962_ sky130_fd_sc_hd__or3_4
XFILLER_0_86_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17574_ _08043_ _08044_ _08062_ VGND VGND VPWR VPWR _08063_ sky130_fd_sc_hd__o21ba_1
X_14786_ _05030_ _05032_ VGND VGND VPWR VPWR _05033_ sky130_fd_sc_hd__xnor2_1
X_11998_ _05213_ _00171_ _02012_ _02013_ VGND VGND VPWR VPWR _02091_ sky130_fd_sc_hd__o2bb2a_1
X_16525_ _06550_ VGND VGND VPWR VPWR _06921_ sky130_fd_sc_hd__clkbuf_4
X_13737_ _03886_ _03722_ VGND VGND VPWR VPWR _03887_ sky130_fd_sc_hd__nor2_1
X_10949_ _00951_ _00950_ VGND VGND VPWR VPWR _01042_ sky130_fd_sc_hd__and2b_1
XFILLER_0_86_888 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16456_ _06845_ VGND VGND VPWR VPWR _06846_ sky130_fd_sc_hd__inv_2
X_13668_ _03622_ _03752_ _03809_ net189 VGND VGND VPWR VPWR _03811_ sky130_fd_sc_hd__a211o_1
XFILLER_0_6_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15407_ _05708_ _05709_ VGND VGND VPWR VPWR _05710_ sky130_fd_sc_hd__or2b_1
X_12619_ _02691_ _02711_ VGND VGND VPWR VPWR _02712_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16387_ _06769_ _06770_ VGND VGND VPWR VPWR _06771_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13599_ _03733_ _03735_ VGND VGND VPWR VPWR _03736_ sky130_fd_sc_hd__xor2_1
X_18126_ _08663_ _08570_ _08568_ VGND VGND VPWR VPWR _08664_ sky130_fd_sc_hd__o21ai_1
X_15338_ _02991_ _09351_ _07123_ _00318_ VGND VGND VPWR VPWR _05634_ sky130_fd_sc_hd__nand4_2
XFILLER_0_41_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18057_ _08418_ _08587_ _08588_ VGND VGND VPWR VPWR _08589_ sky130_fd_sc_hd__o21a_1
X_15269_ _09351_ _00318_ _05758_ _03322_ VGND VGND VPWR VPWR _05559_ sky130_fd_sc_hd__a22o_1
XFILLER_0_111_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17008_ _07443_ _07444_ _07381_ _07336_ VGND VGND VPWR VPWR _07446_ sky130_fd_sc_hd__o211a_1
XTAP_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09830_ _07613_ VGND VGND VPWR VPWR _07657_ sky130_fd_sc_hd__buf_4
XTAP_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09761_ _06895_ VGND VGND VPWR VPWR _06906_ sky130_fd_sc_hd__buf_2
XTAP_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18959_ clknet_4_6_0_clk _09389_ VGND VGND VPWR VPWR salida\[12\] sky130_fd_sc_hd__dfxtp_1
XTAP_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09692_ _05943_ _06138_ _05812_ _05823_ VGND VGND VPWR VPWR _06159_ sky130_fd_sc_hd__a211o_1
Xrebuffer12 _01845_ VGND VGND VPWR VPWR net175 sky130_fd_sc_hd__clkbuf_1
Xrebuffer23 _00336_ VGND VGND VPWR VPWR net186 sky130_fd_sc_hd__buf_1
Xrebuffer34 _06076_ VGND VGND VPWR VPWR net197 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrebuffer45 ApproximateM_inst.lob_16.lob1.genblk1\[11\].genblk1.mux.sel VGND VGND
+ VPWR VPWR net208 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrebuffer56 net218 VGND VGND VPWR VPWR net219 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer67 _05311_ VGND VGND VPWR VPWR net230 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer78 _03376_ VGND VGND VPWR VPWR net241 sky130_fd_sc_hd__clkbuf_1
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer89 _03759_ VGND VGND VPWR VPWR net336 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_0_138_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_119_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_476 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_777 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_142_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_676 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_130_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09959_ _08224_ VGND VGND VPWR VPWR _09059_ sky130_fd_sc_hd__buf_4
X_12970_ _03051_ _03059_ _03062_ VGND VGND VPWR VPWR _03063_ sky130_fd_sc_hd__mux2_1
X_11921_ _02012_ _02013_ ApproximateM_inst.lob_16.lob2.genblk1\[8\].genblk1.mux.sel
+ _00217_ VGND VGND VPWR VPWR _02014_ sky130_fd_sc_hd__and4bb_1
XTAP_2700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14640_ _04871_ VGND VGND VPWR VPWR _04873_ sky130_fd_sc_hd__inv_2
XTAP_2744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11852_ _01944_ VGND VGND VPWR VPWR _01945_ sky130_fd_sc_hd__inv_2
XTAP_2755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10803_ _00273_ _00892_ _00856_ _00891_ VGND VGND VPWR VPWR _00896_ sky130_fd_sc_hd__a211oi_2
XTAP_2788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14571_ _04622_ _04796_ _04797_ VGND VGND VPWR VPWR _04798_ sky130_fd_sc_hd__or3_2
XTAP_2799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11783_ _01872_ _01875_ VGND VGND VPWR VPWR _01876_ sky130_fd_sc_hd__and2_1
XFILLER_0_55_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16310_ _06685_ _06332_ _06686_ VGND VGND VPWR VPWR _06687_ sky130_fd_sc_hd__and3_1
X_13522_ _03449_ _03462_ _03460_ VGND VGND VPWR VPWR _03652_ sky130_fd_sc_hd__a21o_1
X_10734_ _00801_ _00818_ _00825_ _00826_ VGND VGND VPWR VPWR _00827_ sky130_fd_sc_hd__a211o_1
XFILLER_0_55_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17290_ _07750_ _07752_ VGND VGND VPWR VPWR _07753_ sky130_fd_sc_hd__nand2_1
XFILLER_0_94_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16241_ _03027_ _03056_ _00121_ VGND VGND VPWR VPWR _06612_ sky130_fd_sc_hd__a21o_1
X_13453_ _03176_ _03182_ _03048_ VGND VGND VPWR VPWR _03576_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10665_ _00756_ _00590_ _00597_ VGND VGND VPWR VPWR _00758_ sky130_fd_sc_hd__and3_1
X_12404_ _02421_ _02490_ _02488_ VGND VGND VPWR VPWR _02497_ sky130_fd_sc_hd__o21a_1
X_16172_ _03739_ _03804_ VGND VGND VPWR VPWR _06538_ sky130_fd_sc_hd__or2_1
X_13384_ _00107_ _00247_ VGND VGND VPWR VPWR _03501_ sky130_fd_sc_hd__nand2_1
XFILLER_0_63_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10596_ _00676_ _00677_ _00687_ VGND VGND VPWR VPWR _00689_ sky130_fd_sc_hd__nor3b_2
XFILLER_0_140_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15123_ _05180_ _05291_ _05400_ VGND VGND VPWR VPWR _05401_ sky130_fd_sc_hd__a21bo_2
X_12335_ _02355_ _02354_ VGND VGND VPWR VPWR _02428_ sky130_fd_sc_hd__and2b_1
XFILLER_0_106_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15054_ _05312_ _05313_ _05323_ VGND VGND VPWR VPWR _05325_ sky130_fd_sc_hd__and3_1
XFILLER_0_50_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12266_ _05595_ _00180_ _00130_ _06019_ VGND VGND VPWR VPWR _02359_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_687 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14005_ _04178_ _04179_ VGND VGND VPWR VPWR _04180_ sky130_fd_sc_hd__xnor2_1
X_11217_ _01290_ _01308_ _01309_ VGND VGND VPWR VPWR _01310_ sky130_fd_sc_hd__or3_4
Xoutput70 net70 VGND VGND VPWR VPWR leds[0] sky130_fd_sc_hd__buf_2
X_12197_ _02288_ _02203_ _02289_ VGND VGND VPWR VPWR _02290_ sky130_fd_sc_hd__and3_1
XFILLER_0_120_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_128_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput81 net81 VGND VGND VPWR VPWR leds[9] sky130_fd_sc_hd__clkbuf_4
X_18813_ _09298_ _09319_ VGND VGND VPWR VPWR _09320_ sky130_fd_sc_hd__and2_1
Xoutput92 net92 VGND VGND VPWR VPWR o_wb_data[18] sky130_fd_sc_hd__clkbuf_4
X_11148_ _00702_ _00169_ _07559_ _07602_ VGND VGND VPWR VPWR _01241_ sky130_fd_sc_hd__and4_1
XFILLER_0_128_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18744_ _09265_ VGND VGND VPWR VPWR _00073_ sky130_fd_sc_hd__clkbuf_1
X_11079_ _04646_ _04373_ _03432_ _00205_ VGND VGND VPWR VPWR _01172_ sky130_fd_sc_hd__nand4_2
X_15956_ _06200_ _06246_ VGND VGND VPWR VPWR _06303_ sky130_fd_sc_hd__nand2_1
X_14907_ _05163_ _05164_ VGND VGND VPWR VPWR _05165_ sky130_fd_sc_hd__nor2_1
X_18675_ _02259_ _09190_ _09191_ VGND VGND VPWR VPWR _09215_ sky130_fd_sc_hd__a21oi_1
X_15887_ _04828_ _05307_ _06229_ _03039_ VGND VGND VPWR VPWR _06230_ sky130_fd_sc_hd__o22a_1
X_17626_ _08009_ _08042_ _08118_ VGND VGND VPWR VPWR _08120_ sky130_fd_sc_hd__nor3_2
XFILLER_0_59_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14838_ _03539_ _05089_ VGND VGND VPWR VPWR _05090_ sky130_fd_sc_hd__nor2_1
XFILLER_0_58_332 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_129_710 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17557_ _07942_ _07949_ VGND VGND VPWR VPWR _08044_ sky130_fd_sc_hd__nor2_1
X_14769_ _04867_ _04968_ _05012_ _05013_ VGND VGND VPWR VPWR _05014_ sky130_fd_sc_hd__a211o_1
XFILLER_0_46_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16508_ _06834_ _06900_ VGND VGND VPWR VPWR _06902_ sky130_fd_sc_hd__or2b_1
X_17488_ _07965_ _07967_ VGND VGND VPWR VPWR _07969_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_129_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_128_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16439_ _06825_ _06826_ VGND VGND VPWR VPWR _06827_ sky130_fd_sc_hd__nand2_1
XFILLER_0_144_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18109_ _08636_ _08644_ VGND VGND VPWR VPWR _08645_ sky130_fd_sc_hd__xor2_1
XFILLER_0_78_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09813_ _07330_ _07461_ VGND VGND VPWR VPWR _07472_ sky130_fd_sc_hd__xnor2_2
X_09744_ cla_inst.in1\[24\] VGND VGND VPWR VPWR _06722_ sky130_fd_sc_hd__clkbuf_4
X_09675_ _05964_ VGND VGND VPWR VPWR _05975_ sky130_fd_sc_hd__clkbuf_8
XTAP_2007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_696 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_147_540 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_622 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_107_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10450_ _00356_ _00364_ _00355_ VGND VGND VPWR VPWR _00543_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_122_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_150_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10381_ _00472_ _00473_ VGND VGND VPWR VPWR _00474_ sky130_fd_sc_hd__nor2_1
XFILLER_0_60_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12120_ _02211_ _02212_ _05671_ _00205_ VGND VGND VPWR VPWR _02213_ sky130_fd_sc_hd__and4b_1
XFILLER_0_103_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12051_ _02140_ _02142_ VGND VGND VPWR VPWR _02144_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_2_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11002_ _07069_ net232 net221 _07984_ VGND VGND VPWR VPWR _01095_ sky130_fd_sc_hd__a22o_1
X_15810_ _03536_ _06146_ _03123_ VGND VGND VPWR VPWR _06147_ sky130_fd_sc_hd__a21o_1
X_16790_ _06762_ _06947_ _07207_ _06655_ VGND VGND VPWR VPWR _07208_ sky130_fd_sc_hd__a22o_1
X_15741_ _06006_ _06010_ _06070_ VGND VGND VPWR VPWR _06072_ sky130_fd_sc_hd__or3_1
X_12953_ _03024_ _03045_ VGND VGND VPWR VPWR _03046_ sky130_fd_sc_hd__nand2_1
X_11904_ _01992_ _01994_ VGND VGND VPWR VPWR _01997_ sky130_fd_sc_hd__xnor2_4
X_15672_ _05991_ _05996_ VGND VGND VPWR VPWR _05998_ sky130_fd_sc_hd__or2_2
X_18460_ _02938_ _09023_ _09024_ VGND VGND VPWR VPWR _09025_ sky130_fd_sc_hd__a21oi_2
X_12884_ _07091_ VGND VGND VPWR VPWR _02977_ sky130_fd_sc_hd__buf_4
XTAP_2530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14623_ _04714_ _04717_ _04715_ VGND VGND VPWR VPWR _04855_ sky130_fd_sc_hd__o21ba_1
XTAP_2563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17411_ _07742_ _07747_ _07884_ VGND VGND VPWR VPWR _07885_ sky130_fd_sc_hd__a21oi_1
X_11835_ _01926_ _01927_ VGND VGND VPWR VPWR _01928_ sky130_fd_sc_hd__nor2_1
X_18391_ _04853_ _08895_ _08896_ _08948_ _08949_ VGND VGND VPWR VPWR _08950_ sky130_fd_sc_hd__a221o_1
XTAP_2574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17342_ _02200_ _06547_ _06550_ VGND VGND VPWR VPWR _07811_ sky130_fd_sc_hd__a21o_1
X_14554_ _00115_ _01866_ _04658_ _04656_ VGND VGND VPWR VPWR _04780_ sky130_fd_sc_hd__a31o_1
XTAP_1873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11766_ _01845_ _01858_ VGND VGND VPWR VPWR _01859_ sky130_fd_sc_hd__or2_4
XTAP_1884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13505_ _05508_ _05366_ _07374_ _07406_ VGND VGND VPWR VPWR _03633_ sky130_fd_sc_hd__nand4_2
X_10717_ _00805_ _00809_ VGND VGND VPWR VPWR _00810_ sky130_fd_sc_hd__and2_1
X_17273_ _07731_ _07734_ VGND VGND VPWR VPWR _07735_ sky130_fd_sc_hd__or2b_1
X_14485_ _04584_ _04585_ _04595_ VGND VGND VPWR VPWR _04704_ sky130_fd_sc_hd__nor3_1
XFILLER_0_99_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11697_ _01760_ _01769_ _01236_ _01789_ VGND VGND VPWR VPWR _01790_ sky130_fd_sc_hd__o211a_4
XFILLER_0_126_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19012_ clknet_4_9_0_clk _00102_ VGND VGND VPWR VPWR op_code\[1\] sky130_fd_sc_hd__dfxtp_1
X_16224_ _06551_ VGND VGND VPWR VPWR _06594_ sky130_fd_sc_hd__clkbuf_4
X_13436_ _03539_ _03548_ _03557_ VGND VGND VPWR VPWR _03558_ sky130_fd_sc_hd__a21oi_1
X_10648_ _00529_ _00699_ _00739_ _00740_ VGND VGND VPWR VPWR _00741_ sky130_fd_sc_hd__o211a_1
XFILLER_0_70_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrebuffer3 _06548_ VGND VGND VPWR VPWR net166 sky130_fd_sc_hd__buf_1
XFILLER_0_130_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16155_ _01151_ ApproximateM_inst.lob_16.lob2.genblk1\[14\].genblk1.mux.sel _04340_
+ _04362_ VGND VGND VPWR VPWR _06519_ sky130_fd_sc_hd__or4_1
X_13367_ _03480_ _03481_ VGND VGND VPWR VPWR _03482_ sky130_fd_sc_hd__or2_1
X_10579_ _00667_ _00670_ _00671_ VGND VGND VPWR VPWR _00672_ sky130_fd_sc_hd__and3_1
XFILLER_0_106_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15106_ _01873_ _03149_ _05380_ VGND VGND VPWR VPWR _05382_ sky130_fd_sc_hd__a21o_1
X_12318_ _02405_ _02409_ _02410_ VGND VGND VPWR VPWR _02411_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_23_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16086_ _04336_ _03041_ _06443_ VGND VGND VPWR VPWR _06444_ sky130_fd_sc_hd__and3_1
X_13298_ _03393_ _03394_ _03405_ VGND VGND VPWR VPWR _03406_ sky130_fd_sc_hd__o21ai_2
X_15037_ _03117_ _03199_ VGND VGND VPWR VPWR _05307_ sky130_fd_sc_hd__nand2_4
X_12249_ _02339_ _02341_ VGND VGND VPWR VPWR _02342_ sky130_fd_sc_hd__nand2_1
XFILLER_0_139_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_88 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16988_ _07415_ _07423_ VGND VGND VPWR VPWR _07424_ sky130_fd_sc_hd__xor2_1
XFILLER_0_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18727_ _06477_ net35 _09251_ VGND VGND VPWR VPWR _09252_ sky130_fd_sc_hd__mux2_1
X_15939_ _06219_ _06260_ VGND VGND VPWR VPWR _06285_ sky130_fd_sc_hd__or2_1
X_09460_ _03345_ VGND VGND VPWR VPWR _03629_ sky130_fd_sc_hd__buf_4
X_18658_ _09176_ _09201_ VGND VGND VPWR VPWR _09202_ sky130_fd_sc_hd__and2_1
X_17609_ _08099_ _08100_ VGND VGND VPWR VPWR _08101_ sky130_fd_sc_hd__or2_1
X_18589_ salida\[14\] _09141_ _09142_ salida\[46\] _09146_ VGND VGND VPWR VPWR _09150_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_19_538 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_563 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_140_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09727_ _06373_ _06515_ _06504_ VGND VGND VPWR VPWR _06537_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_69_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09658_ _05725_ _05780_ VGND VGND VPWR VPWR _05791_ sky130_fd_sc_hd__nor2_1
XFILLER_0_69_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09589_ _05028_ VGND VGND VPWR VPWR _05039_ sky130_fd_sc_hd__buf_6
XTAP_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11620_ _01192_ _01711_ _01712_ VGND VGND VPWR VPWR _01713_ sky130_fd_sc_hd__nand3_2
XFILLER_0_154_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_148_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11551_ _07243_ ApproximateM_inst.lob_16.lob1.genblk2.mux_final.sel ApproximateM_inst.lob_16.lob1.genblk1\[14\].genblk1.mux.sel
+ _07221_ VGND VGND VPWR VPWR _01644_ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10502_ _00587_ _00588_ _00427_ _00430_ VGND VGND VPWR VPWR _00595_ sky130_fd_sc_hd__a211oi_1
X_14270_ _04461_ _04462_ _04467_ VGND VGND VPWR VPWR _04469_ sky130_fd_sc_hd__a21o_1
XFILLER_0_123_705 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11482_ _08409_ VGND VGND VPWR VPWR _01575_ sky130_fd_sc_hd__buf_8
X_13221_ _03321_ _00212_ _00206_ _03322_ VGND VGND VPWR VPWR _03323_ sky130_fd_sc_hd__a22oi_1
X_10433_ _00524_ _00525_ VGND VGND VPWR VPWR _00526_ sky130_fd_sc_hd__nand2_2
XFILLER_0_33_596 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13152_ _00645_ _07156_ _06732_ _05453_ VGND VGND VPWR VPWR _03250_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10364_ _00453_ _00455_ _00454_ VGND VGND VPWR VPWR _00457_ sky130_fd_sc_hd__a21o_1
XFILLER_0_103_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12103_ _02193_ _02194_ VGND VGND VPWR VPWR _02196_ sky130_fd_sc_hd__nand2_1
XTAP_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13083_ _03025_ _03101_ VGND VGND VPWR VPWR _03175_ sky130_fd_sc_hd__and2_1
X_17960_ _08363_ _08450_ _08481_ VGND VGND VPWR VPWR _08483_ sky130_fd_sc_hd__nand3_1
X_10295_ _00109_ _09349_ _00177_ _00146_ VGND VGND VPWR VPWR _00388_ sky130_fd_sc_hd__and4_1
X_12034_ _00715_ VGND VGND VPWR VPWR _02127_ sky130_fd_sc_hd__clkinv_4
X_16911_ _07231_ _07239_ _07229_ VGND VGND VPWR VPWR _07340_ sky130_fd_sc_hd__o21ai_1
X_17891_ _08405_ _08407_ VGND VGND VPWR VPWR _08408_ sky130_fd_sc_hd__xor2_1
X_16842_ _06358_ _06356_ _06357_ _07264_ VGND VGND VPWR VPWR _07266_ sky130_fd_sc_hd__o31a_1
X_13985_ _04151_ _04155_ _04157_ VGND VGND VPWR VPWR _04158_ sky130_fd_sc_hd__or3_1
X_16773_ _03094_ _06463_ _07190_ VGND VGND VPWR VPWR _09416_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_87_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18512_ _07256_ _09078_ _09079_ VGND VGND VPWR VPWR _09081_ sky130_fd_sc_hd__and3_1
X_15724_ _06052_ _06053_ VGND VGND VPWR VPWR _06054_ sky130_fd_sc_hd__nor2_1
X_12936_ _01357_ VGND VGND VPWR VPWR _03029_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_76_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18443_ _09004_ _09006_ VGND VGND VPWR VPWR _09007_ sky130_fd_sc_hd__or2_1
X_15655_ _01356_ _00665_ _05974_ _05976_ VGND VGND VPWR VPWR _05979_ sky130_fd_sc_hd__a22o_1
X_12867_ _02918_ _02937_ _02936_ VGND VGND VPWR VPWR _02960_ sky130_fd_sc_hd__a21oi_1
XTAP_2360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14606_ _01521_ _07112_ _04707_ _04708_ VGND VGND VPWR VPWR _04836_ sky130_fd_sc_hd__and4_1
X_11818_ _01909_ _01910_ VGND VGND VPWR VPWR _01911_ sky130_fd_sc_hd__nor2_1
X_15586_ _05895_ _05902_ VGND VGND VPWR VPWR _05904_ sky130_fd_sc_hd__nor2_1
X_18374_ _02892_ _08878_ VGND VGND VPWR VPWR _08933_ sky130_fd_sc_hd__nand2_2
XTAP_1670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12798_ _02172_ _02470_ _02851_ _02882_ _02890_ VGND VGND VPWR VPWR _02891_ sky130_fd_sc_hd__o311a_4
XFILLER_0_56_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14537_ _00189_ _00191_ _05257_ _05486_ VGND VGND VPWR VPWR _04761_ sky130_fd_sc_hd__and4_1
X_17325_ _07790_ _07791_ VGND VGND VPWR VPWR _07792_ sky130_fd_sc_hd__and2b_1
X_11749_ _01676_ _01679_ _01680_ _01670_ VGND VGND VPWR VPWR _01842_ sky130_fd_sc_hd__o31a_1
XFILLER_0_154_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14468_ _04683_ _04684_ _04685_ VGND VGND VPWR VPWR _04686_ sky130_fd_sc_hd__nor3_2
XFILLER_0_119_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17256_ _07714_ _07715_ VGND VGND VPWR VPWR _07716_ sky130_fd_sc_hd__xor2_1
XFILLER_0_36_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16207_ _04121_ _03717_ _04351_ VGND VGND VPWR VPWR _06575_ sky130_fd_sc_hd__or3_4
X_13419_ _03538_ VGND VGND VPWR VPWR _03539_ sky130_fd_sc_hd__clkbuf_4
X_17187_ _07502_ _07640_ VGND VGND VPWR VPWR _07641_ sky130_fd_sc_hd__xnor2_1
X_14399_ _04464_ _04465_ VGND VGND VPWR VPWR _04610_ sky130_fd_sc_hd__and2_1
XFILLER_0_113_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_141_568 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16138_ _01108_ _03136_ VGND VGND VPWR VPWR _06500_ sky130_fd_sc_hd__or2_1
XFILLER_0_12_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_76 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_122_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16069_ _06424_ VGND VGND VPWR VPWR _06425_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_121_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09512_ _03684_ _03585_ _03640_ VGND VGND VPWR VPWR _04198_ sky130_fd_sc_hd__nand3_1
XFILLER_0_78_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09443_ _03356_ _03377_ _03410_ _03432_ VGND VGND VPWR VPWR _03443_ sky130_fd_sc_hd__nand4_1
XPHY_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_136_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_117_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_131_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_749 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_104_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10080_ cla_inst.in2\[24\] VGND VGND VPWR VPWR _00173_ sky130_fd_sc_hd__clkbuf_4
X_13770_ _03538_ _03915_ _03922_ _06765_ VGND VGND VPWR VPWR _03923_ sky130_fd_sc_hd__o211a_1
X_10982_ _01072_ _01073_ _01061_ _01068_ VGND VGND VPWR VPWR _01075_ sky130_fd_sc_hd__a211o_1
X_12721_ _02804_ _02813_ VGND VGND VPWR VPWR _02814_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_69_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15440_ _05743_ _05744_ VGND VGND VPWR VPWR _05745_ sky130_fd_sc_hd__xnor2_1
X_12652_ _02742_ _02744_ VGND VGND VPWR VPWR _02745_ sky130_fd_sc_hd__and2_1
XFILLER_0_139_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11603_ _00515_ _01692_ VGND VGND VPWR VPWR _01696_ sky130_fd_sc_hd__nor2_4
X_15371_ _05668_ _05669_ VGND VGND VPWR VPWR _05670_ sky130_fd_sc_hd__or2_1
X_12583_ _01082_ _01081_ ApproximateM_inst.lob_16.lob1.genblk1\[1\].genblk1.mux.sel
+ VGND VGND VPWR VPWR _02676_ sky130_fd_sc_hd__and3_1
XFILLER_0_53_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14322_ _04512_ _04513_ _04524_ VGND VGND VPWR VPWR _04527_ sky130_fd_sc_hd__or3_1
X_17110_ _07345_ _07349_ _07447_ _07448_ VGND VGND VPWR VPWR _07557_ sky130_fd_sc_hd__o31a_1
XFILLER_0_135_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11534_ _05736_ _01005_ VGND VGND VPWR VPWR _01627_ sky130_fd_sc_hd__nand2_1
X_18090_ _08622_ _08623_ VGND VGND VPWR VPWR _08624_ sky130_fd_sc_hd__nand2_1
XFILLER_0_151_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17041_ _07481_ VGND VGND VPWR VPWR _09388_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14253_ _04515_ _04438_ _07755_ _07722_ VGND VGND VPWR VPWR _04451_ sky130_fd_sc_hd__and4_1
XFILLER_0_80_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11465_ _01159_ _01508_ VGND VGND VPWR VPWR _01558_ sky130_fd_sc_hd__nand2_1
XFILLER_0_151_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13204_ _01745_ _00716_ _03304_ VGND VGND VPWR VPWR _03305_ sky130_fd_sc_hd__nand3_1
XFILLER_0_21_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10416_ cla_inst.in1\[31\] VGND VGND VPWR VPWR _00509_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_33_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14184_ _04355_ _04356_ _04375_ VGND VGND VPWR VPWR _04376_ sky130_fd_sc_hd__a21o_1
X_11396_ _01466_ _01467_ _01394_ _01413_ VGND VGND VPWR VPWR _01489_ sky130_fd_sc_hd__a211o_1
XFILLER_0_60_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13135_ _05017_ _00308_ _03229_ _03230_ VGND VGND VPWR VPWR _03232_ sky130_fd_sc_hd__a22o_1
X_10347_ _03881_ _05028_ _00439_ VGND VGND VPWR VPWR _00440_ sky130_fd_sc_hd__and3_1
XFILLER_0_103_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18992_ clknet_4_6_0_clk _09358_ VGND VGND VPWR VPWR salida\[45\] sky130_fd_sc_hd__dfxtp_1
XTAP_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13066_ _03152_ _03157_ VGND VGND VPWR VPWR _03158_ sky130_fd_sc_hd__or2_1
X_17943_ _08458_ _08462_ VGND VGND VPWR VPWR _08465_ sky130_fd_sc_hd__or2_1
X_10278_ _00369_ _00368_ _08984_ _08930_ VGND VGND VPWR VPWR _00371_ sky130_fd_sc_hd__o211ai_2
X_12017_ _01082_ _01081_ _03388_ _00949_ VGND VGND VPWR VPWR _02110_ sky130_fd_sc_hd__and4_1
X_17874_ _08301_ _08303_ _08299_ VGND VGND VPWR VPWR _08390_ sky130_fd_sc_hd__a21bo_1
X_16825_ _07245_ _07246_ VGND VGND VPWR VPWR _07247_ sky130_fd_sc_hd__xor2_1
Xmax_cap1 _04218_ VGND VGND VPWR VPWR net319 sky130_fd_sc_hd__clkbuf_1
X_16756_ _02533_ _03094_ VGND VGND VPWR VPWR _07172_ sky130_fd_sc_hd__nand2_1
X_13968_ _04128_ _04129_ _04138_ VGND VGND VPWR VPWR _04139_ sky130_fd_sc_hd__a21oi_1
X_15707_ _05976_ _05978_ VGND VGND VPWR VPWR _06035_ sky130_fd_sc_hd__nand2_1
X_12919_ _07668_ VGND VGND VPWR VPWR _03012_ sky130_fd_sc_hd__buf_2
X_13899_ _03897_ _03899_ _04063_ VGND VGND VPWR VPWR _04064_ sky130_fd_sc_hd__a21oi_1
X_16687_ _06990_ _06991_ _06989_ VGND VGND VPWR VPWR _07097_ sky130_fd_sc_hd__a21o_1
XFILLER_0_61_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18426_ _06408_ _06449_ _06425_ VGND VGND VPWR VPWR _08989_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15638_ _03012_ _03142_ _03055_ _03010_ VGND VGND VPWR VPWR _05960_ sky130_fd_sc_hd__a22o_1
XTAP_2190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_146_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18357_ _08912_ _08913_ VGND VGND VPWR VPWR _08914_ sky130_fd_sc_hd__and2_1
X_15569_ _05883_ _03142_ _03015_ _05884_ VGND VGND VPWR VPWR _05885_ sky130_fd_sc_hd__and4b_1
XFILLER_0_127_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17308_ _07641_ _07620_ VGND VGND VPWR VPWR _07773_ sky130_fd_sc_hd__or2b_1
XFILLER_0_16_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_34 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18288_ _08835_ _08837_ _08838_ VGND VGND VPWR VPWR _08839_ sky130_fd_sc_hd__o21a_2
XFILLER_0_142_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17239_ _00786_ _06367_ _06369_ _07084_ _07697_ VGND VGND VPWR VPWR _07698_ sky130_fd_sc_hd__a311o_1
XFILLER_0_24_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_566 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09992_ _09287_ _09295_ _09318_ VGND VGND VPWR VPWR _09326_ sky130_fd_sc_hd__nand3_2
XFILLER_0_86_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_4_15_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_15_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_19_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09426_ _03217_ op_code\[2\] op_code\[3\] VGND VGND VPWR VPWR _03260_ sky130_fd_sc_hd__and3_1
XFILLER_0_75_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_820 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11250_ cla_inst.in2\[23\] _01031_ ApproximateM_inst.lob_16.lob1.genblk1\[1\].genblk1.mux.sel
+ cla_inst.in2\[24\] VGND VGND VPWR VPWR _01343_ sky130_fd_sc_hd__a22o_1
XFILLER_0_132_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10201_ _04416_ VGND VGND VPWR VPWR _00294_ sky130_fd_sc_hd__buf_6
XFILLER_0_30_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11181_ _00967_ _00976_ _00977_ VGND VGND VPWR VPWR _01274_ sky130_fd_sc_hd__nor3_1
XFILLER_0_31_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10132_ _00222_ _00224_ VGND VGND VPWR VPWR _00225_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_101_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10063_ _00144_ _00155_ VGND VGND VPWR VPWR _00156_ sky130_fd_sc_hd__xor2_1
X_14940_ _05078_ _05074_ _05075_ VGND VGND VPWR VPWR _05201_ sky130_fd_sc_hd__a21o_1
X_14871_ _03008_ _07515_ _06471_ _04591_ VGND VGND VPWR VPWR _05125_ sky130_fd_sc_hd__and4_1
XFILLER_0_98_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16610_ _02829_ _02828_ VGND VGND VPWR VPWR _07013_ sky130_fd_sc_hd__nand2_1
X_13822_ _03965_ _03978_ VGND VGND VPWR VPWR _03980_ sky130_fd_sc_hd__xnor2_1
X_17590_ _07950_ _07953_ VGND VGND VPWR VPWR _08080_ sky130_fd_sc_hd__and2_1
XFILLER_0_58_717 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13753_ _03738_ _03747_ _03902_ _02969_ VGND VGND VPWR VPWR _03905_ sky130_fd_sc_hd__a31o_1
X_16541_ _06756_ VGND VGND VPWR VPWR _06937_ sky130_fd_sc_hd__buf_2
X_10965_ _05213_ _04482_ VGND VGND VPWR VPWR _01058_ sky130_fd_sc_hd__nand2_2
X_12704_ _02772_ _02796_ VGND VGND VPWR VPWR _02797_ sky130_fd_sc_hd__nor2_1
XFILLER_0_128_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13684_ _03642_ _03644_ _03827_ VGND VGND VPWR VPWR _03829_ sky130_fd_sc_hd__or3_1
X_16472_ _06836_ _06842_ _06860_ _06862_ VGND VGND VPWR VPWR _06864_ sky130_fd_sc_hd__o211a_1
X_10896_ _00985_ _00988_ VGND VGND VPWR VPWR _00989_ sky130_fd_sc_hd__and2_1
X_18211_ _08753_ _08754_ _08755_ VGND VGND VPWR VPWR _08756_ sky130_fd_sc_hd__o21a_1
X_15423_ _05724_ _05726_ VGND VGND VPWR VPWR _05727_ sky130_fd_sc_hd__xnor2_1
X_12635_ _06084_ VGND VGND VPWR VPWR _02728_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_122_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15354_ _04125_ VGND VGND VPWR VPWR _05652_ sky130_fd_sc_hd__clkbuf_4
X_18142_ _02997_ _03052_ VGND VGND VPWR VPWR _08682_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12566_ _02615_ _02619_ _02621_ VGND VGND VPWR VPWR _02659_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_124_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14305_ _04494_ _04347_ _04506_ VGND VGND VPWR VPWR _04508_ sky130_fd_sc_hd__and3_1
X_11517_ _01607_ _01608_ _01609_ VGND VGND VPWR VPWR _01610_ sky130_fd_sc_hd__and3_2
X_15285_ _02996_ _09059_ _00322_ _02993_ VGND VGND VPWR VPWR _05577_ sky130_fd_sc_hd__a22oi_2
X_18073_ _02998_ _06511_ _01136_ VGND VGND VPWR VPWR _08607_ sky130_fd_sc_hd__a21o_1
XFILLER_0_81_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12497_ _02531_ _02583_ VGND VGND VPWR VPWR _02590_ sky130_fd_sc_hd__xnor2_2
X_14236_ _01521_ _05715_ _04430_ _04431_ VGND VGND VPWR VPWR _04432_ sky130_fd_sc_hd__and4_1
XFILLER_0_40_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17024_ _07462_ _07463_ _06507_ VGND VGND VPWR VPWR _07464_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_123_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11448_ _04504_ _00294_ _00205_ _00217_ VGND VGND VPWR VPWR _01541_ sky130_fd_sc_hd__nand4_2
XFILLER_0_151_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14167_ _04197_ _04203_ VGND VGND VPWR VPWR _04357_ sky130_fd_sc_hd__and2b_1
XFILLER_0_0_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11379_ _00865_ _01471_ VGND VGND VPWR VPWR _01472_ sky130_fd_sc_hd__nor2_2
XFILLER_0_21_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13118_ _03210_ _03211_ _03212_ VGND VGND VPWR VPWR _03213_ sky130_fd_sc_hd__nand3_1
XTAP_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14098_ _04279_ _04280_ VGND VGND VPWR VPWR _04281_ sky130_fd_sc_hd__xor2_1
X_18975_ clknet_4_5_0_clk _09406_ VGND VGND VPWR VPWR salida\[28\] sky130_fd_sc_hd__dfxtp_1
XTAP_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17926_ _08422_ _08426_ _08446_ _06723_ _01692_ VGND VGND VPWR VPWR _09398_ sky130_fd_sc_hd__o32a_1
X_13049_ _01108_ _03140_ _03023_ VGND VGND VPWR VPWR _03141_ sky130_fd_sc_hd__o21a_1
X_17857_ _07109_ _07780_ VGND VGND VPWR VPWR _08371_ sky130_fd_sc_hd__nand2_1
X_16808_ _07205_ _07227_ VGND VGND VPWR VPWR _07228_ sky130_fd_sc_hd__xnor2_1
X_17788_ _08194_ _08195_ _08295_ VGND VGND VPWR VPWR _08296_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_89_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16739_ _06749_ _06969_ _07055_ _07053_ VGND VGND VPWR VPWR _07153_ sky130_fd_sc_hd__a31o_1
XFILLER_0_89_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18409_ _08968_ _08967_ VGND VGND VPWR VPWR _08970_ sky130_fd_sc_hd__and2b_1
XFILLER_0_8_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_539 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_130_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_130_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09975_ _09166_ _09172_ _09188_ _07591_ VGND VGND VPWR VPWR _09197_ sky130_fd_sc_hd__and4_1
XFILLER_0_110_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10750_ _00842_ _00840_ _00837_ VGND VGND VPWR VPWR _00843_ sky130_fd_sc_hd__or3b_1
XFILLER_0_137_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10681_ ApproximateM_inst.lob_16.lob1.genblk1\[6\].genblk1.mux.sel VGND VGND VPWR
+ VPWR _00774_ sky130_fd_sc_hd__buf_4
XFILLER_0_82_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12420_ _02510_ _02512_ VGND VGND VPWR VPWR _02513_ sky130_fd_sc_hd__and2_1
XFILLER_0_137_479 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12351_ _02376_ _02442_ _02411_ VGND VGND VPWR VPWR _02444_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_62_274 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11302_ _01392_ _01393_ _01290_ _01379_ VGND VGND VPWR VPWR _01395_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_105_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15070_ _05330_ _05341_ VGND VGND VPWR VPWR _05342_ sky130_fd_sc_hd__nand2_1
X_12282_ _02260_ _02371_ VGND VGND VPWR VPWR _02375_ sky130_fd_sc_hd__and2_1
XFILLER_0_22_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14021_ _03987_ _03989_ VGND VGND VPWR VPWR _04197_ sky130_fd_sc_hd__nor2_1
X_11233_ _01085_ _01092_ _01325_ VGND VGND VPWR VPWR _01326_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_132_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11164_ _01255_ _01256_ VGND VGND VPWR VPWR _01257_ sky130_fd_sc_hd__nand2_1
X_10115_ _00188_ _00201_ VGND VGND VPWR VPWR _00208_ sky130_fd_sc_hd__xnor2_1
X_18760_ _09273_ _09277_ VGND VGND VPWR VPWR _09278_ sky130_fd_sc_hd__and2_1
X_11095_ _01056_ _01182_ _01186_ VGND VGND VPWR VPWR _01188_ sky130_fd_sc_hd__a21o_1
X_15972_ _06308_ _06310_ VGND VGND VPWR VPWR _06320_ sky130_fd_sc_hd__nand2_1
X_17711_ _08102_ _08110_ _08101_ VGND VGND VPWR VPWR _08212_ sky130_fd_sc_hd__a21boi_2
X_14923_ _05180_ _05182_ VGND VGND VPWR VPWR _05183_ sky130_fd_sc_hd__nor2_1
X_10046_ _00123_ _00138_ VGND VGND VPWR VPWR _00139_ sky130_fd_sc_hd__or2_1
X_18691_ _09209_ _09224_ VGND VGND VPWR VPWR _09225_ sky130_fd_sc_hd__and2_1
XFILLER_0_26_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17642_ _06382_ _06380_ _06381_ _07084_ _08136_ VGND VGND VPWR VPWR _08138_ sky130_fd_sc_hd__a311o_1
Xhold92 net92 VGND VGND VPWR VPWR net255 sky130_fd_sc_hd__dlygate4sd3_1
X_14854_ _02984_ _01520_ _07733_ _08158_ VGND VGND VPWR VPWR _05107_ sky130_fd_sc_hd__and4_1
XFILLER_0_26_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13805_ _03949_ _03950_ _03960_ VGND VGND VPWR VPWR _03961_ sky130_fd_sc_hd__o21ai_2
X_17573_ _08054_ _08061_ VGND VGND VPWR VPWR _08062_ sky130_fd_sc_hd__xnor2_1
X_14785_ _04906_ _04914_ _05031_ VGND VGND VPWR VPWR _05032_ sky130_fd_sc_hd__a21oi_1
X_11997_ _02088_ _02089_ VGND VGND VPWR VPWR _02090_ sky130_fd_sc_hd__nor2_1
XFILLER_0_86_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16524_ _06547_ VGND VGND VPWR VPWR _06920_ sky130_fd_sc_hd__clkbuf_4
X_13736_ _03434_ _03586_ _03671_ _03672_ VGND VGND VPWR VPWR _03886_ sky130_fd_sc_hd__o211a_1
X_10948_ ApproximateM_inst.lob_16.lob2.genblk1\[11\].genblk1.mux.sel _03837_ VGND
+ VGND VPWR VPWR _01041_ sky130_fd_sc_hd__nand2_4
XFILLER_0_42_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16455_ _03098_ _06467_ _06501_ _06844_ VGND VGND VPWR VPWR _06845_ sky130_fd_sc_hd__a31o_1
X_13667_ _03786_ _03787_ _03807_ _03808_ VGND VGND VPWR VPWR _03810_ sky130_fd_sc_hd__and4bb_1
X_10879_ _00970_ _00971_ VGND VGND VPWR VPWR _00972_ sky130_fd_sc_hd__nor2_1
XFILLER_0_73_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15406_ _05626_ _05628_ _05707_ VGND VGND VPWR VPWR _05709_ sky130_fd_sc_hd__a21o_1
XFILLER_0_143_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12618_ _02683_ _02684_ _02690_ VGND VGND VPWR VPWR _02711_ sky130_fd_sc_hd__o21ai_1
X_13598_ _03482_ _03483_ _03486_ _03734_ VGND VGND VPWR VPWR _03735_ sky130_fd_sc_hd__a31oi_2
X_16386_ _06757_ _06768_ VGND VGND VPWR VPWR _06770_ sky130_fd_sc_hd__or2_1
XFILLER_0_26_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_606 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18125_ _08490_ VGND VGND VPWR VPWR _08663_ sky130_fd_sc_hd__inv_2
XFILLER_0_143_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15337_ _09351_ _07123_ _00318_ _02991_ VGND VGND VPWR VPWR _05633_ sky130_fd_sc_hd__a22o_1
X_12549_ _02602_ _02601_ _02598_ VGND VGND VPWR VPWR _02642_ sky130_fd_sc_hd__a21o_1
XFILLER_0_41_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18056_ _08410_ _08447_ _08504_ VGND VGND VPWR VPWR _08588_ sky130_fd_sc_hd__o21ai_1
XANTENNA_1 _00042_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15268_ _03322_ _09351_ _00309_ VGND VGND VPWR VPWR _05558_ sky130_fd_sc_hd__and3_1
XFILLER_0_77_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17007_ _07381_ _07336_ _07443_ _07444_ VGND VGND VPWR VPWR _07445_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_1_544 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_112_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14219_ _03034_ _03100_ _03081_ VGND VGND VPWR VPWR _04413_ sky130_fd_sc_hd__mux2_1
X_15199_ _05481_ _05482_ VGND VGND VPWR VPWR _05483_ sky130_fd_sc_hd__nor2_1
XFILLER_0_111_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09760_ _06548_ _06863_ _06873_ _06884_ VGND VGND VPWR VPWR _06895_ sky130_fd_sc_hd__and4b_1
XTAP_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18958_ clknet_4_6_0_clk _09388_ VGND VGND VPWR VPWR salida\[11\] sky130_fd_sc_hd__dfxtp_1
XTAP_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17909_ _07355_ VGND VGND VPWR VPWR _08428_ sky130_fd_sc_hd__buf_2
X_09691_ _05812_ _05823_ _05943_ _06138_ VGND VGND VPWR VPWR _06149_ sky130_fd_sc_hd__o211ai_2
X_18889_ clknet_4_9_0_clk _00043_ VGND VGND VPWR VPWR ApproximateM_inst.lob_16.lob1.genblk1\[7\].genblk1.mux.sel
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_83_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrebuffer13 _01957_ VGND VGND VPWR VPWR net176 sky130_fd_sc_hd__clkbuf_1
Xrebuffer24 _02118_ VGND VGND VPWR VPWR net187 sky130_fd_sc_hd__clkbuf_1
Xrebuffer35 _01769_ VGND VGND VPWR VPWR net198 sky130_fd_sc_hd__buf_2
Xrebuffer46 ApproximateM_inst.lob_16.lob1.genblk1\[11\].genblk1.mux.sel VGND VGND
+ VPWR VPWR net209 sky130_fd_sc_hd__clkbuf_1
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer57 _00980_ VGND VGND VPWR VPWR net220 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer68 net233 VGND VGND VPWR VPWR net231 sky130_fd_sc_hd__clkbuf_1
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer79 net172 VGND VGND VPWR VPWR net242 sky130_fd_sc_hd__buf_1
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_789 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_130_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09958_ _07330_ _07461_ VGND VGND VPWR VPWR _09048_ sky130_fd_sc_hd__nand2_1
X_09889_ _06906_ _06928_ _05181_ _06181_ VGND VGND VPWR VPWR _08300_ sky130_fd_sc_hd__o211ai_1
X_11920_ _05290_ _00176_ _00145_ _00806_ VGND VGND VPWR VPWR _02013_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_87_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11851_ _01919_ _01941_ _01943_ VGND VGND VPWR VPWR _01944_ sky130_fd_sc_hd__a21oi_2
XTAP_2734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10802_ _00231_ _00857_ _00894_ _00859_ _00888_ VGND VGND VPWR VPWR _00895_ sky130_fd_sc_hd__a32o_1
XTAP_2778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14570_ _04794_ _04795_ _04775_ VGND VGND VPWR VPWR _04797_ sky130_fd_sc_hd__o21a_1
XFILLER_0_79_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11782_ _01742_ _01874_ VGND VGND VPWR VPWR _01875_ sky130_fd_sc_hd__nor2_1
XTAP_2789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13521_ _03647_ _03648_ _03408_ _03433_ VGND VGND VPWR VPWR _03650_ sky130_fd_sc_hd__o211a_1
X_10733_ _08126_ _08137_ _08256_ VGND VGND VPWR VPWR _00826_ sky130_fd_sc_hd__and3_1
XFILLER_0_82_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16240_ _06467_ _06610_ VGND VGND VPWR VPWR _06611_ sky130_fd_sc_hd__nand2_1
X_13452_ _03171_ _03174_ _03048_ VGND VGND VPWR VPWR _03575_ sky130_fd_sc_hd__mux2_1
X_10664_ _00590_ _00597_ _00756_ VGND VGND VPWR VPWR _00757_ sky130_fd_sc_hd__a21oi_1
X_12403_ _02495_ VGND VGND VPWR VPWR _02496_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13383_ _03497_ _03499_ VGND VGND VPWR VPWR _03500_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16171_ _03281_ sel_op\[3\] VGND VGND VPWR VPWR _06536_ sky130_fd_sc_hd__or2b_1
X_10595_ _00676_ _00677_ _00687_ VGND VGND VPWR VPWR _00688_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_152_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15122_ _05289_ _05288_ VGND VGND VPWR VPWR _05400_ sky130_fd_sc_hd__or2b_1
X_12334_ _07352_ _00211_ VGND VGND VPWR VPWR _02427_ sky130_fd_sc_hd__nand2_1
XFILLER_0_50_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15053_ _05312_ _05313_ _05323_ VGND VGND VPWR VPWR _05324_ sky130_fd_sc_hd__a21oi_1
X_12265_ ApproximateM_inst.lob_16.lob2.genblk1\[5\].genblk1.mux.sel _00909_ VGND VGND
+ VPWR VPWR _02358_ sky130_fd_sc_hd__and2_2
XFILLER_0_120_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14004_ _00253_ _06482_ VGND VGND VPWR VPWR _04179_ sky130_fd_sc_hd__nand2_1
X_11216_ _01288_ _01289_ _00967_ _01274_ VGND VGND VPWR VPWR _01309_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_121_699 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12196_ _02144_ _02145_ VGND VGND VPWR VPWR _02289_ sky130_fd_sc_hd__or2_1
Xoutput71 net71 VGND VGND VPWR VPWR leds[10] sky130_fd_sc_hd__buf_2
Xoutput82 net82 VGND VGND VPWR VPWR o_wb_ack sky130_fd_sc_hd__clkbuf_4
X_18812_ _02992_ net54 _09301_ VGND VGND VPWR VPWR _09319_ sky130_fd_sc_hd__mux2_1
X_11147_ _01239_ VGND VGND VPWR VPWR _01240_ sky130_fd_sc_hd__inv_2
Xoutput93 net93 VGND VGND VPWR VPWR o_wb_data[19] sky130_fd_sc_hd__clkbuf_4
X_18743_ _09245_ _09264_ VGND VGND VPWR VPWR _09265_ sky130_fd_sc_hd__and2_1
X_11078_ _01167_ _01170_ VGND VGND VPWR VPWR _01171_ sky130_fd_sc_hd__xor2_2
X_15955_ _06248_ VGND VGND VPWR VPWR _06302_ sky130_fd_sc_hd__inv_2
X_14906_ _00190_ _05986_ _05162_ VGND VGND VPWR VPWR _05164_ sky130_fd_sc_hd__and3_1
X_10029_ _07853_ _00119_ _00121_ VGND VGND VPWR VPWR _00122_ sky130_fd_sc_hd__nand3_4
X_18674_ _09214_ VGND VGND VPWR VPWR _00047_ sky130_fd_sc_hd__buf_1
XFILLER_0_78_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15886_ _04826_ _04827_ _03537_ VGND VGND VPWR VPWR _06229_ sky130_fd_sc_hd__mux2_1
X_17625_ _08009_ _08042_ _08118_ VGND VGND VPWR VPWR _08119_ sky130_fd_sc_hd__o21a_1
X_14837_ _05087_ _05088_ _03916_ VGND VGND VPWR VPWR _05089_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_480 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17556_ _07938_ _07941_ VGND VGND VPWR VPWR _08043_ sky130_fd_sc_hd__nor2_1
X_14768_ _04999_ _05000_ _05011_ VGND VGND VPWR VPWR _05013_ sky130_fd_sc_hd__and3_1
XFILLER_0_58_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16507_ _06866_ _06900_ VGND VGND VPWR VPWR _06901_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_128_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13719_ _03865_ _03866_ VGND VGND VPWR VPWR _03867_ sky130_fd_sc_hd__nor2_1
X_17487_ _07965_ _07967_ VGND VGND VPWR VPWR _07968_ sky130_fd_sc_hd__or2_1
X_14699_ _04936_ _04937_ VGND VGND VPWR VPWR _04938_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_129_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16438_ _06749_ _06763_ VGND VGND VPWR VPWR _06826_ sky130_fd_sc_hd__nand2_2
XFILLER_0_144_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_144_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16369_ _04121_ _03281_ VGND VGND VPWR VPWR _06751_ sky130_fd_sc_hd__and2_1
XFILLER_0_82_892 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18108_ _08641_ _08643_ VGND VGND VPWR VPWR _08644_ sky130_fd_sc_hd__nor2_1
XFILLER_0_143_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18039_ _08477_ _08566_ _08567_ VGND VGND VPWR VPWR _08569_ sky130_fd_sc_hd__nand3_1
XFILLER_0_41_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09812_ _07341_ _07450_ VGND VGND VPWR VPWR _07461_ sky130_fd_sc_hd__xor2_2
XFILLER_0_10_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09743_ _05671_ VGND VGND VPWR VPWR _06711_ sky130_fd_sc_hd__buf_4
X_09674_ _05606_ VGND VGND VPWR VPWR _05964_ sky130_fd_sc_hd__buf_4
XTAP_2008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_720 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_119_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_107_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_391 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10380_ _05235_ _07134_ _00470_ _00471_ VGND VGND VPWR VPWR _00473_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_32_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12050_ _02140_ _02142_ VGND VGND VPWR VPWR _02143_ sky130_fd_sc_hd__and2b_1
X_11001_ _07036_ _07069_ _08049_ net221 VGND VGND VPWR VPWR _01094_ sky130_fd_sc_hd__nand4_2
X_15740_ _06006_ _06010_ _06070_ VGND VGND VPWR VPWR _06071_ sky130_fd_sc_hd__o21ai_2
X_12952_ _03027_ _03044_ _01696_ VGND VGND VPWR VPWR _03045_ sky130_fd_sc_hd__a21o_1
X_11903_ _01810_ _01903_ VGND VGND VPWR VPWR _01996_ sky130_fd_sc_hd__nor2_1
XFILLER_0_59_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15671_ _05994_ _05995_ VGND VGND VPWR VPWR _05996_ sky130_fd_sc_hd__nand2_1
XTAP_2520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12883_ _02975_ VGND VGND VPWR VPWR _02976_ sky130_fd_sc_hd__buf_2
XTAP_2531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17410_ _07738_ _07764_ _07762_ VGND VGND VPWR VPWR _07884_ sky130_fd_sc_hd__a21oi_1
X_14622_ _04849_ _04850_ _04851_ VGND VGND VPWR VPWR _04854_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_68_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11834_ _01920_ _01921_ _01925_ VGND VGND VPWR VPWR _01927_ sky130_fd_sc_hd__o21ba_1
X_18390_ _08896_ _08947_ VGND VGND VPWR VPWR _08949_ sky130_fd_sc_hd__nor2_1
XTAP_2564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17341_ _06440_ _07808_ VGND VGND VPWR VPWR _07809_ sky130_fd_sc_hd__nor2_1
X_14553_ _04653_ _04661_ VGND VGND VPWR VPWR _04779_ sky130_fd_sc_hd__and2_1
XFILLER_0_68_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11765_ _01848_ _01856_ _01857_ VGND VGND VPWR VPWR _01858_ sky130_fd_sc_hd__a21oi_1
XTAP_1874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13504_ _05301_ cla_inst.in1\[27\] _07004_ _05279_ VGND VGND VPWR VPWR _03632_ sky130_fd_sc_hd__a22o_1
X_10716_ _08724_ _06482_ _00807_ _00808_ VGND VGND VPWR VPWR _00809_ sky130_fd_sc_hd__a31o_1
XFILLER_0_71_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_126_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_138_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17272_ _07703_ _07704_ _07732_ VGND VGND VPWR VPWR _07734_ sky130_fd_sc_hd__or3b_1
X_14484_ _04586_ _04594_ VGND VGND VPWR VPWR _04703_ sky130_fd_sc_hd__nand2_1
X_11696_ _01233_ _01234_ _01235_ _01204_ VGND VGND VPWR VPWR _01789_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_36_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19011_ clknet_4_9_0_clk _00101_ VGND VGND VPWR VPWR op_code\[0\] sky130_fd_sc_hd__dfxtp_2
X_16223_ _06592_ VGND VGND VPWR VPWR _06593_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_153_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10647_ _00737_ _00738_ _00718_ VGND VGND VPWR VPWR _00740_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_64_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13435_ _03538_ _03556_ VGND VGND VPWR VPWR _03557_ sky130_fd_sc_hd__nor2_1
XFILLER_0_126_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_130_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer4 net166 VGND VGND VPWR VPWR net167 sky130_fd_sc_hd__buf_1
X_13366_ _00877_ _03311_ VGND VGND VPWR VPWR _03481_ sky130_fd_sc_hd__nand2_1
X_16154_ _05213_ _03004_ _03019_ _06517_ VGND VGND VPWR VPWR _06518_ sky130_fd_sc_hd__or4_1
X_10578_ _06982_ _00509_ _00668_ _00669_ VGND VGND VPWR VPWR _00671_ sky130_fd_sc_hd__a22o_1
X_15105_ _00591_ _03149_ _05380_ VGND VGND VPWR VPWR _05381_ sky130_fd_sc_hd__nand3_1
XFILLER_0_51_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12317_ _02339_ _02341_ VGND VGND VPWR VPWR _02410_ sky130_fd_sc_hd__xnor2_1
X_13297_ _03395_ _03404_ VGND VGND VPWR VPWR _03405_ sky130_fd_sc_hd__xnor2_2
X_16085_ _01678_ _06442_ VGND VGND VPWR VPWR _06443_ sky130_fd_sc_hd__and2_1
XFILLER_0_121_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12248_ _02340_ _02335_ VGND VGND VPWR VPWR _02341_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_121_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15036_ _04243_ _04245_ _04247_ VGND VGND VPWR VPWR _05306_ sky130_fd_sc_hd__mux2_2
XFILLER_0_139_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12179_ _01113_ _02045_ VGND VGND VPWR VPWR _02272_ sky130_fd_sc_hd__nor2_2
X_16987_ _07421_ _07422_ VGND VGND VPWR VPWR _07423_ sky130_fd_sc_hd__xnor2_1
X_18726_ _09250_ VGND VGND VPWR VPWR _09251_ sky130_fd_sc_hd__clkbuf_4
X_15938_ _06282_ _06283_ VGND VGND VPWR VPWR _06284_ sky130_fd_sc_hd__or2_2
X_18657_ net63 _03169_ _09193_ VGND VGND VPWR VPWR _09201_ sky130_fd_sc_hd__mux2_1
X_15869_ _06095_ _06165_ _06167_ VGND VGND VPWR VPWR _06210_ sky130_fd_sc_hd__o21a_1
X_17608_ _07969_ _07994_ _07968_ VGND VGND VPWR VPWR _08100_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_149_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18588_ net299 _09140_ _09149_ _09144_ VGND VGND VPWR VPWR _00017_ sky130_fd_sc_hd__o211a_1
XFILLER_0_148_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17539_ _08023_ _08024_ VGND VGND VPWR VPWR _08025_ sky130_fd_sc_hd__and2_1
XFILLER_0_74_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_129_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_105_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_496 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09726_ _06373_ _06504_ _06515_ VGND VGND VPWR VPWR _06526_ sky130_fd_sc_hd__and3_1
XFILLER_0_97_704 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09657_ _05747_ _05758_ _05769_ _05660_ VGND VGND VPWR VPWR _05780_ sky130_fd_sc_hd__a22oi_1
XTAP_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09588_ cla_inst.in1\[17\] VGND VGND VPWR VPWR _05028_ sky130_fd_sc_hd__buf_4
XTAP_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11550_ _07984_ _07973_ _04449_ _04471_ VGND VGND VPWR VPWR _01643_ sky130_fd_sc_hd__nand4_2
XFILLER_0_107_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10501_ _00592_ _00593_ _00413_ _00412_ VGND VGND VPWR VPWR _00594_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_108_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11481_ _01568_ _01569_ _01572_ VGND VGND VPWR VPWR _01574_ sky130_fd_sc_hd__a21o_1
XFILLER_0_107_257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_135_566 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_150_503 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_123_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13220_ _00151_ VGND VGND VPWR VPWR _03322_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_122_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10432_ _00519_ _00523_ VGND VGND VPWR VPWR _00525_ sky130_fd_sc_hd__or2_1
X_13151_ _08724_ _07123_ _00647_ _00648_ VGND VGND VPWR VPWR _03249_ sky130_fd_sc_hd__and4_1
XFILLER_0_20_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10363_ _00453_ _00454_ _00455_ VGND VGND VPWR VPWR _00456_ sky130_fd_sc_hd__and3_1
X_12102_ _02193_ _02194_ VGND VGND VPWR VPWR _02195_ sky130_fd_sc_hd__or2_1
XFILLER_0_131_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13082_ _02607_ _03173_ _03040_ VGND VGND VPWR VPWR _03174_ sky130_fd_sc_hd__o21ai_1
X_10294_ _00125_ _00178_ _00181_ _00151_ VGND VGND VPWR VPWR _00387_ sky130_fd_sc_hd__a22oi_1
X_12033_ _07711_ _02124_ _02125_ VGND VGND VPWR VPWR _02126_ sky130_fd_sc_hd__and3_2
X_16910_ _07331_ _07338_ VGND VGND VPWR VPWR _07339_ sky130_fd_sc_hd__xor2_1
X_17890_ _08296_ _08310_ _08406_ VGND VGND VPWR VPWR _08407_ sky130_fd_sc_hd__a21bo_1
X_16841_ _06598_ _07263_ VGND VGND VPWR VPWR _07264_ sky130_fd_sc_hd__nor2_1
X_16772_ _07160_ _07161_ _07164_ _07188_ VGND VGND VPWR VPWR _07190_ sky130_fd_sc_hd__o211a_1
X_13984_ _03014_ _00399_ _04153_ _04156_ VGND VGND VPWR VPWR _04157_ sky130_fd_sc_hd__a22oi_1
X_18511_ _09075_ _09056_ _09077_ VGND VGND VPWR VPWR _09079_ sky130_fd_sc_hd__o21ai_1
X_15723_ _06048_ _06050_ VGND VGND VPWR VPWR _06053_ sky130_fd_sc_hd__and2_1
XFILLER_0_88_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12935_ _02505_ VGND VGND VPWR VPWR _03028_ sky130_fd_sc_hd__buf_4
XFILLER_0_87_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18442_ _08955_ _08958_ _09003_ VGND VGND VPWR VPWR _09006_ sky130_fd_sc_hd__and3_1
X_15654_ _05977_ VGND VGND VPWR VPWR _05978_ sky130_fd_sc_hd__inv_2
XTAP_2350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12866_ _01502_ _02891_ _02894_ _02940_ _02958_ VGND VGND VPWR VPWR _02959_ sky130_fd_sc_hd__o311ai_4
XTAP_2361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14605_ _02984_ _01520_ _07015_ _07962_ VGND VGND VPWR VPWR _04835_ sky130_fd_sc_hd__and4_1
XTAP_2383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11817_ _04362_ _00196_ _00871_ _04340_ VGND VGND VPWR VPWR _01910_ sky130_fd_sc_hd__a22oi_1
X_18373_ _01502_ _02888_ VGND VGND VPWR VPWR _08932_ sky130_fd_sc_hd__nor2_2
XTAP_2394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15585_ _05895_ _05902_ VGND VGND VPWR VPWR _05903_ sky130_fd_sc_hd__and2_1
XTAP_1660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12797_ _02889_ VGND VGND VPWR VPWR _02890_ sky130_fd_sc_hd__inv_2
XTAP_1682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17324_ _07701_ _07702_ _07789_ VGND VGND VPWR VPWR _07791_ sky130_fd_sc_hd__nand3_1
X_14536_ _00191_ _00460_ _05486_ _00189_ VGND VGND VPWR VPWR _04760_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_56_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11748_ _01836_ _01839_ _01828_ _01840_ VGND VGND VPWR VPWR _01841_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_153_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17255_ _06766_ _07387_ VGND VGND VPWR VPWR _07715_ sky130_fd_sc_hd__nor2_1
X_14467_ _04508_ _04510_ _04507_ VGND VGND VPWR VPWR _04685_ sky130_fd_sc_hd__o21ba_1
X_11679_ _01733_ _01734_ _01736_ VGND VGND VPWR VPWR _01772_ sky130_fd_sc_hd__nor3b_1
XFILLER_0_141_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16206_ net212 _03019_ _06517_ VGND VGND VPWR VPWR _06574_ sky130_fd_sc_hd__or3_1
X_13418_ _03537_ VGND VGND VPWR VPWR _03538_ sky130_fd_sc_hd__clkbuf_4
X_17186_ _07629_ _07639_ VGND VGND VPWR VPWR _07640_ sky130_fd_sc_hd__xnor2_1
X_14398_ _04461_ _04468_ _04606_ _04607_ VGND VGND VPWR VPWR _04609_ sky130_fd_sc_hd__a211o_4
XFILLER_0_12_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16137_ _01220_ _03134_ VGND VGND VPWR VPWR _06499_ sky130_fd_sc_hd__or2_1
X_13349_ _03460_ _03461_ VGND VGND VPWR VPWR _03462_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16068_ _06423_ VGND VGND VPWR VPWR _06424_ sky130_fd_sc_hd__buf_2
XFILLER_0_20_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15019_ _05285_ _05286_ VGND VGND VPWR VPWR _05287_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_45_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09511_ _04023_ _04176_ VGND VGND VPWR VPWR _04187_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_79_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18709_ _09237_ VGND VGND VPWR VPWR _00062_ sky130_fd_sc_hd__buf_1
XFILLER_0_79_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09442_ _03421_ VGND VGND VPWR VPWR _03432_ sky130_fd_sc_hd__clkbuf_8
XPHY_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_148_157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_145_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09709_ _06267_ _06319_ _06329_ VGND VGND VPWR VPWR _06340_ sky130_fd_sc_hd__nand3_2
X_10981_ _01061_ _01068_ _01072_ _01073_ VGND VGND VPWR VPWR _01074_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_69_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12720_ _02810_ _02812_ VGND VGND VPWR VPWR _02813_ sky130_fd_sc_hd__nor2_1
XFILLER_0_139_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12651_ _02735_ _02742_ _02743_ VGND VGND VPWR VPWR _02744_ sky130_fd_sc_hd__nand3_1
XFILLER_0_84_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11602_ _05856_ VGND VGND VPWR VPWR _01695_ sky130_fd_sc_hd__buf_4
X_15370_ _00591_ _05652_ _05667_ VGND VGND VPWR VPWR _05669_ sky130_fd_sc_hd__a21oi_1
X_12582_ _02638_ _02636_ _02637_ VGND VGND VPWR VPWR _02675_ sky130_fd_sc_hd__nand3_1
XFILLER_0_154_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_154_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14321_ _04512_ _04513_ _04524_ VGND VGND VPWR VPWR _04525_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_92_272 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11533_ _01622_ _01623_ _01624_ VGND VGND VPWR VPWR _01626_ sky130_fd_sc_hd__a21o_1
X_17040_ _00593_ _06463_ _07453_ _07480_ VGND VGND VPWR VPWR _07481_ sky130_fd_sc_hd__a22o_1
XFILLER_0_135_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14252_ _02188_ _09303_ _00498_ _04515_ VGND VGND VPWR VPWR _04450_ sky130_fd_sc_hd__a22oi_1
X_11464_ _01160_ _01161_ VGND VGND VPWR VPWR _01557_ sky130_fd_sc_hd__or2b_1
XFILLER_0_40_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_150_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10415_ _00506_ _00492_ _00493_ VGND VGND VPWR VPWR _00508_ sky130_fd_sc_hd__and3_1
X_13203_ _03302_ _03303_ VGND VGND VPWR VPWR _03304_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_151_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14183_ _04372_ _04374_ VGND VGND VPWR VPWR _04375_ sky130_fd_sc_hd__nand2_1
X_11395_ _01486_ _01487_ VGND VGND VPWR VPWR _01488_ sky130_fd_sc_hd__xor2_1
X_13134_ _04558_ _05715_ _03229_ _03230_ VGND VGND VPWR VPWR _03231_ sky130_fd_sc_hd__nand4_1
X_10346_ cla_inst.in1\[16\] VGND VGND VPWR VPWR _00439_ sky130_fd_sc_hd__clkbuf_4
X_18991_ clknet_4_6_0_clk _09357_ VGND VGND VPWR VPWR salida\[44\] sky130_fd_sc_hd__dfxtp_1
XTAP_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13065_ _07766_ _03156_ _03024_ VGND VGND VPWR VPWR _03157_ sky130_fd_sc_hd__o21ai_1
X_17942_ _08458_ _08462_ VGND VGND VPWR VPWR _08464_ sky130_fd_sc_hd__nand2_1
X_10277_ _08930_ _08984_ _00368_ _00369_ VGND VGND VPWR VPWR _00370_ sky130_fd_sc_hd__a211o_2
X_12016_ _01081_ _03388_ _00949_ _01082_ VGND VGND VPWR VPWR _02109_ sky130_fd_sc_hd__a22o_1
X_17873_ _08386_ _08388_ VGND VGND VPWR VPWR _08389_ sky130_fd_sc_hd__nor2_1
X_16824_ _07140_ _07141_ _07146_ VGND VGND VPWR VPWR _07246_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_45_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_cap2 _03204_ VGND VGND VPWR VPWR net320 sky130_fd_sc_hd__buf_1
X_16755_ _07168_ _07170_ VGND VGND VPWR VPWR _07171_ sky130_fd_sc_hd__xor2_1
X_13967_ _04136_ _04137_ VGND VGND VPWR VPWR _04138_ sky130_fd_sc_hd__xor2_1
XFILLER_0_45_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15706_ _06032_ _06033_ VGND VGND VPWR VPWR _06034_ sky130_fd_sc_hd__and2_1
X_12918_ _03010_ VGND VGND VPWR VPWR _03011_ sky130_fd_sc_hd__clkbuf_4
X_16686_ _07094_ _07095_ VGND VGND VPWR VPWR _07096_ sky130_fd_sc_hd__and2b_1
X_13898_ _03896_ _03895_ VGND VGND VPWR VPWR _04063_ sky130_fd_sc_hd__and2b_1
XFILLER_0_88_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18425_ _06024_ _06409_ _06407_ _06330_ VGND VGND VPWR VPWR _08988_ sky130_fd_sc_hd__o211a_1
XFILLER_0_119_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15637_ _03010_ _03012_ _03142_ _03055_ VGND VGND VPWR VPWR _05959_ sky130_fd_sc_hd__and4_1
XTAP_2180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12849_ _00592_ _00167_ _00228_ _00227_ VGND VGND VPWR VPWR _02942_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_75_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18356_ _08856_ _08859_ _08911_ VGND VGND VPWR VPWR _08913_ sky130_fd_sc_hd__or3_1
X_15568_ _07668_ _00119_ _01317_ _03009_ VGND VGND VPWR VPWR _05884_ sky130_fd_sc_hd__a22o_1
XTAP_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17307_ _07502_ _07640_ VGND VGND VPWR VPWR _07772_ sky130_fd_sc_hd__and2_1
X_14519_ _04598_ _04701_ _04739_ _04740_ VGND VGND VPWR VPWR _04741_ sky130_fd_sc_hd__a211o_4
X_18287_ _08835_ _08837_ _06836_ VGND VGND VPWR VPWR _08838_ sky130_fd_sc_hd__a21oi_1
X_15499_ _05685_ _05732_ VGND VGND VPWR VPWR _05809_ sky130_fd_sc_hd__and2b_1
XFILLER_0_4_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_136 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_127_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17238_ _00786_ _06369_ _06367_ VGND VGND VPWR VPWR _07697_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_9_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_153_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17169_ _00716_ _06889_ VGND VGND VPWR VPWR _07621_ sky130_fd_sc_hd__nand2_4
XFILLER_0_12_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09991_ _07711_ _09311_ _09263_ VGND VGND VPWR VPWR _09318_ sky130_fd_sc_hd__a21o_1
XFILLER_0_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09425_ _03184_ _03206_ _03228_ _03239_ VGND VGND VPWR VPWR _00002_ sky130_fd_sc_hd__a22o_1
XFILLER_0_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_149_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_902 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10200_ _04558_ _05257_ VGND VGND VPWR VPWR _00293_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_120_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11180_ _01238_ _01271_ _01272_ VGND VGND VPWR VPWR _01273_ sky130_fd_sc_hd__nor3_1
XFILLER_0_101_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_386 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10131_ _00190_ _00192_ _00223_ _00193_ _00186_ VGND VGND VPWR VPWR _00224_ sky130_fd_sc_hd__a41o_1
XFILLER_0_100_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10062_ _00153_ _00154_ VGND VGND VPWR VPWR _00155_ sky130_fd_sc_hd__and2_1
X_14870_ _03006_ _03107_ VGND VGND VPWR VPWR _05124_ sky130_fd_sc_hd__nand2_1
X_13821_ _03967_ _03977_ VGND VGND VPWR VPWR _03978_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_98_843 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16540_ _06749_ _06762_ _06893_ VGND VGND VPWR VPWR _06936_ sky130_fd_sc_hd__and3_1
X_13752_ _03738_ _03747_ _03902_ VGND VGND VPWR VPWR _03904_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_97_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10964_ _01054_ _01056_ VGND VGND VPWR VPWR _01057_ sky130_fd_sc_hd__and2_1
XFILLER_0_58_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12703_ _02769_ _02771_ VGND VGND VPWR VPWR _02796_ sky130_fd_sc_hd__nor2_1
X_16471_ _02826_ _02968_ _06861_ VGND VGND VPWR VPWR _06862_ sky130_fd_sc_hd__or3_1
X_13683_ _03642_ _03644_ _03827_ VGND VGND VPWR VPWR _03828_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_85_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10895_ _05224_ _08409_ _00986_ _00987_ VGND VGND VPWR VPWR _00988_ sky130_fd_sc_hd__a31o_1
X_18210_ _08753_ _08754_ _06836_ VGND VGND VPWR VPWR _08755_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_127_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15422_ _00115_ _09059_ VGND VGND VPWR VPWR _05726_ sky130_fd_sc_hd__nand2_1
XFILLER_0_54_902 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12634_ _02712_ _02726_ VGND VGND VPWR VPWR _02727_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_31_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_127_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18141_ _08675_ _08679_ _08677_ VGND VGND VPWR VPWR _08680_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_143_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15353_ _05646_ _05650_ VGND VGND VPWR VPWR _05651_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_25_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12565_ _02655_ _02657_ VGND VGND VPWR VPWR _02658_ sky130_fd_sc_hd__nor2_1
XFILLER_0_108_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14304_ _04494_ _04347_ _04506_ VGND VGND VPWR VPWR _04507_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_123_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11516_ _01556_ _01559_ _01519_ _01557_ VGND VGND VPWR VPWR _01609_ sky130_fd_sc_hd__a22o_1
XFILLER_0_80_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18072_ _06543_ _08599_ _08600_ _08604_ VGND VGND VPWR VPWR _08606_ sky130_fd_sc_hd__a31o_1
X_15284_ _03000_ _00339_ _05489_ VGND VGND VPWR VPWR _05576_ sky130_fd_sc_hd__nand3_1
XFILLER_0_41_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12496_ _02587_ _02588_ VGND VGND VPWR VPWR _02589_ sky130_fd_sc_hd__or2_2
XFILLER_0_34_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17023_ _07357_ _07360_ _07356_ VGND VGND VPWR VPWR _07463_ sky130_fd_sc_hd__a21boi_2
X_14235_ _03651_ _03662_ _06722_ _06689_ VGND VGND VPWR VPWR _04431_ sky130_fd_sc_hd__nand4_2
XFILLER_0_40_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11447_ _01526_ _01539_ VGND VGND VPWR VPWR _01540_ sky130_fd_sc_hd__nand2_2
XFILLER_0_111_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_528 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14166_ _04195_ _04206_ VGND VGND VPWR VPWR _04356_ sky130_fd_sc_hd__nand2_1
X_11378_ _00863_ _00864_ VGND VGND VPWR VPWR _01471_ sky130_fd_sc_hd__and2_1
X_13117_ _00604_ _00606_ _00605_ VGND VGND VPWR VPWR _03212_ sky130_fd_sc_hd__a21bo_1
XTAP_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10329_ _00418_ _00419_ _00420_ VGND VGND VPWR VPWR _00422_ sky130_fd_sc_hd__a21o_1
XTAP_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14097_ _02059_ _07025_ VGND VGND VPWR VPWR _04280_ sky130_fd_sc_hd__nand2_1
X_18974_ clknet_4_4_0_clk _09405_ VGND VGND VPWR VPWR salida\[27\] sky130_fd_sc_hd__dfxtp_1
XTAP_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17925_ _07256_ _08432_ _08433_ _08445_ VGND VGND VPWR VPWR _08446_ sky130_fd_sc_hd__a31o_1
X_13048_ _02505_ _06776_ VGND VGND VPWR VPWR _03140_ sky130_fd_sc_hd__nor2_1
X_17856_ _08368_ _08369_ VGND VGND VPWR VPWR _08370_ sky130_fd_sc_hd__nor2_1
X_16807_ _07224_ _07226_ VGND VGND VPWR VPWR _07227_ sky130_fd_sc_hd__xor2_1
X_17787_ _08188_ _08196_ VGND VGND VPWR VPWR _08295_ sky130_fd_sc_hd__or2b_1
X_14999_ _00191_ _00318_ _05758_ _00189_ VGND VGND VPWR VPWR _05265_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_49_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16738_ _07149_ _07151_ VGND VGND VPWR VPWR _07152_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_48_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16669_ _03790_ _06593_ _06594_ VGND VGND VPWR VPWR _07077_ sky130_fd_sc_hd__a21o_1
XFILLER_0_8_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18408_ _08967_ _08968_ VGND VGND VPWR VPWR _08969_ sky130_fd_sc_hd__and2b_1
XFILLER_0_118_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18339_ _08864_ _08866_ VGND VGND VPWR VPWR _08894_ sky130_fd_sc_hd__and2_1
XFILLER_0_154_480 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_331 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_130_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09974_ _09179_ VGND VGND VPWR VPWR _09188_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_0_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10680_ net169 _04220_ _00772_ net228 VGND VGND VPWR VPWR _00773_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_137_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12350_ _02376_ _02411_ _02442_ VGND VGND VPWR VPWR _02443_ sky130_fd_sc_hd__and3_2
XFILLER_0_50_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_105_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11301_ _01290_ _01379_ _01392_ _01393_ VGND VGND VPWR VPWR _01394_ sky130_fd_sc_hd__o211a_2
XFILLER_0_62_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12281_ _00846_ _00399_ _02373_ VGND VGND VPWR VPWR _02374_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_132_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14020_ _09353_ _00716_ _04033_ _04032_ VGND VGND VPWR VPWR _04196_ sky130_fd_sc_hd__a31o_1
X_11232_ _01086_ _01091_ VGND VGND VPWR VPWR _01325_ sky130_fd_sc_hd__or2b_1
XFILLER_0_31_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11163_ _00174_ _07548_ _07581_ cla_inst.in2\[24\] VGND VGND VPWR VPWR _01256_ sky130_fd_sc_hd__a22o_1
XFILLER_0_101_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10114_ _00206_ VGND VGND VPWR VPWR _00207_ sky130_fd_sc_hd__buf_4
X_11094_ _01056_ _01182_ _01186_ VGND VGND VPWR VPWR _01187_ sky130_fd_sc_hd__nand3_4
X_15971_ _06313_ _06315_ _06317_ _03124_ _06318_ VGND VGND VPWR VPWR _09376_ sky130_fd_sc_hd__a221o_1
X_17710_ _08208_ _08210_ VGND VGND VPWR VPWR _08211_ sky130_fd_sc_hd__xor2_1
X_14922_ _05140_ _05056_ _05179_ VGND VGND VPWR VPWR _05182_ sky130_fd_sc_hd__and3_1
X_10045_ _00124_ _00137_ VGND VGND VPWR VPWR _00138_ sky130_fd_sc_hd__xor2_1
X_18690_ net45 _03041_ _09193_ VGND VGND VPWR VPWR _09224_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold82 ApproximateM_inst.lob_16.lob1.mux.sel VGND VGND VPWR VPWR net245 sky130_fd_sc_hd__dlygate4sd3_1
X_17641_ _06382_ _06381_ _06380_ VGND VGND VPWR VPWR _08136_ sky130_fd_sc_hd__a21oi_1
X_14853_ _05103_ _05105_ VGND VGND VPWR VPWR _05106_ sky130_fd_sc_hd__or2_2
Xhold93 _00022_ VGND VGND VPWR VPWR net256 sky130_fd_sc_hd__dlygate4sd3_1
X_13804_ _03951_ _03959_ VGND VGND VPWR VPWR _03960_ sky130_fd_sc_hd__xnor2_1
X_17572_ _08058_ _08059_ VGND VGND VPWR VPWR _08061_ sky130_fd_sc_hd__nor2_1
X_14784_ _04913_ _04907_ VGND VGND VPWR VPWR _05031_ sky130_fd_sc_hd__and2b_1
XFILLER_0_86_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_98_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11996_ _02017_ _02020_ VGND VGND VPWR VPWR _02089_ sky130_fd_sc_hd__xnor2_1
X_16523_ _02974_ _06915_ _06918_ _06645_ VGND VGND VPWR VPWR _06919_ sky130_fd_sc_hd__a211o_1
X_13735_ _03834_ _03835_ _03882_ _03883_ VGND VGND VPWR VPWR _03885_ sky130_fd_sc_hd__o22a_1
XFILLER_0_129_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10947_ _04984_ _00206_ _01025_ _01024_ VGND VGND VPWR VPWR _01040_ sky130_fd_sc_hd__a31o_2
XFILLER_0_133_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16454_ _03060_ _06492_ VGND VGND VPWR VPWR _06844_ sky130_fd_sc_hd__nor2_1
X_13666_ _03786_ _03787_ _03807_ _03808_ VGND VGND VPWR VPWR _03809_ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_0_42_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10878_ _04438_ _04864_ _04143_ _04646_ VGND VGND VPWR VPWR _00971_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_128_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15405_ _05626_ _05628_ _05707_ VGND VGND VPWR VPWR _05708_ sky130_fd_sc_hd__and3_1
XFILLER_0_128_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12617_ _02694_ _02709_ VGND VGND VPWR VPWR _02710_ sky130_fd_sc_hd__xor2_1
X_16385_ _06757_ _06768_ VGND VGND VPWR VPWR _06769_ sky130_fd_sc_hd__nand2_1
XFILLER_0_53_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13597_ _00592_ _03108_ _03488_ VGND VGND VPWR VPWR _03734_ sky130_fd_sc_hd__and3_1
Xclkbuf_4_14_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_14_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_53_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18124_ _08660_ _08661_ VGND VGND VPWR VPWR _08662_ sky130_fd_sc_hd__or2_1
X_15336_ _05449_ _01139_ _05539_ _05538_ VGND VGND VPWR VPWR _05632_ sky130_fd_sc_hd__a31o_1
XFILLER_0_53_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12548_ _02597_ _02639_ _02640_ VGND VGND VPWR VPWR _02641_ sky130_fd_sc_hd__and3_1
X_18055_ _08413_ _08505_ VGND VGND VPWR VPWR _08587_ sky130_fd_sc_hd__or2b_1
X_15267_ _09353_ _00119_ VGND VGND VPWR VPWR _05557_ sky130_fd_sc_hd__nand2_2
XANTENNA_2 _00100_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12479_ _02566_ _02542_ VGND VGND VPWR VPWR _02572_ sky130_fd_sc_hd__and2b_1
XFILLER_0_112_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17006_ _07382_ _07383_ _07442_ VGND VGND VPWR VPWR _07444_ sky130_fd_sc_hd__and3_1
X_14218_ _03125_ _04257_ _04265_ _03199_ _04412_ VGND VGND VPWR VPWR _09383_ sky130_fd_sc_hd__a221o_1
XFILLER_0_10_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15198_ _00190_ _00192_ _07025_ _08876_ VGND VGND VPWR VPWR _05482_ sky130_fd_sc_hd__and4_1
XFILLER_0_111_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14149_ _01873_ _04336_ VGND VGND VPWR VPWR _04337_ sky130_fd_sc_hd__nand2_2
XTAP_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18957_ clknet_4_6_0_clk _09387_ VGND VGND VPWR VPWR salida\[10\] sky130_fd_sc_hd__dfxtp_1
XTAP_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17908_ _03368_ _06511_ _01692_ VGND VGND VPWR VPWR _08427_ sky130_fd_sc_hd__a21o_1
X_09690_ _05943_ _05954_ _06127_ VGND VGND VPWR VPWR _06138_ sky130_fd_sc_hd__nand3_4
X_18888_ clknet_4_12_0_clk _00042_ VGND VGND VPWR VPWR ApproximateM_inst.lob_16.lob1.genblk1\[6\].genblk1.mux.sel
+ sky130_fd_sc_hd__dfxtp_2
Xrebuffer14 _04683_ VGND VGND VPWR VPWR net177 sky130_fd_sc_hd__clkbuf_1
X_17839_ _07751_ _07489_ _07596_ _07039_ VGND VGND VPWR VPWR _08351_ sky130_fd_sc_hd__a22o_1
Xrebuffer25 _04599_ VGND VGND VPWR VPWR net188 sky130_fd_sc_hd__buf_1
XFILLER_0_89_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrebuffer36 _01859_ VGND VGND VPWR VPWR net199 sky130_fd_sc_hd__buf_1
Xrebuffer47 _01803_ VGND VGND VPWR VPWR net210 sky130_fd_sc_hd__clkbuf_1
Xrebuffer58 _05377_ VGND VGND VPWR VPWR net221 sky130_fd_sc_hd__buf_1
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer69 net233 VGND VGND VPWR VPWR net232 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_172 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09957_ _07341_ _07450_ VGND VGND VPWR VPWR _09037_ sky130_fd_sc_hd__nand2_1
XTAP_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09888_ _08126_ _08267_ _07919_ _07930_ VGND VGND VPWR VPWR _08289_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_99_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11850_ _01884_ _01942_ VGND VGND VPWR VPWR _01943_ sky130_fd_sc_hd__nand2_1
XTAP_2735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10801_ _00162_ _00230_ VGND VGND VPWR VPWR _00894_ sky130_fd_sc_hd__or2_1
XTAP_2768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11781_ _01873_ _01357_ _01680_ VGND VGND VPWR VPWR _01874_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_68_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13520_ _03408_ _03433_ _03647_ _03648_ VGND VGND VPWR VPWR _03649_ sky130_fd_sc_hd__a211oi_4
X_10732_ _08126_ _08137_ _08256_ VGND VGND VPWR VPWR _00825_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_12_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13451_ _03569_ _03572_ _03547_ VGND VGND VPWR VPWR _03573_ sky130_fd_sc_hd__mux2_1
X_10663_ _00754_ _00755_ VGND VGND VPWR VPWR _00756_ sky130_fd_sc_hd__or2_1
XFILLER_0_24_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12402_ _02492_ _02493_ _02494_ VGND VGND VPWR VPWR _02495_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_137_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16170_ _00181_ _06532_ _06533_ _06534_ _03313_ VGND VGND VPWR VPWR _06535_ sky130_fd_sc_hd__o32a_1
XFILLER_0_35_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13382_ _00112_ _03321_ _00165_ _00212_ VGND VGND VPWR VPWR _03499_ sky130_fd_sc_hd__and4_1
X_10594_ _00684_ _00686_ VGND VGND VPWR VPWR _00687_ sky130_fd_sc_hd__xor2_2
X_15121_ _05396_ _05397_ VGND VGND VPWR VPWR _05398_ sky130_fd_sc_hd__nand2_2
XFILLER_0_50_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12333_ _02423_ _02425_ VGND VGND VPWR VPWR _02426_ sky130_fd_sc_hd__nor2_1
XFILLER_0_121_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15052_ _05320_ _05321_ VGND VGND VPWR VPWR _05323_ sky130_fd_sc_hd__or2_1
XFILLER_0_133_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12264_ _06019_ _08039_ _00180_ _00130_ VGND VGND VPWR VPWR _02357_ sky130_fd_sc_hd__and4_1
XFILLER_0_31_470 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14003_ _04175_ _04177_ VGND VGND VPWR VPWR _04178_ sky130_fd_sc_hd__nor2_1
X_11215_ _01306_ _01307_ VGND VGND VPWR VPWR _01308_ sky130_fd_sc_hd__nand2_1
X_12195_ _02144_ _02145_ VGND VGND VPWR VPWR _02288_ sky130_fd_sc_hd__nand2_1
XFILLER_0_102_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput72 net72 VGND VGND VPWR VPWR leds[11] sky130_fd_sc_hd__buf_2
X_18811_ _09317_ VGND VGND VPWR VPWR _00094_ sky130_fd_sc_hd__clkbuf_1
X_11146_ _00253_ cla_inst.in2\[21\] _07570_ _07613_ VGND VGND VPWR VPWR _01239_ sky130_fd_sc_hd__and4_1
Xoutput83 net83 VGND VGND VPWR VPWR o_wb_data[0] sky130_fd_sc_hd__clkbuf_4
Xoutput94 net94 VGND VGND VPWR VPWR o_wb_data[1] sky130_fd_sc_hd__clkbuf_4
X_11077_ _01168_ _01169_ VGND VGND VPWR VPWR _01170_ sky130_fd_sc_hd__xnor2_2
X_18742_ _03036_ net62 _09251_ VGND VGND VPWR VPWR _09264_ sky130_fd_sc_hd__mux2_1
X_15954_ _06300_ VGND VGND VPWR VPWR _06301_ sky130_fd_sc_hd__inv_2
X_14905_ _00190_ _05986_ _05162_ VGND VGND VPWR VPWR _05163_ sky130_fd_sc_hd__a21oi_1
X_10028_ _00120_ _08158_ VGND VGND VPWR VPWR _00121_ sky130_fd_sc_hd__and2_4
X_18673_ _09209_ _09213_ VGND VGND VPWR VPWR _09214_ sky130_fd_sc_hd__and2_1
X_15885_ _06192_ _06226_ _02969_ VGND VGND VPWR VPWR _06228_ sky130_fd_sc_hd__a21o_1
X_17624_ _08116_ _08117_ VGND VGND VPWR VPWR _08118_ sky130_fd_sc_hd__nor2_1
X_14836_ _03051_ _03114_ _02981_ VGND VGND VPWR VPWR _05088_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17555_ _08011_ _08012_ VGND VGND VPWR VPWR _08042_ sky130_fd_sc_hd__nor2_1
XFILLER_0_98_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14767_ _04999_ _05000_ _05011_ VGND VGND VPWR VPWR _05012_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_86_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11979_ _01973_ _01974_ _01975_ _01944_ VGND VGND VPWR VPWR _02072_ sky130_fd_sc_hd__o22a_1
X_16506_ _06826_ _06899_ VGND VGND VPWR VPWR _06900_ sky130_fd_sc_hd__xor2_2
X_13718_ cla_inst.in2\[27\] cla_inst.in2\[26\] _03837_ _03410_ VGND VGND VPWR VPWR
+ _03866_ sky130_fd_sc_hd__and4_1
XFILLER_0_85_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17486_ _07840_ _07849_ _07966_ VGND VGND VPWR VPWR _07967_ sky130_fd_sc_hd__a21oi_1
X_14698_ _04807_ _04808_ _04805_ VGND VGND VPWR VPWR _04937_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_128_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16437_ _06657_ _06749_ _06763_ VGND VGND VPWR VPWR _06825_ sky130_fd_sc_hd__a21o_1
X_13649_ _06040_ VGND VGND VPWR VPWR _03790_ sky130_fd_sc_hd__buf_4
XFILLER_0_144_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_116_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16368_ _06749_ VGND VGND VPWR VPWR _06750_ sky130_fd_sc_hd__buf_4
XFILLER_0_5_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18107_ _07106_ _07861_ _08642_ _08639_ VGND VGND VPWR VPWR _08643_ sky130_fd_sc_hd__o22a_1
X_15319_ _05612_ _05613_ VGND VGND VPWR VPWR _05614_ sky130_fd_sc_hd__nand2_2
XFILLER_0_5_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_152_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16299_ _06513_ _06587_ _06586_ VGND VGND VPWR VPWR _06675_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_75_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18038_ _08477_ _08566_ _08567_ VGND VGND VPWR VPWR _08568_ sky130_fd_sc_hd__a21o_1
XFILLER_0_112_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09811_ _07395_ _07439_ VGND VGND VPWR VPWR _07450_ sky130_fd_sc_hd__xnor2_2
X_09742_ _05649_ _05704_ _06689_ _06029_ VGND VGND VPWR VPWR _06700_ sky130_fd_sc_hd__a22o_1
XFILLER_0_94_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09673_ _05529_ _05867_ _05932_ VGND VGND VPWR VPWR _05954_ sky130_fd_sc_hd__a21o_1
XTAP_2009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11000_ _01085_ _01092_ VGND VGND VPWR VPWR _01093_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_99_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12951_ _01223_ VGND VGND VPWR VPWR _03044_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_88_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11902_ _01992_ _01994_ VGND VGND VPWR VPWR _01995_ sky130_fd_sc_hd__or2_1
X_15670_ _05920_ _05993_ VGND VGND VPWR VPWR _05995_ sky130_fd_sc_hd__or2_1
XFILLER_0_87_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12882_ _02974_ VGND VGND VPWR VPWR _02975_ sky130_fd_sc_hd__buf_4
XTAP_2521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14621_ _04849_ _04850_ _04851_ VGND VGND VPWR VPWR _04852_ sky130_fd_sc_hd__and3_1
XTAP_2543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11833_ _01920_ _01921_ _01925_ VGND VGND VPWR VPWR _01926_ sky130_fd_sc_hd__nor3b_2
XTAP_2554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17340_ _06368_ _06438_ _03311_ VGND VGND VPWR VPWR _07808_ sky130_fd_sc_hd__a21oi_1
XTAP_2587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14552_ _04654_ _04660_ VGND VGND VPWR VPWR _04778_ sky130_fd_sc_hd__and2b_1
XTAP_1853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11764_ _01852_ _01855_ VGND VGND VPWR VPWR _01857_ sky130_fd_sc_hd__and2_1
XTAP_1864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13503_ _03418_ VGND VGND VPWR VPWR _03631_ sky130_fd_sc_hd__inv_2
XTAP_1886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17271_ _07729_ _07730_ VGND VGND VPWR VPWR _07732_ sky130_fd_sc_hd__nand2_1
X_10715_ _00806_ _06591_ _04569_ _04449_ VGND VGND VPWR VPWR _00808_ sky130_fd_sc_hd__and4_1
XTAP_1897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14483_ _04587_ _04593_ VGND VGND VPWR VPWR _04702_ sky130_fd_sc_hd__nand2_1
XFILLER_0_153_512 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11695_ _01748_ _01778_ VGND VGND VPWR VPWR _01788_ sky130_fd_sc_hd__and2b_1
X_19010_ clknet_4_1_0_clk _09378_ VGND VGND VPWR VPWR salida\[63\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16222_ _06547_ VGND VGND VPWR VPWR _06592_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_125_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13434_ _03551_ _03555_ _02780_ VGND VGND VPWR VPWR _03556_ sky130_fd_sc_hd__mux2_1
X_10646_ _00718_ _00737_ _00738_ VGND VGND VPWR VPWR _00739_ sky130_fd_sc_hd__or3_2
XFILLER_0_153_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16153_ _03771_ ApproximateM_inst.lob_16.lob2.genblk1\[14\].genblk1.mux.sel _03184_
+ VGND VGND VPWR VPWR _06517_ sky130_fd_sc_hd__or3b_2
Xrebuffer5 _06541_ VGND VGND VPWR VPWR net168 sky130_fd_sc_hd__buf_1
XFILLER_0_141_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13365_ _03478_ _03479_ VGND VGND VPWR VPWR _03480_ sky130_fd_sc_hd__xor2_1
X_10577_ _07363_ _00509_ _00668_ _00669_ VGND VGND VPWR VPWR _00670_ sky130_fd_sc_hd__nand4_1
XFILLER_0_134_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_140_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15104_ _05378_ _05379_ VGND VGND VPWR VPWR _05380_ sky130_fd_sc_hd__xnor2_1
X_12316_ _02360_ _02406_ _02408_ VGND VGND VPWR VPWR _02409_ sky130_fd_sc_hd__or3_1
XFILLER_0_23_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16084_ _03111_ _03693_ _06441_ VGND VGND VPWR VPWR _06442_ sky130_fd_sc_hd__and3_1
X_13296_ _03402_ _03403_ VGND VGND VPWR VPWR _03404_ sky130_fd_sc_hd__and2b_1
XFILLER_0_139_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15035_ _05302_ _05303_ _04823_ VGND VGND VPWR VPWR _05305_ sky130_fd_sc_hd__o21ai_1
X_12247_ _02208_ _02331_ VGND VGND VPWR VPWR _02340_ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_121_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12178_ _02128_ _02258_ VGND VGND VPWR VPWR _02271_ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11129_ _01137_ _01221_ VGND VGND VPWR VPWR _01222_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16986_ _07304_ _07306_ _07301_ VGND VGND VPWR VPWR _07422_ sky130_fd_sc_hd__o21ba_1
X_18725_ _09110_ _09115_ _09178_ VGND VGND VPWR VPWR _09250_ sky130_fd_sc_hd__nor3_4
X_15937_ _06242_ _06254_ _06281_ VGND VGND VPWR VPWR _06283_ sky130_fd_sc_hd__and3_1
X_15868_ _06207_ _06208_ VGND VGND VPWR VPWR _06209_ sky130_fd_sc_hd__nand2_1
X_18656_ _09200_ VGND VGND VPWR VPWR _00041_ sky130_fd_sc_hd__buf_1
XFILLER_0_78_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17607_ _08083_ _08098_ VGND VGND VPWR VPWR _08099_ sky130_fd_sc_hd__xnor2_1
X_14819_ _04932_ _04964_ _05067_ _05068_ VGND VGND VPWR VPWR _05069_ sky130_fd_sc_hd__o211ai_4
X_15799_ _06134_ VGND VGND VPWR VPWR _06135_ sky130_fd_sc_hd__inv_2
XFILLER_0_80_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18587_ salida\[13\] _09141_ _09142_ salida\[45\] _09146_ VGND VGND VPWR VPWR _09149_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_148_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17538_ _03693_ _07355_ _02989_ VGND VGND VPWR VPWR _08024_ sky130_fd_sc_hd__or3b_1
XFILLER_0_47_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17469_ _07945_ _07946_ VGND VGND VPWR VPWR _07948_ sky130_fd_sc_hd__and2_1
XFILLER_0_15_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_707 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_735 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09725_ _06340_ _06351_ _06362_ VGND VGND VPWR VPWR _06515_ sky130_fd_sc_hd__a21o_1
X_09656_ _05627_ VGND VGND VPWR VPWR _05769_ sky130_fd_sc_hd__inv_2
XTAP_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09587_ ApproximateM_inst.lob_16.lob2.genblk1\[11\].genblk1.mux.sel VGND VGND VPWR
+ VPWR _05017_ sky130_fd_sc_hd__buf_4
XTAP_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_443 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_135_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_540 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_107_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_523 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10500_ _00399_ VGND VGND VPWR VPWR _00593_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_107_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11480_ _01568_ _01569_ _01572_ VGND VGND VPWR VPWR _01573_ sky130_fd_sc_hd__nand3_1
XFILLER_0_135_578 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_150_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10431_ _00519_ _00523_ VGND VGND VPWR VPWR _00524_ sky130_fd_sc_hd__nand2_1
XFILLER_0_123_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13150_ _00644_ _00645_ _07134_ _00309_ VGND VGND VPWR VPWR _03248_ sky130_fd_sc_hd__and4_1
X_10362_ _04690_ _08757_ _00451_ _00452_ VGND VGND VPWR VPWR _00455_ sky130_fd_sc_hd__a22o_1
X_12101_ _02098_ _02101_ VGND VGND VPWR VPWR _02194_ sky130_fd_sc_hd__xnor2_1
X_10293_ _09197_ _09226_ VGND VGND VPWR VPWR _00386_ sky130_fd_sc_hd__nor2_1
X_13081_ _03025_ _03094_ VGND VGND VPWR VPWR _03173_ sky130_fd_sc_hd__and2_1
X_12032_ _00514_ _02044_ VGND VGND VPWR VPWR _02125_ sky130_fd_sc_hd__nor2_2
X_16840_ _06358_ _06357_ _06356_ VGND VGND VPWR VPWR _07263_ sky130_fd_sc_hd__o21a_1
X_16771_ _06508_ _07171_ _07187_ VGND VGND VPWR VPWR _07188_ sky130_fd_sc_hd__a21oi_1
X_13983_ net218 VGND VGND VPWR VPWR _04156_ sky130_fd_sc_hd__inv_2
X_15722_ _06048_ _06050_ VGND VGND VPWR VPWR _06052_ sky130_fd_sc_hd__nor2_1
X_18510_ _09075_ _09056_ _09077_ VGND VGND VPWR VPWR _09078_ sky130_fd_sc_hd__or3_1
X_12934_ _03026_ VGND VGND VPWR VPWR _03027_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_34_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15653_ _00115_ _00665_ _05974_ _05976_ VGND VGND VPWR VPWR _05977_ sky130_fd_sc_hd__and4_1
X_18441_ _08955_ _08958_ _09003_ VGND VGND VPWR VPWR _09004_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_34_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12865_ _02957_ VGND VGND VPWR VPWR _02958_ sky130_fd_sc_hd__inv_2
XTAP_2340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14604_ _04723_ _04724_ _04734_ VGND VGND VPWR VPWR _04834_ sky130_fd_sc_hd__nor3_2
XTAP_2373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18372_ _08927_ _08928_ VGND VGND VPWR VPWR _08931_ sky130_fd_sc_hd__nand2_1
X_11816_ _04493_ _04416_ _00129_ ApproximateM_inst.lob_16.lob1.genblk1\[2\].genblk1.mux.sel
+ VGND VGND VPWR VPWR _01909_ sky130_fd_sc_hd__and4_1
XTAP_2384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15584_ _05900_ _05901_ VGND VGND VPWR VPWR _05902_ sky130_fd_sc_hd__xnor2_1
XTAP_1650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_410 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12796_ _02887_ _01502_ _02888_ VGND VGND VPWR VPWR _02889_ sky130_fd_sc_hd__or3_4
XTAP_2395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17323_ _07701_ _07702_ _07789_ VGND VGND VPWR VPWR _07790_ sky130_fd_sc_hd__a21oi_1
X_14535_ _04754_ _04757_ _04609_ _04699_ VGND VGND VPWR VPWR _04759_ sky130_fd_sc_hd__o211ai_2
XTAP_1683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11747_ _01820_ _01826_ _01827_ VGND VGND VPWR VPWR _01840_ sky130_fd_sc_hd__nand3_2
XFILLER_0_139_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17254_ _07712_ _07713_ VGND VGND VPWR VPWR _07714_ sky130_fd_sc_hd__nor2_1
X_14466_ _04681_ _04682_ _04564_ _04565_ VGND VGND VPWR VPWR _04684_ sky130_fd_sc_hd__o211a_2
XFILLER_0_50_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11678_ _01721_ _01739_ net198 _01770_ VGND VGND VPWR VPWR _01771_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_126_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16205_ _06084_ _06711_ _06524_ VGND VGND VPWR VPWR _06573_ sky130_fd_sc_hd__or3_1
XFILLER_0_52_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13417_ _03536_ VGND VGND VPWR VPWR _03537_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_153_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10629_ _00544_ _00551_ VGND VGND VPWR VPWR _00722_ sky130_fd_sc_hd__nand2_1
X_17185_ _07637_ _07638_ VGND VGND VPWR VPWR _07639_ sky130_fd_sc_hd__xor2_1
X_14397_ _04606_ _04607_ _04461_ _04468_ VGND VGND VPWR VPWR _04608_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_52_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16136_ _02983_ _06495_ _06497_ _06467_ VGND VGND VPWR VPWR _06498_ sky130_fd_sc_hd__o211a_1
X_13348_ _03450_ _03451_ _03459_ VGND VGND VPWR VPWR _03461_ sky130_fd_sc_hd__and3_1
XFILLER_0_12_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16067_ _06418_ _06422_ VGND VGND VPWR VPWR _06423_ sky130_fd_sc_hd__or2_1
X_13279_ _03892_ _06613_ _08049_ _03881_ VGND VGND VPWR VPWR _03385_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15018_ _05161_ _05178_ _05158_ VGND VGND VPWR VPWR _05286_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_20_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16969_ _07288_ _07291_ _07402_ VGND VGND VPWR VPWR _07403_ sky130_fd_sc_hd__a21o_1
X_09510_ _04110_ _04165_ VGND VGND VPWR VPWR _04176_ sky130_fd_sc_hd__nor2_2
X_18708_ _09209_ _09236_ VGND VGND VPWR VPWR _09237_ sky130_fd_sc_hd__and2_1
X_09441_ ApproximateM_inst.lob_16.lob1.genblk1\[8\].genblk1.mux.sel VGND VGND VPWR
+ VPWR _03421_ sky130_fd_sc_hd__buf_6
X_18639_ net46 _01746_ _09183_ VGND VGND VPWR VPWR _09186_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_145_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_144_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_762 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09708_ _06234_ _06245_ _06256_ VGND VGND VPWR VPWR _06329_ sky130_fd_sc_hd__a21o_1
X_10980_ _01069_ _01070_ _01071_ VGND VGND VPWR VPWR _01073_ sky130_fd_sc_hd__nand3_1
XFILLER_0_97_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09639_ ApproximateM_inst.lob_16.lob2.genblk1\[6\].genblk1.mux.sel VGND VGND VPWR
+ VPWR _05584_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_69_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12650_ _02740_ _02741_ _02733_ _02739_ VGND VGND VPWR VPWR _02743_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_77_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11601_ _01693_ _01673_ VGND VGND VPWR VPWR _01694_ sky130_fd_sc_hd__and2b_1
X_12581_ _02597_ _02639_ _02640_ VGND VGND VPWR VPWR _02674_ sky130_fd_sc_hd__nand3_1
XFILLER_0_53_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14320_ _04325_ _04523_ VGND VGND VPWR VPWR _04524_ sky130_fd_sc_hd__xor2_1
XFILLER_0_80_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11532_ _01622_ _01623_ _01624_ VGND VGND VPWR VPWR _01625_ sky130_fd_sc_hd__nand3_2
XFILLER_0_93_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_284 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14251_ _02059_ _07025_ _04278_ _04277_ _08876_ VGND VGND VPWR VPWR _04448_ sky130_fd_sc_hd__a32o_1
X_11463_ _01552_ _01555_ VGND VGND VPWR VPWR _01556_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_33_340 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13202_ _01505_ _00399_ _00705_ _00704_ VGND VGND VPWR VPWR _03303_ sky130_fd_sc_hd__a31o_1
X_10414_ _00492_ _00493_ _00506_ VGND VGND VPWR VPWR _00507_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_33_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14182_ _04357_ _04358_ _04371_ VGND VGND VPWR VPWR _04374_ sky130_fd_sc_hd__or3_1
X_11394_ _01358_ _01420_ _01434_ VGND VGND VPWR VPWR _01487_ sky130_fd_sc_hd__a21o_1
XFILLER_0_60_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13133_ _04646_ _04373_ _05606_ _05617_ VGND VGND VPWR VPWR _03230_ sky130_fd_sc_hd__nand4_2
X_10345_ _00435_ _00436_ _00437_ VGND VGND VPWR VPWR _00438_ sky130_fd_sc_hd__nand3_1
X_18990_ clknet_4_3_0_clk _09356_ VGND VGND VPWR VPWR salida\[43\] sky130_fd_sc_hd__dfxtp_1
XTAP_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13064_ _03026_ _03155_ VGND VGND VPWR VPWR _03156_ sky130_fd_sc_hd__and2_1
X_17941_ _08459_ _08461_ VGND VGND VPWR VPWR _08462_ sky130_fd_sc_hd__xnor2_1
X_10276_ _00349_ _00350_ _00367_ VGND VGND VPWR VPWR _00369_ sky130_fd_sc_hd__and3_1
X_12015_ _02031_ _02039_ VGND VGND VPWR VPWR _02108_ sky130_fd_sc_hd__xnor2_1
X_17872_ _07630_ _07861_ _08385_ VGND VGND VPWR VPWR _08388_ sky130_fd_sc_hd__o21a_1
X_16823_ _07240_ _07244_ VGND VGND VPWR VPWR _07245_ sky130_fd_sc_hd__xor2_1
XFILLER_0_136_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_49 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13966_ _03970_ _03973_ _03971_ VGND VGND VPWR VPWR _04137_ sky130_fd_sc_hd__o21ba_1
X_16754_ _06990_ _06991_ _07096_ _07169_ VGND VGND VPWR VPWR _07170_ sky130_fd_sc_hd__a31o_1
Xmax_cap3 _03884_ VGND VGND VPWR VPWR net321 sky130_fd_sc_hd__clkbuf_1
X_12917_ _03009_ VGND VGND VPWR VPWR _03010_ sky130_fd_sc_hd__buf_2
X_15705_ _03007_ _03055_ _06031_ VGND VGND VPWR VPWR _06033_ sky130_fd_sc_hd__a21o_1
X_16685_ _00881_ _06673_ _03790_ VGND VGND VPWR VPWR _07095_ sky130_fd_sc_hd__or3b_1
X_13897_ _04060_ _04061_ VGND VGND VPWR VPWR _04062_ sky130_fd_sc_hd__xor2_1
XFILLER_0_152_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18424_ _02920_ net115 _08986_ VGND VGND VPWR VPWR _08987_ sky130_fd_sc_hd__a21o_1
X_12848_ _02928_ _02929_ _02931_ VGND VGND VPWR VPWR _02941_ sky130_fd_sc_hd__and3_1
X_15636_ _03007_ _04900_ VGND VGND VPWR VPWR _05958_ sky130_fd_sc_hd__nand2_1
XTAP_2170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15567_ _03009_ _07668_ _00119_ _01317_ VGND VGND VPWR VPWR _05883_ sky130_fd_sc_hd__and4_1
XFILLER_0_61_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18355_ _08856_ _08859_ _08911_ VGND VGND VPWR VPWR _08912_ sky130_fd_sc_hd__o21ai_1
XTAP_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12779_ _02853_ _02865_ VGND VGND VPWR VPWR _02872_ sky130_fd_sc_hd__nand2_1
XFILLER_0_127_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14518_ _04737_ _04738_ _04702_ _04703_ VGND VGND VPWR VPWR _04740_ sky130_fd_sc_hd__o211a_1
XFILLER_0_124_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17306_ _07769_ _07770_ VGND VGND VPWR VPWR _07771_ sky130_fd_sc_hd__xnor2_1
X_15498_ _05773_ _05757_ _05759_ VGND VGND VPWR VPWR _05808_ sky130_fd_sc_hd__nand3_1
X_18286_ _08753_ _08754_ _08815_ _08836_ VGND VGND VPWR VPWR _08837_ sky130_fd_sc_hd__a31o_1
XFILLER_0_127_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_154_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_142_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14449_ _04651_ _04652_ _04663_ VGND VGND VPWR VPWR _04665_ sky130_fd_sc_hd__or3_1
X_17237_ _03198_ _05086_ _07693_ _07695_ VGND VGND VPWR VPWR _07696_ sky130_fd_sc_hd__a211o_1
XFILLER_0_141_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17168_ _07518_ _07528_ _07525_ VGND VGND VPWR VPWR _07620_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_141_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16119_ _06470_ _06478_ _03077_ VGND VGND VPWR VPWR _06479_ sky130_fd_sc_hd__a21o_1
X_09990_ _09303_ VGND VGND VPWR VPWR _09311_ sky130_fd_sc_hd__buf_4
X_17099_ _07543_ _07544_ VGND VGND VPWR VPWR _07545_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_86_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09424_ op_code\[0\] VGND VGND VPWR VPWR _03239_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_137_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_149_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_638 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_117_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10130_ _00194_ VGND VGND VPWR VPWR _00223_ sky130_fd_sc_hd__buf_4
XFILLER_0_30_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10061_ _00106_ _00147_ _00150_ _00152_ VGND VGND VPWR VPWR _00154_ sky130_fd_sc_hd__a22o_1
XFILLER_0_100_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13820_ _03969_ _03976_ VGND VGND VPWR VPWR _03977_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_98_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_855 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13751_ _03900_ _03901_ VGND VGND VPWR VPWR _03902_ sky130_fd_sc_hd__xnor2_2
X_10963_ _05213_ _04657_ _01054_ _01055_ VGND VGND VPWR VPWR _01056_ sky130_fd_sc_hd__nand4_4
X_12702_ _02758_ _02791_ _02794_ VGND VGND VPWR VPWR _02795_ sky130_fd_sc_hd__a21oi_2
X_16470_ _02823_ _02825_ VGND VGND VPWR VPWR _06861_ sky130_fd_sc_hd__nor2_1
X_13682_ _03816_ _03825_ VGND VGND VPWR VPWR _03827_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_38_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10894_ ApproximateM_inst.lob_16.lob2.genblk1\[10\].genblk1.mux.sel _05290_ ApproximateM_inst.lob_16.lob1.genblk1\[13\].genblk1.mux.sel
+ ApproximateM_inst.lob_16.lob1.genblk1\[12\].genblk1.mux.sel VGND VGND VPWR VPWR
+ _00987_ sky130_fd_sc_hd__and4_1
XFILLER_0_97_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15421_ _05722_ _05723_ VGND VGND VPWR VPWR _05724_ sky130_fd_sc_hd__nor2_1
X_12633_ _02716_ _02718_ _02719_ _02725_ VGND VGND VPWR VPWR _02726_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_26_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15352_ _05647_ _05648_ VGND VGND VPWR VPWR _05650_ sky130_fd_sc_hd__or2_1
X_18140_ _08676_ VGND VGND VPWR VPWR _08679_ sky130_fd_sc_hd__inv_2
X_12564_ _02611_ _02654_ VGND VGND VPWR VPWR _02657_ sky130_fd_sc_hd__and2_1
XFILLER_0_109_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14303_ _04503_ _04505_ VGND VGND VPWR VPWR _04506_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_124_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_136_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11515_ _01164_ _01163_ _01156_ VGND VGND VPWR VPWR _01608_ sky130_fd_sc_hd__a21o_1
X_18071_ _06462_ _08602_ _08603_ VGND VGND VPWR VPWR _08604_ sky130_fd_sc_hd__or3_1
Xwire131 _03265_ VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__buf_2
X_15283_ _05370_ _05487_ _05485_ VGND VGND VPWR VPWR _05575_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_25_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire142 _00850_ VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__buf_1
X_12495_ _02584_ _02586_ VGND VGND VPWR VPWR _02588_ sky130_fd_sc_hd__nor2_1
X_17022_ _08615_ _07459_ _07460_ VGND VGND VPWR VPWR _07462_ sky130_fd_sc_hd__a21o_1
XFILLER_0_22_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14234_ _03596_ _06722_ _05606_ _03629_ VGND VGND VPWR VPWR _04430_ sky130_fd_sc_hd__a22o_1
XFILLER_0_123_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11446_ _01535_ _01538_ VGND VGND VPWR VPWR _01539_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_80_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14165_ _03993_ _04205_ VGND VGND VPWR VPWR _04355_ sky130_fd_sc_hd__or2_1
X_11377_ _01315_ _01419_ VGND VGND VPWR VPWR _01470_ sky130_fd_sc_hd__and2_1
X_13116_ _03207_ _03208_ _03209_ VGND VGND VPWR VPWR _03211_ sky130_fd_sc_hd__a21o_1
XTAP_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10328_ _00418_ _00419_ _00420_ VGND VGND VPWR VPWR _00421_ sky130_fd_sc_hd__nand3_2
XTAP_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14096_ _07123_ _04277_ _04278_ VGND VGND VPWR VPWR _04279_ sky130_fd_sc_hd__a21bo_1
X_18973_ clknet_4_5_0_clk _09404_ VGND VGND VPWR VPWR salida\[26\] sky130_fd_sc_hd__dfxtp_1
XTAP_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17924_ _08444_ VGND VGND VPWR VPWR _08445_ sky130_fd_sc_hd__inv_2
X_13047_ _03138_ VGND VGND VPWR VPWR _03139_ sky130_fd_sc_hd__inv_2
X_10259_ _07799_ cla_inst.in1\[31\] _09256_ ApproximateM_inst.lob_16.lob2.genblk1\[1\].genblk1.mux.sel
+ VGND VGND VPWR VPWR _00352_ sky130_fd_sc_hd__a22o_1
X_17855_ _07394_ _07604_ _07665_ _07649_ VGND VGND VPWR VPWR _08369_ sky130_fd_sc_hd__and4_1
X_16806_ _07122_ _07132_ _07225_ VGND VGND VPWR VPWR _07226_ sky130_fd_sc_hd__a21o_1
X_17786_ _08292_ _08293_ VGND VGND VPWR VPWR _08294_ sky130_fd_sc_hd__or2_1
X_14998_ _05163_ _05166_ _05164_ VGND VGND VPWR VPWR _05264_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_88_332 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16737_ _07049_ _07057_ _07150_ VGND VGND VPWR VPWR _07151_ sky130_fd_sc_hd__a21o_1
X_13949_ _03954_ _03955_ _04116_ VGND VGND VPWR VPWR _04118_ sky130_fd_sc_hd__nor3_1
XFILLER_0_88_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_218 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_410 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16668_ _00881_ _06433_ VGND VGND VPWR VPWR _07076_ sky130_fd_sc_hd__nor2_1
X_18407_ _08868_ _08917_ VGND VGND VPWR VPWR _08968_ sky130_fd_sc_hd__and2_1
X_15619_ _05938_ _05939_ VGND VGND VPWR VPWR _05940_ sky130_fd_sc_hd__and2_1
XFILLER_0_29_465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16599_ _07000_ VGND VGND VPWR VPWR _07001_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18338_ _08807_ _08870_ VGND VGND VPWR VPWR _08893_ sky130_fd_sc_hd__nor2_1
XFILLER_0_16_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_802 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_127_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18269_ _02869_ _08760_ VGND VGND VPWR VPWR _08819_ sky130_fd_sc_hd__nand2_2
XFILLER_0_154_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_298 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_130_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_141_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09973_ ApproximateM_inst.lob_16.lob1.genblk1\[1\].genblk1.mux.sel VGND VGND VPWR
+ VPWR _09179_ sky130_fd_sc_hd__buf_4
XFILLER_0_79_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11300_ _01389_ _01390_ _01391_ _01382_ VGND VGND VPWR VPWR _01393_ sky130_fd_sc_hd__a22o_1
XFILLER_0_50_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_596 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_132_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12280_ _01113_ _02259_ VGND VGND VPWR VPWR _02373_ sky130_fd_sc_hd__nor2_2
XFILLER_0_62_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11231_ _01319_ _01323_ VGND VGND VPWR VPWR _01324_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_105_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11162_ cla_inst.in2\[24\] _00174_ _07548_ _07581_ VGND VGND VPWR VPWR _01255_ sky130_fd_sc_hd__nand4_1
X_10113_ _00205_ VGND VGND VPWR VPWR _00206_ sky130_fd_sc_hd__clkbuf_8
X_11093_ _01183_ _01184_ _01185_ VGND VGND VPWR VPWR _01186_ sky130_fd_sc_hd__a21bo_1
X_15970_ _04241_ _04079_ _05623_ VGND VGND VPWR VPWR _06318_ sky130_fd_sc_hd__and3_1
X_14921_ _05140_ _05056_ _05179_ VGND VGND VPWR VPWR _05180_ sky130_fd_sc_hd__a21oi_2
X_10044_ _00133_ _00136_ VGND VGND VPWR VPWR _00137_ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17640_ _08132_ _08133_ _08134_ VGND VGND VPWR VPWR _08135_ sky130_fd_sc_hd__o21ai_1
X_14852_ _01521_ _00498_ _05101_ _05102_ VGND VGND VPWR VPWR _05105_ sky130_fd_sc_hd__and4_1
Xhold83 ApproximateM_inst.lob_16.lob1.genblk1\[3\].genblk1.mux.sel VGND VGND VPWR
+ VPWR net246 sky130_fd_sc_hd__dlygate4sd3_1
Xhold94 net96 VGND VGND VPWR VPWR net257 sky130_fd_sc_hd__dlygate4sd3_1
X_13803_ _03952_ _03958_ VGND VGND VPWR VPWR _03959_ sky130_fd_sc_hd__xor2_1
X_14783_ _04877_ _05029_ VGND VGND VPWR VPWR _05030_ sky130_fd_sc_hd__xnor2_1
X_17571_ _07143_ _07387_ _08055_ _08057_ VGND VGND VPWR VPWR _08059_ sky130_fd_sc_hd__o22a_1
X_11995_ _02083_ _02087_ VGND VGND VPWR VPWR _02088_ sky130_fd_sc_hd__or2_1
X_13734_ _03834_ _03835_ _03882_ _03883_ VGND VGND VPWR VPWR _03884_ sky130_fd_sc_hd__nor4_1
X_16522_ _02974_ _06916_ VGND VGND VPWR VPWR _06918_ sky130_fd_sc_hd__nor2_1
X_10946_ _01022_ _01023_ _01038_ VGND VGND VPWR VPWR _01039_ sky130_fd_sc_hd__and3_4
XFILLER_0_85_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13665_ _03805_ _03806_ _03788_ VGND VGND VPWR VPWR _03808_ sky130_fd_sc_hd__a21o_1
X_16453_ _02980_ _06488_ VGND VGND VPWR VPWR _06843_ sky130_fd_sc_hd__or2_1
XFILLER_0_128_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10877_ _04351_ _04373_ _03815_ _03837_ VGND VGND VPWR VPWR _00970_ sky130_fd_sc_hd__and4_1
XFILLER_0_73_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15404_ _05703_ _05706_ VGND VGND VPWR VPWR _05707_ sky130_fd_sc_hd__xor2_1
XFILLER_0_66_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12616_ _02707_ _02708_ VGND VGND VPWR VPWR _02709_ sky130_fd_sc_hd__nor2_1
XFILLER_0_128_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16384_ _06763_ _06767_ VGND VGND VPWR VPWR _06768_ sky130_fd_sc_hd__nor2_1
X_13596_ _03731_ _03732_ VGND VGND VPWR VPWR _03733_ sky130_fd_sc_hd__nor2_1
XFILLER_0_54_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15335_ _01356_ _03055_ _05559_ _05558_ _04900_ VGND VGND VPWR VPWR _05631_ sky130_fd_sc_hd__a32o_1
XFILLER_0_54_766 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18123_ _08616_ _08573_ _08658_ VGND VGND VPWR VPWR _08661_ sky130_fd_sc_hd__and3_1
X_12547_ _00832_ _00180_ _02595_ _02596_ VGND VGND VPWR VPWR _02640_ sky130_fd_sc_hd__a22o_1
XFILLER_0_81_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15266_ _05467_ _05468_ VGND VGND VPWR VPWR _05556_ sky130_fd_sc_hd__or2_1
X_18054_ _08502_ _08585_ VGND VGND VPWR VPWR _08586_ sky130_fd_sc_hd__xnor2_1
X_12478_ _02540_ _02541_ VGND VGND VPWR VPWR _02571_ sky130_fd_sc_hd__or2b_1
XFILLER_0_41_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_3 _00166_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14217_ _04401_ _04410_ _04411_ VGND VGND VPWR VPWR _04412_ sky130_fd_sc_hd__a21oi_2
X_17005_ _07382_ _07383_ _07442_ VGND VGND VPWR VPWR _07443_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_22_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11429_ _01520_ _07559_ _07602_ _01521_ VGND VGND VPWR VPWR _01522_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_112_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15197_ _02996_ _07025_ _00119_ _02993_ VGND VGND VPWR VPWR _05481_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_22_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14148_ _00461_ VGND VGND VPWR VPWR _04336_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_6_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18956_ clknet_4_1_0_clk _09417_ VGND VGND VPWR VPWR salida\[9\] sky130_fd_sc_hd__dfxtp_1
X_14079_ _02979_ _04259_ VGND VGND VPWR VPWR _04260_ sky130_fd_sc_hd__or2_1
XTAP_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17907_ _02173_ _08423_ _08425_ VGND VGND VPWR VPWR _08426_ sky130_fd_sc_hd__a21oi_4
X_18887_ clknet_4_11_0_clk _00041_ VGND VGND VPWR VPWR ApproximateM_inst.lob_16.lob1.genblk1\[5\].genblk1.mux.sel
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_83_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17838_ _08265_ _08273_ VGND VGND VPWR VPWR _08350_ sky130_fd_sc_hd__or2_1
XFILLER_0_83_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer15 _04574_ VGND VGND VPWR VPWR net178 sky130_fd_sc_hd__clkbuf_1
Xrebuffer26 _03810_ VGND VGND VPWR VPWR net189 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_107_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_77 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xrebuffer37 _04432_ VGND VGND VPWR VPWR net200 sky130_fd_sc_hd__clkbuf_1
Xrebuffer48 _03004_ VGND VGND VPWR VPWR net211 sky130_fd_sc_hd__clkbuf_1
X_17769_ _08259_ _08166_ _08274_ VGND VGND VPWR VPWR _08275_ sky130_fd_sc_hd__o21a_1
Xrebuffer59 _05377_ VGND VGND VPWR VPWR net222 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_84 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_146_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09956_ net166 _06906_ _09005_ _09016_ VGND VGND VPWR VPWR _09027_ sky130_fd_sc_hd__o211a_1
XTAP_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09887_ _07919_ _07930_ _08126_ _08267_ VGND VGND VPWR VPWR _08278_ sky130_fd_sc_hd__o211a_1
XFILLER_0_99_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10800_ _00856_ _00891_ _00273_ _00892_ VGND VGND VPWR VPWR _00893_ sky130_fd_sc_hd__o211ai_4
XTAP_2758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11780_ _00164_ VGND VGND VPWR VPWR _01873_ sky130_fd_sc_hd__buf_6
XFILLER_0_138_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10731_ _00797_ _00821_ _06181_ _00822_ VGND VGND VPWR VPWR _00824_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_137_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13450_ _03164_ _03571_ VGND VGND VPWR VPWR _03572_ sky130_fd_sc_hd__or2_1
X_10662_ _00752_ _00753_ _00572_ _00598_ VGND VGND VPWR VPWR _00755_ sky130_fd_sc_hd__o211a_1
XFILLER_0_153_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12401_ _07984_ _07973_ _00909_ _00145_ VGND VGND VPWR VPWR _02494_ sky130_fd_sc_hd__nand4_2
XFILLER_0_35_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13381_ _03321_ _00165_ _00212_ _03322_ VGND VGND VPWR VPWR _03497_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_35_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10593_ _00685_ _00108_ _00511_ VGND VGND VPWR VPWR _00686_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15120_ _05310_ _05395_ VGND VGND VPWR VPWR _05397_ sky130_fd_sc_hd__or2_1
XFILLER_0_90_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12332_ _02423_ _02424_ _05671_ _00146_ VGND VGND VPWR VPWR _02425_ sky130_fd_sc_hd__and4b_1
XFILLER_0_23_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15051_ _05212_ _05314_ _05319_ VGND VGND VPWR VPWR _05321_ sky130_fd_sc_hd__nor3_1
X_12263_ _06993_ _00213_ _02354_ _02355_ VGND VGND VPWR VPWR _02356_ sky130_fd_sc_hd__a31o_1
X_14002_ _00195_ _00702_ _08452_ _04700_ VGND VGND VPWR VPWR _04177_ sky130_fd_sc_hd__and4_1
X_11214_ _01304_ _01305_ _01291_ _01292_ VGND VGND VPWR VPWR _01307_ sky130_fd_sc_hd__a211o_1
XFILLER_0_31_482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12194_ _02268_ _02275_ _02285_ _02286_ VGND VGND VPWR VPWR _02287_ sky130_fd_sc_hd__a211oi_2
X_18810_ _09298_ _09316_ VGND VGND VPWR VPWR _09317_ sky130_fd_sc_hd__and2_1
XFILLER_0_102_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11145_ _01147_ _01148_ _01237_ VGND VGND VPWR VPWR _01238_ sky130_fd_sc_hd__and3_1
Xoutput73 net73 VGND VGND VPWR VPWR leds[1] sky130_fd_sc_hd__buf_2
Xoutput84 net84 VGND VGND VPWR VPWR o_wb_data[10] sky130_fd_sc_hd__clkbuf_4
Xoutput95 net95 VGND VGND VPWR VPWR o_wb_data[20] sky130_fd_sc_hd__clkbuf_4
X_18741_ _09262_ VGND VGND VPWR VPWR _00072_ sky130_fd_sc_hd__buf_1
X_11076_ _01046_ _01045_ VGND VGND VPWR VPWR _01169_ sky130_fd_sc_hd__and2b_1
X_15953_ _06284_ _06285_ _06287_ _06269_ VGND VGND VPWR VPWR _06300_ sky130_fd_sc_hd__a2bb2o_1
X_14904_ _00191_ _05715_ VGND VGND VPWR VPWR _05162_ sky130_fd_sc_hd__and2_1
X_10027_ _07799_ VGND VGND VPWR VPWR _00120_ sky130_fd_sc_hd__clkbuf_4
X_18672_ net37 _00593_ _09193_ VGND VGND VPWR VPWR _09213_ sky130_fd_sc_hd__mux2_1
X_15884_ _06192_ _06226_ VGND VGND VPWR VPWR _06227_ sky130_fd_sc_hd__nor2_1
X_17623_ _08113_ _08114_ VGND VGND VPWR VPWR _08117_ sky130_fd_sc_hd__nor2_1
X_14835_ _03059_ _03076_ _03164_ VGND VGND VPWR VPWR _05087_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17554_ _08020_ _08022_ _08041_ _06723_ _01862_ VGND VGND VPWR VPWR _09393_ sky130_fd_sc_hd__o32a_1
X_14766_ _05009_ _05010_ VGND VGND VPWR VPWR _05011_ sky130_fd_sc_hd__and2_1
X_11978_ _01944_ _01973_ _01974_ _01975_ VGND VGND VPWR VPWR _02071_ sky130_fd_sc_hd__nor4_1
X_16505_ _06897_ _06898_ VGND VGND VPWR VPWR _06899_ sky130_fd_sc_hd__xor2_2
X_13717_ _00125_ _04143_ _04154_ _00151_ VGND VGND VPWR VPWR _03865_ sky130_fd_sc_hd__a22oi_1
X_10929_ _00939_ _00931_ _00938_ VGND VGND VPWR VPWR _01022_ sky130_fd_sc_hd__nand3_1
X_14697_ _04934_ _04935_ VGND VGND VPWR VPWR _04936_ sky130_fd_sc_hd__xor2_2
X_17485_ _07823_ _07839_ VGND VGND VPWR VPWR _07966_ sky130_fd_sc_hd__nor2_1
XFILLER_0_73_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16436_ _06822_ _06823_ VGND VGND VPWR VPWR _06824_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13648_ _03609_ _03616_ _03615_ VGND VGND VPWR VPWR _03789_ sky130_fd_sc_hd__a21o_1
XFILLER_0_73_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13579_ _03697_ _03698_ _03712_ VGND VGND VPWR VPWR _03714_ sky130_fd_sc_hd__and3_1
XFILLER_0_5_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16367_ _06660_ _06663_ _00494_ VGND VGND VPWR VPWR _06749_ sky130_fd_sc_hd__o21a_4
XFILLER_0_42_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18106_ _08640_ VGND VGND VPWR VPWR _08642_ sky130_fd_sc_hd__inv_2
XFILLER_0_143_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15318_ _05524_ _05525_ _05611_ VGND VGND VPWR VPWR _05613_ sky130_fd_sc_hd__nand3_1
X_16298_ _02489_ _00108_ _06673_ VGND VGND VPWR VPWR _06674_ sky130_fd_sc_hd__or3_1
XFILLER_0_2_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18037_ _07303_ _07861_ _08384_ VGND VGND VPWR VPWR _08567_ sky130_fd_sc_hd__or3_1
XFILLER_0_151_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15249_ _03006_ _01695_ VGND VGND VPWR VPWR _05537_ sky130_fd_sc_hd__nand2_1
XFILLER_0_111_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09810_ _07417_ _07428_ VGND VGND VPWR VPWR _07439_ sky130_fd_sc_hd__and2b_1
XFILLER_0_120_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09741_ cla_inst.in1\[22\] VGND VGND VPWR VPWR _06689_ sky130_fd_sc_hd__buf_4
X_18939_ clknet_4_2_0_clk _00093_ VGND VGND VPWR VPWR cla_inst.in2\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_94_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09672_ _05529_ _05867_ _05932_ VGND VGND VPWR VPWR _05943_ sky130_fd_sc_hd__nand3_4
XFILLER_0_118_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_80 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_119_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_298 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_123 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09939_ _05649_ _06722_ _05704_ _05573_ VGND VGND VPWR VPWR _08843_ sky130_fd_sc_hd__a22o_1
Xclkbuf_4_13_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_13_0_clk sky130_fd_sc_hd__clkbuf_8
X_12950_ _03040_ _03042_ VGND VGND VPWR VPWR _03043_ sky130_fd_sc_hd__nand2_1
X_11901_ _01747_ _01993_ VGND VGND VPWR VPWR _01994_ sky130_fd_sc_hd__xor2_2
X_12881_ _02973_ VGND VGND VPWR VPWR _02974_ sky130_fd_sc_hd__clkbuf_4
XTAP_2500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14620_ _04713_ _04718_ _04712_ VGND VGND VPWR VPWR _04851_ sky130_fd_sc_hd__a21bo_1
X_11832_ _01922_ _01923_ _01924_ VGND VGND VPWR VPWR _01925_ sky130_fd_sc_hd__a21bo_1
XTAP_2544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14551_ _04480_ _04662_ VGND VGND VPWR VPWR _04776_ sky130_fd_sc_hd__or2_1
XTAP_1843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11763_ _01852_ _01855_ VGND VGND VPWR VPWR _01856_ sky130_fd_sc_hd__xor2_1
XTAP_1854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_102 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13502_ _03627_ _03628_ VGND VGND VPWR VPWR _03630_ sky130_fd_sc_hd__xnor2_1
X_10714_ _06591_ _04569_ _04449_ _00806_ VGND VGND VPWR VPWR _00807_ sky130_fd_sc_hd__a22o_1
XTAP_1887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17270_ _07703_ _07704_ _07729_ _07730_ VGND VGND VPWR VPWR _07731_ sky130_fd_sc_hd__o211a_1
X_14482_ _04598_ _04599_ _04605_ VGND VGND VPWR VPWR _04701_ sky130_fd_sc_hd__nand3_2
XTAP_1898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11694_ _01751_ _01785_ _01783_ _01786_ VGND VGND VPWR VPWR _01787_ sky130_fd_sc_hd__o211a_1
XFILLER_0_153_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16221_ _06513_ _06586_ _06587_ _06588_ _06589_ VGND VGND VPWR VPWR _06590_ sky130_fd_sc_hd__a311o_1
XFILLER_0_126_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13433_ _03552_ _03554_ _02489_ VGND VGND VPWR VPWR _03555_ sky130_fd_sc_hd__mux2_1
X_10645_ _00735_ _00736_ _00719_ _00720_ VGND VGND VPWR VPWR _00738_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_125_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_894 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16152_ op_code\[2\] op_code\[3\] VGND VGND VPWR VPWR _06516_ sky130_fd_sc_hd__and2_2
X_13364_ _01505_ _00557_ _03300_ _03299_ VGND VGND VPWR VPWR _03479_ sky130_fd_sc_hd__a31o_1
X_10576_ _07047_ _07080_ _09256_ _09303_ VGND VGND VPWR VPWR _00669_ sky130_fd_sc_hd__nand4_2
Xrebuffer6 _03498_ VGND VGND VPWR VPWR net169 sky130_fd_sc_hd__buf_4
XFILLER_0_24_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15103_ _05273_ _05274_ _05271_ VGND VGND VPWR VPWR _05379_ sky130_fd_sc_hd__o21ai_1
X_12315_ _02407_ _02359_ _02358_ VGND VGND VPWR VPWR _02408_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_133_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16083_ _03107_ _06440_ VGND VGND VPWR VPWR _06441_ sky130_fd_sc_hd__and2_1
X_13295_ _03400_ _03401_ _03396_ VGND VGND VPWR VPWR _03403_ sky130_fd_sc_hd__a21o_1
X_15034_ _05302_ _05303_ VGND VGND VPWR VPWR _05304_ sky130_fd_sc_hd__and2_1
X_12246_ _02246_ _02338_ VGND VGND VPWR VPWR _02339_ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12177_ _02268_ _02269_ VGND VGND VPWR VPWR _02270_ sky130_fd_sc_hd__nand2_1
X_11128_ _07700_ _05257_ _01220_ VGND VGND VPWR VPWR _01221_ sky130_fd_sc_hd__and3_2
X_16985_ _07419_ _07420_ VGND VGND VPWR VPWR _07421_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_3_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18724_ net59 _09190_ _09249_ VGND VGND VPWR VPWR _00067_ sky130_fd_sc_hd__o21a_1
XFILLER_0_64_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11059_ _04078_ _01151_ _00176_ _00145_ VGND VGND VPWR VPWR _01152_ sky130_fd_sc_hd__and4_1
X_15936_ _06242_ _06254_ _06281_ VGND VGND VPWR VPWR _06282_ sky130_fd_sc_hd__a21oi_1
X_18655_ _09176_ _09199_ VGND VGND VPWR VPWR _09200_ sky130_fd_sc_hd__and2_1
X_15867_ _06157_ _06205_ _06206_ VGND VGND VPWR VPWR _06208_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_154_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17606_ _08084_ _08097_ VGND VGND VPWR VPWR _08098_ sky130_fd_sc_hd__xnor2_1
X_14818_ _05065_ _05066_ _04965_ _04966_ VGND VGND VPWR VPWR _05068_ sky130_fd_sc_hd__a211o_1
X_18586_ net297 _09140_ _09148_ _09144_ VGND VGND VPWR VPWR _00016_ sky130_fd_sc_hd__o211a_1
XFILLER_0_148_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15798_ _06065_ _06068_ _06133_ VGND VGND VPWR VPWR _06134_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_86_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17537_ _02989_ _06510_ _01862_ VGND VGND VPWR VPWR _08023_ sky130_fd_sc_hd__a21o_1
X_14749_ _04989_ _04990_ _04991_ VGND VGND VPWR VPWR _04992_ sky130_fd_sc_hd__nand3_1
XFILLER_0_46_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_129_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17468_ _07945_ _07946_ VGND VGND VPWR VPWR _07947_ sky130_fd_sc_hd__nor2_1
XFILLER_0_74_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16419_ _01151_ ApproximateM_inst.lob_16.lob2.genblk1\[14\].genblk1.mux.sel _03184_
+ VGND VGND VPWR VPWR _06805_ sky130_fd_sc_hd__o21a_1
XFILLER_0_116_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_500 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17399_ _07753_ _07754_ _07750_ VGND VGND VPWR VPWR _07872_ sky130_fd_sc_hd__o21a_1
XFILLER_0_55_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_719 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_144_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_747 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_663 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09724_ _06450_ _06493_ VGND VGND VPWR VPWR _06504_ sky130_fd_sc_hd__xnor2_2
X_09655_ _05715_ VGND VGND VPWR VPWR _05758_ sky130_fd_sc_hd__buf_4
X_09586_ _04995_ _03935_ _03925_ VGND VGND VPWR VPWR _05006_ sky130_fd_sc_hd__a21oi_2
XTAP_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_307 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_108_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_535 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_135_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10430_ _00521_ _00522_ VGND VGND VPWR VPWR _00523_ sky130_fd_sc_hd__xor2_1
XFILLER_0_73_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_104_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10361_ _00282_ _00285_ _00283_ VGND VGND VPWR VPWR _00454_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_115_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_216 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12100_ _02190_ _02192_ VGND VGND VPWR VPWR _02193_ sky130_fd_sc_hd__or2_1
X_13080_ _03168_ _03171_ _03048_ VGND VGND VPWR VPWR _03172_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10292_ _09353_ _00223_ _00238_ _00237_ VGND VGND VPWR VPWR _00385_ sky130_fd_sc_hd__a31o_1
XFILLER_0_131_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12031_ _01575_ VGND VGND VPWR VPWR _02124_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_109_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16770_ _03198_ _04257_ _07182_ _07186_ VGND VGND VPWR VPWR _07187_ sky130_fd_sc_hd__a211o_1
X_13982_ _04152_ _00398_ _07526_ _04153_ VGND VGND VPWR VPWR _04155_ sky130_fd_sc_hd__and4b_1
X_15721_ _06049_ _05985_ VGND VGND VPWR VPWR _06050_ sky130_fd_sc_hd__or2_1
X_12933_ _03025_ VGND VGND VPWR VPWR _03026_ sky130_fd_sc_hd__clkbuf_4
X_18440_ _08999_ _09002_ VGND VGND VPWR VPWR _09003_ sky130_fd_sc_hd__xnor2_1
X_15652_ _02991_ _09351_ _00495_ _07744_ VGND VGND VPWR VPWR _05976_ sky130_fd_sc_hd__nand4_1
XTAP_2330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12864_ _02951_ _02956_ VGND VGND VPWR VPWR _02957_ sky130_fd_sc_hd__or2b_1
XTAP_2341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_806 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14603_ _04726_ _04732_ VGND VGND VPWR VPWR _04833_ sky130_fd_sc_hd__nand2_2
XTAP_2363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18371_ _08927_ _08928_ VGND VGND VPWR VPWR _08929_ sky130_fd_sc_hd__or2_1
X_11815_ _01905_ _01907_ VGND VGND VPWR VPWR _01908_ sky130_fd_sc_hd__xnor2_1
XTAP_2374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15583_ _00115_ _00495_ VGND VGND VPWR VPWR _05901_ sky130_fd_sc_hd__nand2_1
X_12795_ _01500_ _01499_ _01450_ _01447_ VGND VGND VPWR VPWR _02888_ sky130_fd_sc_hd__o211a_2
XTAP_1640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_422 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17322_ _07786_ _07787_ VGND VGND VPWR VPWR _07789_ sky130_fd_sc_hd__or2b_1
X_14534_ _04609_ _04699_ _04754_ _04757_ VGND VGND VPWR VPWR _04758_ sky130_fd_sc_hd__a211o_1
X_11746_ _01837_ _01838_ VGND VGND VPWR VPWR _01839_ sky130_fd_sc_hd__and2_1
XFILLER_0_50_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17253_ _06653_ _07486_ _07593_ net331 VGND VGND VPWR VPWR _07713_ sky130_fd_sc_hd__o22a_1
XFILLER_0_154_855 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14465_ _04564_ _04565_ net217 _04682_ VGND VGND VPWR VPWR _04683_ sky130_fd_sc_hd__a211oi_4
X_11677_ _01760_ _01761_ _01768_ VGND VGND VPWR VPWR _01770_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_154_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16204_ _06571_ VGND VGND VPWR VPWR _06572_ sky130_fd_sc_hd__clkbuf_4
X_10628_ _00545_ _00550_ VGND VGND VPWR VPWR _00721_ sky130_fd_sc_hd__nand2_1
X_13416_ _03535_ VGND VGND VPWR VPWR _03536_ sky130_fd_sc_hd__buf_4
XFILLER_0_126_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14396_ _04598_ net188 _04605_ VGND VGND VPWR VPWR _04607_ sky130_fd_sc_hd__a21oi_2
X_17184_ _07630_ _07130_ _07521_ _07519_ VGND VGND VPWR VPWR _07638_ sky130_fd_sc_hd__o31a_1
XFILLER_0_52_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13347_ _03450_ _03451_ _03459_ VGND VGND VPWR VPWR _03460_ sky130_fd_sc_hd__a21oi_1
X_16135_ _03089_ _06496_ VGND VGND VPWR VPWR _06497_ sky130_fd_sc_hd__or2_1
X_10559_ _00649_ _00650_ _00646_ _00472_ VGND VGND VPWR VPWR _00652_ sky130_fd_sc_hd__a211o_1
XFILLER_0_59_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13278_ _03881_ _03782_ _08049_ VGND VGND VPWR VPWR _03384_ sky130_fd_sc_hd__and3_1
X_16066_ _03239_ _03217_ VGND VGND VPWR VPWR _06422_ sky130_fd_sc_hd__nand2_2
X_15017_ _05283_ _05284_ VGND VGND VPWR VPWR _05285_ sky130_fd_sc_hd__nand2_1
X_12229_ _02160_ _02159_ VGND VGND VPWR VPWR _02322_ sky130_fd_sc_hd__nor2_1
XFILLER_0_121_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16968_ _06657_ _07108_ _07292_ VGND VGND VPWR VPWR _07402_ sky130_fd_sc_hd__and3_1
X_18707_ net53 _03143_ _09182_ VGND VGND VPWR VPWR _09236_ sky130_fd_sc_hd__mux2_1
X_15919_ _06232_ _06235_ _06263_ VGND VGND VPWR VPWR _06264_ sky130_fd_sc_hd__and3_1
XFILLER_0_78_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16899_ _07324_ _07326_ VGND VGND VPWR VPWR _07327_ sky130_fd_sc_hd__xnor2_1
X_09440_ _03399_ VGND VGND VPWR VPWR _03410_ sky130_fd_sc_hd__buf_6
X_18638_ _09185_ VGND VGND VPWR VPWR _00036_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_148_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18569_ net261 _09098_ _09135_ _09126_ VGND VGND VPWR VPWR _00010_ sky130_fd_sc_hd__o211a_1
XFILLER_0_86_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_131_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09707_ _06277_ _06309_ VGND VGND VPWR VPWR _06319_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_97_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09638_ _05562_ VGND VGND VPWR VPWR _05573_ sky130_fd_sc_hd__buf_2
XFILLER_0_97_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09569_ _04777_ _04799_ _04788_ VGND VGND VPWR VPWR _04821_ sky130_fd_sc_hd__a21o_1
X_11600_ _01105_ _00514_ _01692_ _05845_ VGND VGND VPWR VPWR _01693_ sky130_fd_sc_hd__or4b_4
XFILLER_0_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12580_ _02644_ _02645_ _02651_ VGND VGND VPWR VPWR _02673_ sky130_fd_sc_hd__a21o_1
XFILLER_0_136_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_764 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11531_ _01566_ _01567_ _01565_ VGND VGND VPWR VPWR _01624_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_81_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14250_ _04289_ _04291_ VGND VGND VPWR VPWR _04447_ sky130_fd_sc_hd__nand2_1
XFILLER_0_92_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_123_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11462_ _01553_ _01554_ VGND VGND VPWR VPWR _01555_ sky130_fd_sc_hd__nand2_1
XFILLER_0_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13201_ _03300_ _03301_ VGND VGND VPWR VPWR _03302_ sky130_fd_sc_hd__xor2_1
XFILLER_0_33_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10413_ _00496_ _00505_ VGND VGND VPWR VPWR _00506_ sky130_fd_sc_hd__xnor2_2
X_14181_ _04357_ _04358_ _04371_ VGND VGND VPWR VPWR _04372_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_21_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11393_ _01469_ _01485_ VGND VGND VPWR VPWR _01486_ sky130_fd_sc_hd__xnor2_1
X_13132_ _00294_ _05606_ _05617_ _04351_ VGND VGND VPWR VPWR _03229_ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10344_ _00276_ _00277_ _00275_ VGND VGND VPWR VPWR _00437_ sky130_fd_sc_hd__a21bo_1
XTAP_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13063_ _03154_ VGND VGND VPWR VPWR _03155_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_103_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17940_ _08357_ _08460_ VGND VGND VPWR VPWR _08461_ sky130_fd_sc_hd__nand2_1
X_10275_ _00349_ _00350_ _00367_ VGND VGND VPWR VPWR _00368_ sky130_fd_sc_hd__a21oi_1
X_12014_ _02090_ _02105_ _02106_ _02050_ VGND VGND VPWR VPWR _02107_ sky130_fd_sc_hd__o211a_4
X_17871_ _07630_ _07861_ _08385_ VGND VGND VPWR VPWR _08386_ sky130_fd_sc_hd__nor3_1
X_16822_ _07241_ _07148_ _07242_ VGND VGND VPWR VPWR _07244_ sky130_fd_sc_hd__a21o_1
XFILLER_0_45_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16753_ _06989_ _07094_ _07095_ VGND VGND VPWR VPWR _07169_ sky130_fd_sc_hd__o21a_1
X_13965_ _04134_ _04135_ VGND VGND VPWR VPWR _04136_ sky130_fd_sc_hd__xnor2_1
Xmax_cap4 _02293_ VGND VGND VPWR VPWR net322 sky130_fd_sc_hd__clkbuf_1
X_15704_ _03007_ _03055_ _06031_ VGND VGND VPWR VPWR _06032_ sky130_fd_sc_hd__nand3_1
X_12916_ _03008_ VGND VGND VPWR VPWR _03009_ sky130_fd_sc_hd__buf_2
X_16684_ _03790_ _06509_ _02214_ VGND VGND VPWR VPWR _07094_ sky130_fd_sc_hd__a21oi_1
X_13896_ _03847_ _03849_ _03852_ _03854_ VGND VGND VPWR VPWR _04061_ sky130_fd_sc_hd__a31oi_2
X_18423_ _02920_ net115 _03201_ VGND VGND VPWR VPWR _08986_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_152_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15635_ _05929_ VGND VGND VPWR VPWR _05957_ sky130_fd_sc_hd__inv_2
XTAP_2160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12847_ _02939_ VGND VGND VPWR VPWR _02940_ sky130_fd_sc_hd__inv_2
XTAP_2171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18354_ _08909_ _08910_ VGND VGND VPWR VPWR _08911_ sky130_fd_sc_hd__xnor2_1
X_15566_ _03007_ _01112_ VGND VGND VPWR VPWR _05882_ sky130_fd_sc_hd__nand2_1
XTAP_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12778_ _02869_ _02870_ VGND VGND VPWR VPWR _02871_ sky130_fd_sc_hd__and2_1
XFILLER_0_28_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17305_ _07618_ _07642_ _07617_ VGND VGND VPWR VPWR _07770_ sky130_fd_sc_hd__o21ba_1
X_14517_ _04702_ _04703_ _04737_ _04738_ VGND VGND VPWR VPWR _04739_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_84_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18285_ _08751_ _08813_ _08814_ VGND VGND VPWR VPWR _08836_ sky130_fd_sc_hd__o21ba_1
X_11729_ ApproximateM_inst.lob_16.lob2.genblk1\[11\].genblk1.mux.sel _00177_ VGND
+ VGND VPWR VPWR _01822_ sky130_fd_sc_hd__nand2_1
X_15497_ _02975_ _05805_ _05806_ VGND VGND VPWR VPWR _05807_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_127_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17236_ _06368_ _06438_ _07694_ VGND VGND VPWR VPWR _07695_ sky130_fd_sc_hd__o21a_1
XFILLER_0_117_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14448_ _04651_ _04652_ _04663_ VGND VGND VPWR VPWR _04664_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_142_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17167_ _07617_ _07618_ VGND VGND VPWR VPWR _07619_ sky130_fd_sc_hd__nor2_1
XFILLER_0_25_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14379_ _02188_ _09256_ _07755_ VGND VGND VPWR VPWR _04588_ sky130_fd_sc_hd__and3_1
XFILLER_0_4_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16118_ _03029_ _01746_ _01503_ _03083_ _06477_ _03161_ VGND VGND VPWR VPWR _06478_
+ sky130_fd_sc_hd__mux4_1
X_17098_ _06665_ _07314_ VGND VGND VPWR VPWR _07544_ sky130_fd_sc_hd__nor2_1
XFILLER_0_110_744 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16049_ _01417_ _03143_ VGND VGND VPWR VPWR _06403_ sky130_fd_sc_hd__or2_2
XFILLER_0_79_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09423_ _03217_ _03206_ VGND VGND VPWR VPWR _03228_ sky130_fd_sc_hd__nor2_1
XFILLER_0_149_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_118_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_91 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_144_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10060_ _09352_ _00147_ _00150_ _00152_ VGND VGND VPWR VPWR _00153_ sky130_fd_sc_hd__nand4_1
X_13750_ _03732_ _03735_ _03731_ VGND VGND VPWR VPWR _03901_ sky130_fd_sc_hd__o21ba_2
X_10962_ _06591_ _03804_ _03826_ _00806_ VGND VGND VPWR VPWR _01055_ sky130_fd_sc_hd__a22o_1
XFILLER_0_98_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12701_ _02792_ _02793_ VGND VGND VPWR VPWR _02794_ sky130_fd_sc_hd__and2_1
X_13681_ _03823_ _03824_ VGND VGND VPWR VPWR _03825_ sky130_fd_sc_hd__and2_1
X_10893_ _05290_ _03739_ _03804_ ApproximateM_inst.lob_16.lob2.genblk1\[10\].genblk1.mux.sel
+ VGND VGND VPWR VPWR _00986_ sky130_fd_sc_hd__a22o_1
X_15420_ _02991_ _08876_ _05721_ VGND VGND VPWR VPWR _05723_ sky130_fd_sc_hd__and3_1
XFILLER_0_109_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12632_ _02722_ _02723_ _02724_ VGND VGND VPWR VPWR _02725_ sky130_fd_sc_hd__or3_1
XFILLER_0_93_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15351_ _05569_ _05567_ VGND VGND VPWR VPWR _05648_ sky130_fd_sc_hd__and2b_1
XFILLER_0_108_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12563_ _02618_ _02625_ VGND VGND VPWR VPWR _02656_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_25_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14302_ _01745_ _04336_ VGND VGND VPWR VPWR _04505_ sky130_fd_sc_hd__nand2_1
X_11514_ _01164_ _01156_ _01163_ VGND VGND VPWR VPWR _01607_ sky130_fd_sc_hd__nand3_1
XFILLER_0_80_222 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18070_ _07002_ _08036_ _03197_ _05881_ VGND VGND VPWR VPWR _08603_ sky130_fd_sc_hd__a2bb2o_1
X_15282_ _05571_ _05572_ VGND VGND VPWR VPWR _05574_ sky130_fd_sc_hd__nand2_1
X_12494_ _02584_ _02586_ VGND VGND VPWR VPWR _02587_ sky130_fd_sc_hd__and2_1
XFILLER_0_124_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire132 _08451_ VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17021_ _07386_ _07355_ _00399_ VGND VGND VPWR VPWR _07460_ sky130_fd_sc_hd__o21a_1
X_14233_ _04283_ net133 _04295_ VGND VGND VPWR VPWR _04429_ sky130_fd_sc_hd__nor3_2
X_11445_ _06460_ _00878_ _01536_ _01537_ _00193_ VGND VGND VPWR VPWR _01538_ sky130_fd_sc_hd__a32o_1
XFILLER_0_123_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14164_ _04337_ _04353_ VGND VGND VPWR VPWR _04354_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_22_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11376_ _01409_ _01411_ _01407_ VGND VGND VPWR VPWR _01469_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13115_ _03207_ _03208_ _03209_ VGND VGND VPWR VPWR _03210_ sky130_fd_sc_hd__nand3_1
X_10327_ _00245_ _00267_ VGND VGND VPWR VPWR _00420_ sky130_fd_sc_hd__nand2_1
X_14095_ _04132_ _07156_ _06732_ _04099_ VGND VGND VPWR VPWR _04278_ sky130_fd_sc_hd__a22o_1
X_18972_ clknet_4_5_0_clk _09403_ VGND VGND VPWR VPWR salida\[25\] sky130_fd_sc_hd__dfxtp_1
XTAP_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17923_ _08434_ _08436_ _08439_ _08443_ VGND VGND VPWR VPWR _08444_ sky130_fd_sc_hd__and4b_1
X_13046_ _03135_ _03137_ _03048_ VGND VGND VPWR VPWR _03138_ sky130_fd_sc_hd__mux2_1
X_10258_ _07700_ _07799_ cla_inst.in1\[31\] _09256_ VGND VGND VPWR VPWR _00351_ sky130_fd_sc_hd__nand4_1
X_17854_ _07608_ _07314_ _07516_ _07195_ VGND VGND VPWR VPWR _08368_ sky130_fd_sc_hd__o22a_1
X_10189_ _04121_ _04580_ _04460_ _04088_ VGND VGND VPWR VPWR _00282_ sky130_fd_sc_hd__a22oi_2
X_16805_ _07121_ _07119_ VGND VGND VPWR VPWR _07225_ sky130_fd_sc_hd__and2b_1
X_17785_ _08257_ _08258_ _08291_ VGND VGND VPWR VPWR _08293_ sky130_fd_sc_hd__and3_1
X_14997_ _05168_ _05167_ VGND VGND VPWR VPWR _05263_ sky130_fd_sc_hd__or2b_1
X_16736_ _07017_ _07048_ VGND VGND VPWR VPWR _07150_ sky130_fd_sc_hd__nor2_1
X_13948_ _03954_ _03955_ _04116_ VGND VGND VPWR VPWR _04117_ sky130_fd_sc_hd__o21a_1
XFILLER_0_88_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16667_ _02800_ _07073_ _07074_ VGND VGND VPWR VPWR _07075_ sky130_fd_sc_hd__o21a_1
X_13879_ _04025_ _04026_ _04040_ VGND VGND VPWR VPWR _04042_ sky130_fd_sc_hd__and3_1
XFILLER_0_29_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18406_ _08965_ _08966_ VGND VGND VPWR VPWR _08967_ sky130_fd_sc_hd__xor2_1
X_15618_ _05861_ net118 _05937_ VGND VGND VPWR VPWR _05939_ sky130_fd_sc_hd__or3b_1
XFILLER_0_57_742 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16598_ _06696_ _06701_ _03060_ VGND VGND VPWR VPWR _07000_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18337_ _03143_ _06464_ _08839_ _08892_ VGND VGND VPWR VPWR _09404_ sky130_fd_sc_hd__o2bb2a_1
X_15549_ _05863_ VGND VGND VPWR VPWR _05864_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_639 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_814 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_154_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18268_ _08815_ _08816_ _08817_ VGND VGND VPWR VPWR _08818_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_21_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_244 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_141_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17219_ _02669_ _02670_ _07562_ VGND VGND VPWR VPWR _07676_ sky130_fd_sc_hd__o21a_1
X_18199_ _08587_ _08742_ VGND VGND VPWR VPWR _08743_ sky130_fd_sc_hd__or2_1
XFILLER_0_141_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_141_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09972_ cla_inst.in2\[29\] VGND VGND VPWR VPWR _09172_ sky130_fd_sc_hd__buf_2
XFILLER_0_12_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_731 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_153_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_195 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11230_ _01320_ _01322_ VGND VGND VPWR VPWR _01323_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_120_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_121_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11161_ cla_inst.in2\[22\] _09212_ VGND VGND VPWR VPWR _01254_ sky130_fd_sc_hd__and2_1
XFILLER_0_113_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10112_ _04220_ VGND VGND VPWR VPWR _00205_ sky130_fd_sc_hd__clkbuf_8
X_11092_ _05508_ _05464_ _04143_ _04056_ VGND VGND VPWR VPWR _01185_ sky130_fd_sc_hd__nand4_1
X_14920_ _05161_ _05178_ VGND VGND VPWR VPWR _05179_ sky130_fd_sc_hd__xnor2_1
X_10043_ _09353_ _00134_ _00135_ _00128_ VGND VGND VPWR VPWR _00136_ sky130_fd_sc_hd__a22oi_1
X_14851_ _02986_ _07733_ _05101_ _05102_ VGND VGND VPWR VPWR _05103_ sky130_fd_sc_hd__a22oi_4
Xhold84 op_code\[1\] VGND VGND VPWR VPWR net247 sky130_fd_sc_hd__buf_1
Xhold95 _00025_ VGND VGND VPWR VPWR net258 sky130_fd_sc_hd__dlygate4sd3_1
X_13802_ _03955_ _03956_ VGND VGND VPWR VPWR _03958_ sky130_fd_sc_hd__or2_1
XFILLER_0_98_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17570_ _07143_ _07387_ _08055_ _08057_ VGND VGND VPWR VPWR _08058_ sky130_fd_sc_hd__nor4_1
X_14782_ _05018_ _05027_ VGND VGND VPWR VPWR _05029_ sky130_fd_sc_hd__xor2_1
XFILLER_0_97_130 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11994_ _02084_ _02085_ _02086_ VGND VGND VPWR VPWR _02087_ sky130_fd_sc_hd__o21ba_1
X_16521_ _06639_ _06632_ _06627_ _06641_ _03080_ _03077_ VGND VGND VPWR VPWR _06916_
+ sky130_fd_sc_hd__mux4_2
X_13733_ _03879_ _03880_ _03836_ _03715_ VGND VGND VPWR VPWR _03883_ sky130_fd_sc_hd__o211a_1
XFILLER_0_58_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10945_ _01028_ _01036_ _01037_ VGND VGND VPWR VPWR _01038_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_97_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16452_ _06839_ _06840_ VGND VGND VPWR VPWR _06842_ sky130_fd_sc_hd__xnor2_1
X_13664_ _03788_ _03805_ _03806_ VGND VGND VPWR VPWR _03807_ sky130_fd_sc_hd__nand3_2
X_10876_ _05017_ _03750_ VGND VGND VPWR VPWR _00969_ sky130_fd_sc_hd__nand2_1
XFILLER_0_27_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15403_ _05705_ _05591_ _05588_ VGND VGND VPWR VPWR _05706_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_54_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12615_ _02705_ _02706_ _02701_ _02704_ VGND VGND VPWR VPWR _02708_ sky130_fd_sc_hd__o211a_1
X_16383_ _06579_ _06653_ _06766_ _06561_ VGND VGND VPWR VPWR _06767_ sky130_fd_sc_hd__o22a_1
X_13595_ _03518_ _03521_ _03730_ VGND VGND VPWR VPWR _03732_ sky130_fd_sc_hd__nor3b_4
XFILLER_0_93_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18122_ _08616_ _08573_ _08658_ VGND VGND VPWR VPWR _08660_ sky130_fd_sc_hd__a21oi_1
X_15334_ _05556_ _05565_ VGND VGND VPWR VPWR _05630_ sky130_fd_sc_hd__and2_1
XFILLER_0_53_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12546_ _02636_ _02637_ _02638_ VGND VGND VPWR VPWR _02639_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_136_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18053_ _08582_ _08584_ VGND VGND VPWR VPWR _08585_ sky130_fd_sc_hd__or2_1
X_15265_ _05476_ _05473_ VGND VGND VPWR VPWR _05555_ sky130_fd_sc_hd__and2b_1
X_12477_ _02568_ _02569_ VGND VGND VPWR VPWR _02570_ sky130_fd_sc_hd__or2_1
XFILLER_0_151_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_4 _00181_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17004_ _07434_ _07441_ VGND VGND VPWR VPWR _07442_ sky130_fd_sc_hd__xnor2_1
X_14216_ _04401_ _04410_ _03202_ VGND VGND VPWR VPWR _04411_ sky130_fd_sc_hd__o21ai_1
X_11428_ _03574_ VGND VGND VPWR VPWR _01521_ sky130_fd_sc_hd__buf_4
X_15196_ _05478_ _05479_ VGND VGND VPWR VPWR _05480_ sky130_fd_sc_hd__nand2_1
XFILLER_0_22_686 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14147_ _04148_ _04163_ VGND VGND VPWR VPWR _04335_ sky130_fd_sc_hd__nand2_1
X_11359_ _01436_ _01416_ VGND VGND VPWR VPWR _01452_ sky130_fd_sc_hd__or2b_1
XFILLER_0_120_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18955_ clknet_4_1_0_clk _09416_ VGND VGND VPWR VPWR salida\[8\] sky130_fd_sc_hd__dfxtp_1
X_14078_ _03567_ _03581_ _02980_ VGND VGND VPWR VPWR _04259_ sky130_fd_sc_hd__mux2_1
XTAP_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13029_ _02976_ _03035_ _03039_ _03118_ _03121_ VGND VGND VPWR VPWR _03122_ sky130_fd_sc_hd__o32a_1
X_17906_ _04238_ _08424_ VGND VGND VPWR VPWR _08425_ sky130_fd_sc_hd__or2_1
X_18886_ clknet_4_13_0_clk _00040_ VGND VGND VPWR VPWR ApproximateM_inst.lob_16.lob1.genblk1\[4\].genblk1.mux.sel
+ sky130_fd_sc_hd__dfxtp_1
X_17837_ _08263_ _08264_ VGND VGND VPWR VPWR _08349_ sky130_fd_sc_hd__nand2_1
XFILLER_0_83_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer16 _04574_ VGND VGND VPWR VPWR net179 sky130_fd_sc_hd__clkbuf_1
Xrebuffer27 net337 VGND VGND VPWR VPWR net190 sky130_fd_sc_hd__clkbuf_1
Xrebuffer38 _04432_ VGND VGND VPWR VPWR net201 sky130_fd_sc_hd__buf_1
XFILLER_0_107_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17768_ _08265_ _08273_ VGND VGND VPWR VPWR _08274_ sky130_fd_sc_hd__xor2_1
XFILLER_0_83_89 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xrebuffer49 _03004_ VGND VGND VPWR VPWR net212 sky130_fd_sc_hd__buf_1
XFILLER_0_107_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16719_ _06579_ _07130_ VGND VGND VPWR VPWR _07131_ sky130_fd_sc_hd__or2_1
XFILLER_0_107_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17699_ _08074_ _08076_ _08197_ VGND VGND VPWR VPWR _08199_ sky130_fd_sc_hd__nor3_1
XFILLER_0_9_603 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_119_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_146_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_712 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_135_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_84_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_130_603 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09955_ _08973_ _08984_ _08995_ _08681_ VGND VGND VPWR VPWR _09016_ sky130_fd_sc_hd__a22o_1
XTAP_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09886_ _08126_ _08137_ _08256_ VGND VGND VPWR VPWR _08267_ sky130_fd_sc_hd__nand3_2
XTAP_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10730_ _00797_ _00821_ _06181_ _00822_ VGND VGND VPWR VPWR _00823_ sky130_fd_sc_hd__o211a_2
XFILLER_0_138_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10661_ _00572_ _00598_ _00752_ _00753_ VGND VGND VPWR VPWR _00754_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_138_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12400_ _07243_ _00176_ _00145_ _07221_ VGND VGND VPWR VPWR _02493_ sky130_fd_sc_hd__a22o_1
X_13380_ _03270_ _03272_ VGND VGND VPWR VPWR _03496_ sky130_fd_sc_hd__or2_1
XFILLER_0_91_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10592_ cla_inst.in2\[31\] _00108_ VGND VGND VPWR VPWR _00685_ sky130_fd_sc_hd__nand2_1
XFILLER_0_36_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12331_ _08039_ _00196_ _09212_ _00992_ VGND VGND VPWR VPWR _02424_ sky130_fd_sc_hd__a22o_1
XFILLER_0_91_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15050_ _05212_ _05314_ _05319_ VGND VGND VPWR VPWR _05320_ sky130_fd_sc_hd__o21a_1
X_12262_ _07984_ _07243_ _04220_ _00774_ VGND VGND VPWR VPWR _02355_ sky130_fd_sc_hd__and4_1
X_11213_ _01291_ _01292_ _01304_ _01305_ VGND VGND VPWR VPWR _01306_ sky130_fd_sc_hd__o211ai_2
X_14001_ _00702_ _08452_ _01005_ _00195_ VGND VGND VPWR VPWR _04175_ sky130_fd_sc_hd__a22oi_2
X_12193_ _02195_ _02198_ _02284_ VGND VGND VPWR VPWR _02286_ sky130_fd_sc_hd__and3_1
XFILLER_0_31_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11144_ _01204_ _01236_ VGND VGND VPWR VPWR _01237_ sky130_fd_sc_hd__or2b_1
Xoutput74 net74 VGND VGND VPWR VPWR leds[2] sky130_fd_sc_hd__clkbuf_4
Xoutput85 net85 VGND VGND VPWR VPWR o_wb_data[11] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_128_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput96 net96 VGND VGND VPWR VPWR o_wb_data[21] sky130_fd_sc_hd__clkbuf_4
X_18740_ _09245_ _09261_ VGND VGND VPWR VPWR _09262_ sky130_fd_sc_hd__and2_1
X_11075_ _04548_ _04056_ VGND VGND VPWR VPWR _01168_ sky130_fd_sc_hd__nand2_1
X_15952_ _06232_ _06235_ _06263_ _06297_ VGND VGND VPWR VPWR _06299_ sky130_fd_sc_hd__a211o_1
X_14903_ _05158_ _05160_ VGND VGND VPWR VPWR _05161_ sky130_fd_sc_hd__nor2_1
X_10026_ _08876_ VGND VGND VPWR VPWR _00119_ sky130_fd_sc_hd__buf_4
X_18671_ _09211_ VGND VGND VPWR VPWR _00046_ sky130_fd_sc_hd__buf_1
X_15883_ _06225_ VGND VGND VPWR VPWR _06226_ sky130_fd_sc_hd__inv_2
X_17622_ _08113_ _08114_ VGND VGND VPWR VPWR _08116_ sky130_fd_sc_hd__and2_1
X_14834_ _03921_ _05085_ VGND VGND VPWR VPWR _05086_ sky130_fd_sc_hd__nor2_1
XFILLER_0_53_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17553_ _07256_ _08027_ _08029_ _08040_ VGND VGND VPWR VPWR _08041_ sky130_fd_sc_hd__a31o_1
X_14765_ _05001_ _05008_ VGND VGND VPWR VPWR _05010_ sky130_fd_sc_hd__nand2_1
XFILLER_0_58_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11977_ _02052_ _02068_ _02069_ VGND VGND VPWR VPWR _02070_ sky130_fd_sc_hd__or3_2
X_16504_ _06824_ _06827_ _06822_ VGND VGND VPWR VPWR _06898_ sky130_fd_sc_hd__o21a_1
X_13716_ _03654_ _03656_ VGND VGND VPWR VPWR _03864_ sky130_fd_sc_hd__or2_1
XFILLER_0_86_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17484_ _07954_ _07964_ VGND VGND VPWR VPWR _07965_ sky130_fd_sc_hd__xnor2_1
X_10928_ _00980_ _01019_ _01018_ VGND VGND VPWR VPWR _01021_ sky130_fd_sc_hd__o21a_1
XFILLER_0_58_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14696_ _04798_ _04801_ VGND VGND VPWR VPWR _04935_ sky130_fd_sc_hd__nand2_1
XFILLER_0_117_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16435_ _06769_ _06821_ VGND VGND VPWR VPWR _06823_ sky130_fd_sc_hd__nand2_1
X_13647_ _03637_ _03639_ VGND VGND VPWR VPWR _03788_ sky130_fd_sc_hd__nand2_1
X_10859_ _04558_ _04045_ _00950_ _00951_ VGND VGND VPWR VPWR _00952_ sky130_fd_sc_hd__a31o_1
XFILLER_0_54_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16366_ _03539_ _06734_ _06747_ _06484_ VGND VGND VPWR VPWR _06748_ sky130_fd_sc_hd__o211a_1
X_13578_ _03697_ _03698_ _03712_ VGND VGND VPWR VPWR _03713_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_81_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18105_ _08639_ _07859_ _07109_ _08640_ VGND VGND VPWR VPWR _08641_ sky130_fd_sc_hd__and4b_1
XFILLER_0_143_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15317_ _05524_ _05525_ _05611_ VGND VGND VPWR VPWR _05612_ sky130_fd_sc_hd__a21o_1
X_12529_ _02615_ _02619_ _02621_ VGND VGND VPWR VPWR _02622_ sky130_fd_sc_hd__and3_1
X_16297_ _06585_ VGND VGND VPWR VPWR _06673_ sky130_fd_sc_hd__buf_2
XFILLER_0_41_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18036_ _08470_ _08479_ VGND VGND VPWR VPWR _08566_ sky130_fd_sc_hd__or2b_1
X_15248_ _05534_ _05535_ VGND VGND VPWR VPWR _05536_ sky130_fd_sc_hd__nor2_1
XFILLER_0_111_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15179_ _05237_ _05359_ VGND VGND VPWR VPWR _05461_ sky130_fd_sc_hd__and2b_1
XFILLER_0_10_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09740_ _05573_ _05595_ _05693_ _05606_ VGND VGND VPWR VPWR _06678_ sky130_fd_sc_hd__and4_1
X_18938_ clknet_4_11_0_clk _00092_ VGND VGND VPWR VPWR cla_inst.in2\[24\] sky130_fd_sc_hd__dfxtp_2
.ends

