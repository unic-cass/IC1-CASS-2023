magic
tech sky130A
magscale 1 2
timestamp 1676037725
<< nwell >>
rect -38 261 1694 582
<< pwell >>
rect 1365 157 1655 203
rect 1 21 1655 157
rect 29 -17 63 21
<< scnmos >>
rect 79 47 109 131
rect 163 47 193 131
rect 258 47 288 119
rect 367 47 397 119
rect 463 47 493 131
rect 571 47 601 131
rect 761 47 791 131
rect 846 47 876 131
rect 1034 47 1064 131
rect 1141 47 1171 119
rect 1251 47 1281 119
rect 1346 47 1376 131
rect 1447 47 1477 177
rect 1531 47 1561 177
<< scpmoshvt >>
rect 79 369 109 497
rect 163 369 193 497
rect 258 413 288 497
rect 342 413 372 497
rect 486 345 516 473
rect 570 345 600 473
rect 758 316 788 424
rect 842 316 872 424
rect 1030 369 1060 497
rect 1165 413 1195 497
rect 1249 413 1279 497
rect 1350 369 1380 497
rect 1447 297 1477 497
rect 1531 297 1561 497
<< ndiff >>
rect 27 119 79 131
rect 27 85 35 119
rect 69 85 79 119
rect 27 47 79 85
rect 109 93 163 131
rect 109 59 119 93
rect 153 59 163 93
rect 109 47 163 59
rect 193 119 243 131
rect 412 119 463 131
rect 193 47 258 119
rect 288 107 367 119
rect 288 73 310 107
rect 344 73 367 107
rect 288 47 367 73
rect 397 47 463 119
rect 493 93 571 131
rect 493 59 514 93
rect 548 59 571 93
rect 493 47 571 59
rect 601 93 655 131
rect 601 59 613 93
rect 647 59 655 93
rect 601 47 655 59
rect 709 119 761 131
rect 709 85 717 119
rect 751 85 761 119
rect 709 47 761 85
rect 791 119 846 131
rect 791 85 802 119
rect 836 85 846 119
rect 791 47 846 85
rect 876 101 928 131
rect 876 67 886 101
rect 920 67 928 101
rect 876 47 928 67
rect 982 93 1034 131
rect 982 59 990 93
rect 1024 59 1034 93
rect 982 47 1034 59
rect 1064 119 1126 131
rect 1391 131 1447 177
rect 1296 119 1346 131
rect 1064 47 1141 119
rect 1171 93 1251 119
rect 1171 59 1194 93
rect 1228 59 1251 93
rect 1171 47 1251 59
rect 1281 47 1346 119
rect 1376 119 1447 131
rect 1376 85 1403 119
rect 1437 85 1447 119
rect 1376 47 1447 85
rect 1477 103 1531 177
rect 1477 69 1487 103
rect 1521 69 1531 103
rect 1477 47 1531 69
rect 1561 161 1629 177
rect 1561 127 1587 161
rect 1621 127 1629 161
rect 1561 93 1629 127
rect 1561 59 1587 93
rect 1621 59 1629 93
rect 1561 47 1629 59
<< pdiff >>
rect 27 459 79 497
rect 27 425 35 459
rect 69 425 79 459
rect 27 369 79 425
rect 109 485 163 497
rect 109 451 119 485
rect 153 451 163 485
rect 109 369 163 451
rect 193 413 258 497
rect 288 459 342 497
rect 288 425 298 459
rect 332 425 342 459
rect 288 413 342 425
rect 372 473 471 497
rect 372 413 486 473
rect 193 369 243 413
rect 428 345 486 413
rect 516 461 570 473
rect 516 427 526 461
rect 560 427 570 461
rect 516 345 570 427
rect 600 391 652 473
rect 978 465 1030 497
rect 978 431 986 465
rect 1020 431 1030 465
rect 600 357 610 391
rect 644 357 652 391
rect 600 345 652 357
rect 706 412 758 424
rect 706 378 714 412
rect 748 378 758 412
rect 706 316 758 378
rect 788 362 842 424
rect 788 328 798 362
rect 832 328 842 362
rect 788 316 842 328
rect 872 363 924 424
rect 978 369 1030 431
rect 1060 413 1165 497
rect 1195 465 1249 497
rect 1195 431 1205 465
rect 1239 431 1249 465
rect 1195 413 1249 431
rect 1279 413 1350 497
rect 1060 369 1110 413
rect 872 329 882 363
rect 916 329 924 363
rect 872 316 924 329
rect 1294 369 1350 413
rect 1380 485 1447 497
rect 1380 451 1403 485
rect 1437 451 1447 485
rect 1380 417 1447 451
rect 1380 383 1403 417
rect 1437 383 1447 417
rect 1380 369 1447 383
rect 1395 297 1447 369
rect 1477 475 1531 497
rect 1477 441 1487 475
rect 1521 441 1531 475
rect 1477 401 1531 441
rect 1477 367 1487 401
rect 1521 367 1531 401
rect 1477 297 1531 367
rect 1561 485 1629 497
rect 1561 451 1587 485
rect 1621 451 1629 485
rect 1561 417 1629 451
rect 1561 383 1587 417
rect 1621 383 1629 417
rect 1561 349 1629 383
rect 1561 315 1587 349
rect 1621 315 1629 349
rect 1561 297 1629 315
<< ndiffc >>
rect 35 85 69 119
rect 119 59 153 93
rect 310 73 344 107
rect 514 59 548 93
rect 613 59 647 93
rect 717 85 751 119
rect 802 85 836 119
rect 886 67 920 101
rect 990 59 1024 93
rect 1194 59 1228 93
rect 1403 85 1437 119
rect 1487 69 1521 103
rect 1587 127 1621 161
rect 1587 59 1621 93
<< pdiffc >>
rect 35 425 69 459
rect 119 451 153 485
rect 298 425 332 459
rect 526 427 560 461
rect 986 431 1020 465
rect 610 357 644 391
rect 714 378 748 412
rect 798 328 832 362
rect 1205 431 1239 465
rect 882 329 916 363
rect 1403 451 1437 485
rect 1403 383 1437 417
rect 1487 441 1521 475
rect 1487 367 1521 401
rect 1587 451 1621 485
rect 1587 383 1621 417
rect 1587 315 1621 349
<< poly >>
rect 79 497 109 523
rect 163 497 193 523
rect 258 497 288 523
rect 342 497 372 523
rect 486 473 516 523
rect 570 493 872 523
rect 1030 497 1060 523
rect 1165 497 1195 523
rect 1249 497 1279 523
rect 1350 497 1380 523
rect 1447 497 1477 523
rect 1531 497 1561 523
rect 570 473 600 493
rect 79 265 109 369
rect 163 343 193 369
rect 21 249 109 265
rect 21 215 31 249
rect 65 215 109 249
rect 162 335 193 343
rect 162 219 192 335
rect 258 323 288 413
rect 342 375 372 413
rect 234 307 288 323
rect 330 365 396 375
rect 330 331 346 365
rect 380 331 396 365
rect 758 424 788 450
rect 842 424 872 493
rect 330 321 396 331
rect 486 330 516 345
rect 234 273 244 307
rect 278 279 288 307
rect 463 300 516 330
rect 278 273 397 279
rect 234 257 397 273
rect 258 249 397 257
rect 21 199 109 215
rect 79 131 109 199
rect 157 203 211 219
rect 157 169 167 203
rect 201 169 211 203
rect 157 153 211 169
rect 258 191 325 207
rect 258 157 281 191
rect 315 157 325 191
rect 163 131 193 153
rect 258 141 325 157
rect 258 119 288 141
rect 367 119 397 249
rect 463 219 493 300
rect 570 219 600 345
rect 1165 375 1195 413
rect 758 272 788 316
rect 842 290 872 316
rect 1030 279 1060 369
rect 1141 365 1207 375
rect 1141 331 1157 365
rect 1191 331 1207 365
rect 1141 321 1207 331
rect 1249 315 1279 413
rect 1249 299 1303 315
rect 1249 279 1259 299
rect 646 262 788 272
rect 646 228 662 262
rect 696 248 788 262
rect 979 263 1064 279
rect 696 228 876 248
rect 454 203 508 219
rect 454 169 464 203
rect 498 169 508 203
rect 454 153 508 169
rect 550 203 604 219
rect 646 218 876 228
rect 550 169 560 203
rect 594 176 604 203
rect 594 169 791 176
rect 550 153 791 169
rect 463 131 493 153
rect 569 146 791 153
rect 571 131 601 146
rect 761 131 791 146
rect 846 131 876 218
rect 979 229 989 263
rect 1023 229 1064 263
rect 979 213 1064 229
rect 1034 131 1064 213
rect 1141 265 1259 279
rect 1293 265 1303 299
rect 1350 265 1380 369
rect 1447 265 1477 297
rect 1531 265 1561 297
rect 1141 249 1303 265
rect 1345 249 1399 265
rect 1141 119 1171 249
rect 1345 215 1355 249
rect 1389 215 1399 249
rect 1213 191 1281 207
rect 1345 199 1399 215
rect 1441 249 1561 265
rect 1441 215 1451 249
rect 1485 215 1561 249
rect 1441 199 1561 215
rect 1213 157 1223 191
rect 1257 157 1281 191
rect 1213 141 1281 157
rect 1251 119 1281 141
rect 1346 131 1376 199
rect 1447 177 1477 199
rect 1531 177 1561 199
rect 79 21 109 47
rect 163 21 193 47
rect 258 21 288 47
rect 367 21 397 47
rect 463 21 493 47
rect 571 21 601 47
rect 761 21 791 47
rect 846 21 876 47
rect 1034 21 1064 47
rect 1141 21 1171 47
rect 1251 21 1281 47
rect 1346 21 1376 47
rect 1447 21 1477 47
rect 1531 21 1561 47
<< polycont >>
rect 31 215 65 249
rect 346 331 380 365
rect 244 273 278 307
rect 167 169 201 203
rect 281 157 315 191
rect 1157 331 1191 365
rect 662 228 696 262
rect 464 169 498 203
rect 560 169 594 203
rect 989 229 1023 263
rect 1259 265 1293 299
rect 1355 215 1389 249
rect 1451 215 1485 249
rect 1223 157 1257 191
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1656 561
rect 103 485 169 527
rect 35 459 69 475
rect 103 451 119 485
rect 153 451 169 485
rect 519 461 565 527
rect 282 425 298 459
rect 332 425 397 459
rect 431 425 448 459
rect 35 417 69 425
rect 35 391 133 417
rect 35 383 305 391
rect 99 357 305 383
rect 339 365 380 391
rect 339 357 346 365
rect 29 323 65 349
rect 63 289 65 323
rect 29 249 65 289
rect 29 215 31 249
rect 29 195 65 215
rect 99 161 133 357
rect 312 331 346 357
rect 201 289 213 323
rect 247 307 278 323
rect 244 257 278 273
rect 312 315 380 331
rect 34 127 133 161
rect 167 203 247 219
rect 312 207 346 315
rect 414 281 448 425
rect 519 427 526 461
rect 560 427 565 461
rect 951 465 1020 527
rect 1403 485 1437 527
rect 519 411 565 427
rect 661 425 673 459
rect 707 425 764 459
rect 713 412 764 425
rect 594 357 610 391
rect 644 357 663 391
rect 713 378 714 412
rect 748 378 764 412
rect 713 362 764 378
rect 629 332 663 357
rect 629 298 683 332
rect 201 169 247 203
rect 167 153 247 169
rect 34 119 69 127
rect 34 85 35 119
rect 34 69 69 85
rect 103 59 119 93
rect 153 59 169 93
rect 204 79 247 153
rect 281 191 346 207
rect 315 157 346 191
rect 281 141 346 157
rect 380 247 448 281
rect 649 278 683 298
rect 380 107 414 247
rect 482 203 523 264
rect 448 169 464 203
rect 498 169 523 203
rect 448 143 523 169
rect 557 203 615 264
rect 557 169 560 203
rect 594 169 615 203
rect 557 143 615 169
rect 649 262 696 278
rect 649 228 662 262
rect 649 212 696 228
rect 294 73 310 107
rect 344 73 414 107
rect 490 93 556 109
rect 649 93 683 212
rect 730 135 764 362
rect 103 17 169 59
rect 490 59 514 93
rect 548 59 556 93
rect 597 59 613 93
rect 647 59 683 93
rect 717 119 764 135
rect 751 85 764 119
rect 717 69 764 85
rect 798 425 857 459
rect 891 425 903 459
rect 951 431 986 465
rect 798 362 836 425
rect 951 401 1020 431
rect 1065 431 1205 465
rect 1239 431 1255 465
rect 832 328 836 362
rect 798 119 836 328
rect 798 85 802 119
rect 798 69 836 85
rect 879 363 917 379
rect 879 329 882 363
rect 916 347 917 363
rect 1065 347 1099 431
rect 1305 425 1317 459
rect 1351 425 1369 459
rect 916 329 1099 347
rect 879 313 1099 329
rect 879 117 913 313
rect 949 263 1023 279
rect 949 229 989 263
rect 949 143 1023 229
rect 879 101 920 117
rect 879 67 886 101
rect 490 17 556 59
rect 879 51 920 67
rect 959 93 1025 109
rect 959 59 990 93
rect 1024 59 1025 93
rect 1065 93 1099 313
rect 1133 391 1191 397
rect 1167 365 1191 391
rect 1133 331 1157 357
rect 1133 207 1191 331
rect 1335 333 1369 425
rect 1403 417 1437 451
rect 1403 367 1437 383
rect 1471 475 1553 491
rect 1471 441 1487 475
rect 1521 441 1553 475
rect 1471 401 1553 441
rect 1471 367 1487 401
rect 1521 367 1553 401
rect 1225 323 1293 329
rect 1259 299 1293 323
rect 1335 299 1457 333
rect 1491 299 1553 367
rect 1587 485 1637 527
rect 1621 451 1637 485
rect 1587 417 1637 451
rect 1621 383 1637 417
rect 1587 349 1637 383
rect 1621 315 1637 349
rect 1587 299 1637 315
rect 1225 265 1259 289
rect 1423 265 1457 299
rect 1225 249 1293 265
rect 1327 249 1389 265
rect 1327 215 1355 249
rect 1133 191 1257 207
rect 1133 157 1223 191
rect 1133 141 1257 157
rect 1307 199 1389 215
rect 1423 249 1485 265
rect 1423 215 1451 249
rect 1423 199 1485 215
rect 1065 59 1194 93
rect 1228 59 1244 93
rect 1307 75 1369 199
rect 1403 119 1453 163
rect 1519 145 1553 299
rect 1437 85 1453 119
rect 959 17 1025 59
rect 1403 17 1453 85
rect 1487 103 1553 145
rect 1521 69 1553 103
rect 1487 53 1553 69
rect 1587 161 1638 177
rect 1621 127 1638 161
rect 1587 93 1638 127
rect 1621 59 1638 93
rect 1587 17 1638 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1656 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 397 425 431 459
rect 305 357 339 391
rect 29 289 63 323
rect 213 307 247 323
rect 213 289 244 307
rect 244 289 247 307
rect 673 425 707 459
rect 857 425 891 459
rect 1317 425 1351 459
rect 1133 365 1167 391
rect 1133 357 1157 365
rect 1157 357 1167 365
rect 1225 289 1259 323
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
<< metal1 >>
rect 0 561 1656 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1656 561
rect 0 496 1656 527
rect 385 459 443 465
rect 385 425 397 459
rect 431 456 443 459
rect 661 459 719 465
rect 661 456 673 459
rect 431 428 673 456
rect 431 425 443 428
rect 385 419 443 425
rect 661 425 673 428
rect 707 425 719 459
rect 661 419 719 425
rect 845 459 903 465
rect 845 425 857 459
rect 891 456 903 459
rect 1305 459 1363 465
rect 1305 456 1317 459
rect 891 428 1317 456
rect 891 425 903 428
rect 845 419 903 425
rect 1305 425 1317 428
rect 1351 425 1363 459
rect 1305 419 1363 425
rect 293 391 351 397
rect 293 357 305 391
rect 339 388 351 391
rect 1121 391 1179 397
rect 1121 388 1133 391
rect 339 360 1133 388
rect 339 357 351 360
rect 293 351 351 357
rect 1121 357 1133 360
rect 1167 357 1179 391
rect 1121 351 1179 357
rect 17 323 75 329
rect 17 289 29 323
rect 63 320 75 323
rect 201 323 259 329
rect 201 320 213 323
rect 63 292 213 320
rect 63 289 75 292
rect 17 283 75 289
rect 201 289 213 292
rect 247 320 259 323
rect 1213 323 1271 329
rect 1213 320 1225 323
rect 247 292 1225 320
rect 247 289 259 292
rect 201 283 259 289
rect 1213 289 1225 292
rect 1259 289 1271 323
rect 1213 283 1271 289
rect 0 17 1656 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1656 17
rect 0 -48 1656 -17
<< labels >>
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 8 nsew ground bidirectional
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 9 nsew power bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 7 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 10 nsew power bidirectional abutment
flabel locali s 1501 357 1535 391 0 FreeSans 400 0 0 0 X
port 11 nsew signal output
flabel locali s 29 221 63 255 0 FreeSans 400 0 0 0 S0
port 5 nsew signal input
flabel locali s 29 289 63 323 0 FreeSans 400 0 0 0 S0
port 5 nsew signal input
flabel locali s 213 153 247 187 0 FreeSans 400 0 0 0 A2
port 3 nsew signal input
flabel locali s 213 85 247 119 0 FreeSans 400 0 0 0 A2
port 3 nsew signal input
flabel locali s 489 153 523 187 0 FreeSans 400 0 0 0 A3
port 4 nsew signal input
flabel locali s 489 221 523 255 0 FreeSans 400 0 0 0 A3
port 4 nsew signal input
flabel locali s 581 221 615 255 0 FreeSans 400 0 0 0 S1
port 6 nsew signal input
flabel locali s 581 153 615 187 0 FreeSans 400 0 0 0 S1
port 6 nsew signal input
flabel locali s 949 221 983 255 0 FreeSans 400 0 0 0 A1
port 2 nsew signal input
flabel locali s 949 153 983 187 0 FreeSans 400 0 0 0 A1
port 2 nsew signal input
flabel locali s 1317 153 1351 187 0 FreeSans 400 0 0 0 A0
port 1 nsew signal input
flabel locali s 1317 85 1351 119 0 FreeSans 400 0 0 0 A0
port 1 nsew signal input
flabel locali s 1501 85 1535 119 0 FreeSans 400 0 0 0 X
port 11 nsew signal output
flabel locali s 1501 425 1535 459 0 FreeSans 400 0 0 0 X
port 11 nsew signal output
rlabel comment s 0 0 0 0 4 mux4_2
rlabel locali s 244 257 278 289 1 S0
port 5 nsew signal input
rlabel locali s 201 289 278 323 1 S0
port 5 nsew signal input
rlabel locali s 1225 249 1293 329 1 S0
port 5 nsew signal input
rlabel metal1 s 1213 320 1271 329 1 S0
port 5 nsew signal input
rlabel metal1 s 1213 283 1271 292 1 S0
port 5 nsew signal input
rlabel metal1 s 201 320 259 329 1 S0
port 5 nsew signal input
rlabel metal1 s 201 283 259 292 1 S0
port 5 nsew signal input
rlabel metal1 s 17 320 75 329 1 S0
port 5 nsew signal input
rlabel metal1 s 17 292 1271 320 1 S0
port 5 nsew signal input
rlabel metal1 s 17 283 75 292 1 S0
port 5 nsew signal input
rlabel metal1 s 0 -48 1656 48 1 VGND
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1656 592 1 VPWR
port 10 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1656 544
string GDS_END 1784296
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1770058
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 13.600 41.400 13.600 
<< end >>
