* NGSPICE file created from egd_top_wrapper.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_2 abstract view
.subckt sky130_fd_sc_hd__a311oi_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_1 abstract view
.subckt sky130_fd_sc_hd__nor2b_1 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

.subckt egd_top_wrapper la_data_in_58_43[0] la_data_in_58_43[10] la_data_in_58_43[11]
+ la_data_in_58_43[12] la_data_in_58_43[13] la_data_in_58_43[14] la_data_in_58_43[15]
+ la_data_in_58_43[1] la_data_in_58_43[2] la_data_in_58_43[3] la_data_in_58_43[4]
+ la_data_in_58_43[5] la_data_in_58_43[6] la_data_in_58_43[7] la_data_in_58_43[8]
+ la_data_in_58_43[9] la_data_in_60_59[0] la_data_in_60_59[1] la_data_in_65 la_data_out_23_16[0]
+ la_data_out_23_16[1] la_data_out_23_16[2] la_data_out_23_16[3] la_data_out_23_16[4]
+ la_data_out_23_16[5] la_data_out_23_16[6] la_data_out_23_16[7] la_data_out_26_24[0]
+ la_data_out_26_24[1] la_data_out_26_24[2] la_data_out_30_27[0] la_data_out_30_27[1]
+ la_data_out_30_27[2] la_data_out_30_27[3] vccd1 vssd1 wb_clk_i
XTAP_188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6845_ net89 _0304_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[121\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_50_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3988_ egd_top.BitStream_buffer.BS_buffer\[20\] vssd1 vssd1 vccd1 vccd1 _0502_ sky130_fd_sc_hd__clkbuf_4
X_6776_ net180 _0235_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[44\]
+ sky130_fd_sc_hd__dfxtp_1
X_5727_ _0602_ _0592_ _0688_ _0595_ _2227_ vssd1 vssd1 vccd1 vccd1 _2228_ sky130_fd_sc_hd__o221a_1
X_5658_ _3163_ _3177_ vssd1 vssd1 vccd1 vccd1 _2160_ sky130_fd_sc_hd__nand2_1
X_4609_ _0611_ _0587_ vssd1 vssd1 vccd1 vccd1 _1119_ sky130_fd_sc_hd__or2_1
X_5589_ _1360_ _0463_ vssd1 vssd1 vccd1 vccd1 _2091_ sky130_fd_sc_hd__or2_1
XFILLER_89_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4960_ _0353_ _0400_ vssd1 vssd1 vccd1 vccd1 _1467_ sky130_fd_sc_hd__nand2_1
XFILLER_51_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3911_ _0424_ vssd1 vssd1 vccd1 vccd1 _0425_ sky130_fd_sc_hd__clkbuf_2
X_4891_ _3300_ _0772_ vssd1 vssd1 vccd1 vccd1 _1399_ sky130_fd_sc_hd__nand2_1
XFILLER_44_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3842_ _0348_ _0350_ _0355_ vssd1 vssd1 vccd1 vccd1 _0356_ sky130_fd_sc_hd__o21ai_1
X_5512_ _0371_ _0869_ vssd1 vssd1 vccd1 vccd1 _2015_ sky130_fd_sc_hd__nand2_1
X_3773_ _3087_ _3297_ vssd1 vssd1 vccd1 vccd1 _3307_ sky130_fd_sc_hd__nand2_2
X_6492_ _2802_ _2853_ vssd1 vssd1 vccd1 vccd1 _2854_ sky130_fd_sc_hd__nand2_1
X_5443_ _3027_ _1944_ _1946_ vssd1 vssd1 vccd1 vccd1 _0287_ sky130_fd_sc_hd__o21a_1
X_5374_ _0676_ _0593_ _0611_ _0599_ _1877_ vssd1 vssd1 vccd1 vccd1 _1878_ sky130_fd_sc_hd__o221a_1
X_4325_ egd_top.BitStream_buffer.BS_buffer\[80\] vssd1 vssd1 vccd1 vccd1 _0837_ sky130_fd_sc_hd__clkbuf_4
XFILLER_86_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4256_ _0767_ _3299_ _0768_ vssd1 vssd1 vccd1 vccd1 _0769_ sky130_fd_sc_hd__o21ai_1
X_4187_ _0532_ _0530_ _0524_ _0533_ vssd1 vssd1 vccd1 vccd1 _0700_ sky130_fd_sc_hd__o22a_1
XFILLER_74_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_386 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6828_ net72 _0287_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BitStream_buffer_output\[5\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_23_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_0__2887_ _2887_ vssd1 vssd1 vccd1 vccd1 clknet_0__2887_ sky130_fd_sc_hd__clkbuf_16
X_6759_ net163 _0218_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[61\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_12_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5090_ _2980_ _3123_ _1595_ vssd1 vssd1 vccd1 vccd1 _1596_ sky130_fd_sc_hd__o21ai_1
X_4110_ _0622_ _0623_ vssd1 vssd1 vccd1 vccd1 _0624_ sky130_fd_sc_hd__nand2_1
X_4041_ _2932_ _3211_ _3034_ vssd1 vssd1 vccd1 vccd1 _0555_ sky130_fd_sc_hd__and3_1
XFILLER_56_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6560__103 clknet_1_1__leaf__2887_ vssd1 vssd1 vccd1 vccd1 net137 sky130_fd_sc_hd__inv_2
X_5992_ _2982_ _2465_ _2458_ _2469_ vssd1 vssd1 vccd1 vccd1 _0261_ sky130_fd_sc_hd__o211a_1
X_4943_ _3167_ egd_top.BitStream_buffer.BS_buffer\[118\] vssd1 vssd1 vccd1 vccd1 _1451_
+ sky130_fd_sc_hd__nand2_1
XFILLER_32_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4874_ _0496_ _0527_ vssd1 vssd1 vccd1 vccd1 _1382_ sky130_fd_sc_hd__nand2_1
X_6613_ clknet_1_1__leaf__2883_ vssd1 vssd1 vccd1 vccd1 _2892_ sky130_fd_sc_hd__buf_1
XFILLER_32_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3825_ _0338_ vssd1 vssd1 vccd1 vccd1 _0339_ sky130_fd_sc_hd__buf_2
X_3756_ _3289_ vssd1 vssd1 vccd1 vccd1 _3290_ sky130_fd_sc_hd__buf_4
X_6475_ _2807_ _2771_ _2804_ vssd1 vssd1 vccd1 vccd1 _2838_ sky130_fd_sc_hd__nand3_1
X_5426_ _0566_ _3137_ _0568_ _3141_ _1929_ vssd1 vssd1 vccd1 vccd1 _1930_ sky130_fd_sc_hd__a221oi_1
X_3687_ egd_top.BitStream_buffer.BS_buffer\[70\] vssd1 vssd1 vccd1 vccd1 _3221_ sky130_fd_sc_hd__clkbuf_4
X_5357_ _0633_ _0523_ _1084_ _0526_ _1860_ vssd1 vssd1 vccd1 vccd1 _1861_ sky130_fd_sc_hd__o221a_1
XFILLER_87_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4308_ _3181_ _0623_ _0741_ _3176_ vssd1 vssd1 vccd1 vccd1 _0820_ sky130_fd_sc_hd__a22o_1
XFILLER_59_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5288_ _0406_ _0436_ vssd1 vssd1 vccd1 vccd1 _1793_ sky130_fd_sc_hd__nand2_1
XFILLER_59_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4239_ _3239_ vssd1 vssd1 vccd1 vccd1 _0752_ sky130_fd_sc_hd__inv_2
XFILLER_74_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3610_ _3143_ vssd1 vssd1 vccd1 vccd1 _3144_ sky130_fd_sc_hd__buf_2
X_4590_ _0474_ _0449_ _1097_ _1098_ _1099_ vssd1 vssd1 vccd1 vccd1 _1100_ sky130_fd_sc_hd__o2111a_1
X_3541_ egd_top.BitStream_buffer.BS_buffer\[110\] vssd1 vssd1 vccd1 vccd1 _3075_ sky130_fd_sc_hd__clkbuf_4
X_3472_ net11 vssd1 vssd1 vccd1 vccd1 _3011_ sky130_fd_sc_hd__buf_4
X_6260_ egd_top.BitStream_buffer.BitStream_buffer_output\[11\] vssd1 vssd1 vccd1 vccd1
+ _2631_ sky130_fd_sc_hd__inv_2
XFILLER_50_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5211_ _0804_ _3055_ _1713_ _1714_ _1715_ vssd1 vssd1 vccd1 vccd1 _1716_ sky130_fd_sc_hd__o2111a_1
X_6191_ _2586_ _2575_ vssd1 vssd1 vccd1 vccd1 _2589_ sky130_fd_sc_hd__and2_1
X_5142_ _0393_ _0342_ _0345_ _0400_ _1647_ vssd1 vssd1 vccd1 vccd1 _1648_ sky130_fd_sc_hd__a221oi_1
XFILLER_69_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5073_ _3293_ _3271_ _3315_ _3275_ _1579_ vssd1 vssd1 vccd1 vccd1 _1580_ sky130_fd_sc_hd__a221oi_1
X_4024_ _0488_ _3077_ vssd1 vssd1 vccd1 vccd1 _0538_ sky130_fd_sc_hd__nor2_2
XFILLER_56_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5975_ _2449_ _0676_ vssd1 vssd1 vccd1 vccd1 _2459_ sky130_fd_sc_hd__nand2_1
X_4926_ _1430_ _3239_ _1431_ _1432_ _1433_ vssd1 vssd1 vccd1 vccd1 _1434_ sky130_fd_sc_hd__o2111a_1
X_4857_ _0564_ _0583_ vssd1 vssd1 vccd1 vccd1 _1365_ sky130_fd_sc_hd__nand2_1
XFILLER_20_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3808_ _3290_ _3079_ vssd1 vssd1 vccd1 vccd1 _0322_ sky130_fd_sc_hd__nor2_2
XFILLER_60_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4788_ egd_top.BitStream_buffer.BS_buffer\[66\] vssd1 vssd1 vccd1 vccd1 _1297_ sky130_fd_sc_hd__clkinv_2
X_3739_ _3071_ _3213_ vssd1 vssd1 vccd1 vccd1 _3273_ sky130_fd_sc_hd__nand2_1
XFILLER_69_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6458_ _2819_ _2821_ vssd1 vssd1 vccd1 vccd1 _2822_ sky130_fd_sc_hd__nor2_1
X_6389_ _2757_ _2758_ _2664_ vssd1 vssd1 vccd1 vccd1 _2759_ sky130_fd_sc_hd__a21o_1
X_5409_ _1899_ _1912_ vssd1 vssd1 vccd1 vccd1 _1913_ sky130_fd_sc_hd__nand2_1
XFILLER_87_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5760_ _3138_ _0726_ _3173_ _3081_ _2260_ vssd1 vssd1 vccd1 vccd1 _2261_ sky130_fd_sc_hd__a221oi_1
X_4711_ _3049_ _0327_ _1219_ vssd1 vssd1 vccd1 vccd1 _1220_ sky130_fd_sc_hd__o21ai_1
X_5691_ _0960_ _0349_ _2191_ vssd1 vssd1 vccd1 vccd1 _2192_ sky130_fd_sc_hd__o21ai_1
X_4642_ _3283_ _3251_ _3276_ _3255_ _1151_ vssd1 vssd1 vccd1 vccd1 _1152_ sky130_fd_sc_hd__a221oi_1
X_4573_ _0375_ _0341_ _0344_ _0379_ _1082_ vssd1 vssd1 vccd1 vccd1 _1083_ sky130_fd_sc_hd__a221oi_1
X_3524_ _3057_ _3031_ _3032_ vssd1 vssd1 vccd1 vccd1 _3058_ sky130_fd_sc_hd__and3_2
X_6312_ _2676_ _2682_ vssd1 vssd1 vccd1 vccd1 _2683_ sky130_fd_sc_hd__nand2_1
X_3455_ net15 vssd1 vssd1 vccd1 vccd1 _2998_ sky130_fd_sc_hd__clkbuf_4
X_6243_ _2608_ _1003_ vssd1 vssd1 vccd1 vccd1 _2618_ sky130_fd_sc_hd__nand2_1
XFILLER_69_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3386_ _2938_ _2939_ egd_top.BitStream_buffer.buffer_index\[6\] vssd1 vssd1 vccd1
+ vccd1 _2940_ sky130_fd_sc_hd__and3_1
X_6174_ _3023_ _2555_ _2570_ _2574_ vssd1 vssd1 vccd1 vccd1 _0184_ sky130_fd_sc_hd__o211a_1
X_5125_ _0776_ _3299_ _1630_ vssd1 vssd1 vccd1 vccd1 _1631_ sky130_fd_sc_hd__o21ai_1
XFILLER_84_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5056_ _0796_ _0327_ _1560_ _1561_ _1562_ vssd1 vssd1 vccd1 vccd1 _1563_ sky130_fd_sc_hd__o2111ai_1
X_4007_ _0484_ _3031_ egd_top.BitStream_buffer.pc\[3\] vssd1 vssd1 vccd1 vccd1 _0521_
+ sky130_fd_sc_hd__and3_1
XFILLER_37_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5958_ _2449_ _0682_ vssd1 vssd1 vccd1 vccd1 _2450_ sky130_fd_sc_hd__nand2_1
X_4909_ _0727_ _3089_ _1414_ _1415_ _1416_ vssd1 vssd1 vccd1 vccd1 _1417_ sky130_fd_sc_hd__o2111a_1
XFILLER_21_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5889_ _0442_ _3230_ vssd1 vssd1 vccd1 vccd1 _2389_ sky130_fd_sc_hd__nand2_1
XFILLER_4_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_5 _1065_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6861_ net105 _0320_ vssd1 vssd1 vccd1 vccd1 net33 sky130_fd_sc_hd__dfxtp_2
X_6792_ net36 _0251_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[28\]
+ sky130_fd_sc_hd__dfxtp_4
X_5812_ _0837_ _3233_ _3236_ _3302_ _2311_ vssd1 vssd1 vccd1 vccd1 _2312_ sky130_fd_sc_hd__a221oi_2
X_5743_ _0869_ _0538_ _0393_ _0541_ _2243_ vssd1 vssd1 vccd1 vccd1 _2244_ sky130_fd_sc_hd__a221oi_1
XFILLER_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5674_ _2986_ _3088_ vssd1 vssd1 vccd1 vccd1 _2176_ sky130_fd_sc_hd__or2_1
XFILLER_30_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4625_ _0543_ _0529_ _0907_ _0525_ vssd1 vssd1 vccd1 vccd1 _1135_ sky130_fd_sc_hd__o22a_1
X_4556_ _3147_ egd_top.BitStream_buffer.BS_buffer\[124\] vssd1 vssd1 vccd1 vccd1 _1067_
+ sky130_fd_sc_hd__nand2_1
X_3507_ _3035_ vssd1 vssd1 vccd1 vccd1 _3041_ sky130_fd_sc_hd__buf_4
XFILLER_89_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4487_ _0365_ _0538_ egd_top.BitStream_buffer.BS_buffer\[34\] _0541_ _0997_ vssd1
+ vssd1 vccd1 vccd1 _0998_ sky130_fd_sc_hd__a221oi_1
X_3438_ net4 vssd1 vssd1 vccd1 vccd1 _2985_ sky130_fd_sc_hd__buf_4
X_6226_ _2608_ _1158_ vssd1 vssd1 vccd1 vccd1 _2609_ sky130_fd_sc_hd__nand2_1
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3369_ net17 vssd1 vssd1 vccd1 vccd1 _2923_ sky130_fd_sc_hd__clkinv_4
X_6157_ _2998_ _2554_ _2558_ _2565_ vssd1 vssd1 vccd1 vccd1 _0192_ sky130_fd_sc_hd__o211a_1
X_5108_ _0673_ _3183_ _1613_ vssd1 vssd1 vccd1 vccd1 _1614_ sky130_fd_sc_hd__o21ai_1
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6088_ _2517_ _0448_ vssd1 vssd1 vccd1 vccd1 _2525_ sky130_fd_sc_hd__nand2_1
X_5039_ _3177_ _3194_ _3197_ _0741_ _1545_ vssd1 vssd1 vccd1 vccd1 _1546_ sky130_fd_sc_hd__a221oi_1
XFILLER_72_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput31 net31 vssd1 vssd1 vccd1 vccd1 la_data_out_30_27[0] sky130_fd_sc_hd__buf_12
Xoutput20 net20 vssd1 vssd1 vccd1 vccd1 la_data_out_23_16[0] sky130_fd_sc_hd__buf_12
XFILLER_88_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1__f__2884_ clknet_0__2884_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__2884_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_48_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4410_ egd_top.BitStream_buffer.BS_buffer\[17\] vssd1 vssd1 vccd1 vccd1 _0922_ sky130_fd_sc_hd__inv_2
X_5390_ _0854_ _3319_ vssd1 vssd1 vccd1 vccd1 _1894_ sky130_fd_sc_hd__or2_1
X_4341_ _0330_ _3324_ _3326_ _0785_ _0852_ vssd1 vssd1 vccd1 vccd1 _0853_ sky130_fd_sc_hd__a221oi_1
X_4272_ egd_top.BitStream_buffer.BS_buffer\[93\] vssd1 vssd1 vccd1 vccd1 _0785_ sky130_fd_sc_hd__clkbuf_4
X_6011_ _2471_ _0524_ vssd1 vssd1 vccd1 vccd1 _2480_ sky130_fd_sc_hd__nand2_1
XTAP_189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6844_ net88 _0303_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[122\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_50_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3987_ egd_top.BitStream_buffer.BS_buffer\[16\] _0487_ egd_top.BitStream_buffer.BS_buffer\[17\]
+ _0490_ _0500_ vssd1 vssd1 vccd1 vccd1 _0501_ sky130_fd_sc_hd__a221oi_1
XFILLER_10_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6775_ net179 _0234_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[45\]
+ sky130_fd_sc_hd__dfxtp_1
X_5726_ _0685_ _0598_ vssd1 vssd1 vccd1 vccd1 _2227_ sky130_fd_sc_hd__or2_1
X_6529__75 clknet_1_1__leaf__2884_ vssd1 vssd1 vccd1 vccd1 net109 sky130_fd_sc_hd__inv_2
X_5657_ _0566_ _3144_ _0568_ _3148_ _2158_ vssd1 vssd1 vccd1 vccd1 _2159_ sky130_fd_sc_hd__a221oi_1
X_4608_ _0581_ egd_top.BitStream_buffer.BS_buffer\[14\] vssd1 vssd1 vccd1 vccd1 _1118_
+ sky130_fd_sc_hd__nand2_1
XFILLER_2_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6544__89 clknet_1_0__leaf__2885_ vssd1 vssd1 vccd1 vccd1 net123 sky130_fd_sc_hd__inv_2
X_5588_ _0457_ _3221_ vssd1 vssd1 vccd1 vccd1 _2090_ sky130_fd_sc_hd__nand2_1
X_4539_ _3250_ egd_top.BitStream_buffer.BS_buffer\[77\] vssd1 vssd1 vccd1 vccd1 _1050_
+ sky130_fd_sc_hd__nand2_1
XFILLER_89_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6209_ _2902_ egd_top.BitStream_buffer.pc\[1\] vssd1 vssd1 vccd1 vccd1 _2598_ sky130_fd_sc_hd__nand2_1
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3910_ _3033_ _2934_ vssd1 vssd1 vccd1 vccd1 _0424_ sky130_fd_sc_hd__nand2_1
XFILLER_32_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4890_ _3291_ egd_top.BitStream_buffer.BS_buffer\[88\] vssd1 vssd1 vccd1 vccd1 _1398_
+ sky130_fd_sc_hd__nand2_1
X_3841_ _0353_ _0354_ vssd1 vssd1 vccd1 vccd1 _0355_ sky130_fd_sc_hd__nand2_1
XFILLER_80_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3772_ egd_top.BitStream_buffer.BS_buffer\[87\] vssd1 vssd1 vccd1 vccd1 _3306_ sky130_fd_sc_hd__clkinv_2
X_5511_ _0642_ _0342_ _0345_ _0874_ _2013_ vssd1 vssd1 vccd1 vccd1 _2014_ sky130_fd_sc_hd__a221oi_1
X_6491_ _2840_ _2805_ vssd1 vssd1 vccd1 vccd1 _2853_ sky130_fd_sc_hd__nor2_1
X_5442_ _1945_ _3027_ _2905_ vssd1 vssd1 vccd1 vccd1 _1946_ sky130_fd_sc_hd__a21oi_1
X_5373_ _0574_ _0596_ vssd1 vssd1 vccd1 vccd1 _1877_ sky130_fd_sc_hd__or2_1
X_4324_ _3268_ _3251_ _3272_ _3255_ _0835_ vssd1 vssd1 vccd1 vccd1 _0836_ sky130_fd_sc_hd__a221oi_1
XFILLER_59_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4255_ _3301_ _3288_ vssd1 vssd1 vccd1 vccd1 _0768_ sky130_fd_sc_hd__nand2_1
X_4186_ egd_top.BitStream_buffer.BS_buffer\[28\] vssd1 vssd1 vccd1 vccd1 _0699_ sky130_fd_sc_hd__inv_2
XFILLER_67_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6827_ net71 _0286_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BitStream_buffer_output\[4\]
+ sky130_fd_sc_hd__dfxtp_2
Xclkbuf_0__2886_ _2886_ vssd1 vssd1 vccd1 vccd1 clknet_0__2886_ sky130_fd_sc_hd__clkbuf_16
X_6758_ net162 _0217_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[62\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_10_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5709_ _0755_ _0464_ _2207_ _2208_ _2209_ vssd1 vssd1 vccd1 vccd1 _2210_ sky130_fd_sc_hd__o2111a_1
XFILLER_12_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_104 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4040_ _0553_ vssd1 vssd1 vccd1 vccd1 _0554_ sky130_fd_sc_hd__inv_2
XFILLER_1_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5991_ _2466_ _0492_ vssd1 vssd1 vccd1 vccd1 _2469_ sky130_fd_sc_hd__nand2_1
XFILLER_24_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4942_ _3155_ egd_top.BitStream_buffer.BS_buffer\[120\] vssd1 vssd1 vccd1 vccd1 _1450_
+ sky130_fd_sc_hd__nand2_1
XFILLER_52_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4873_ _0489_ _0509_ vssd1 vssd1 vccd1 vccd1 _1381_ sky130_fd_sc_hd__nand2_1
XFILLER_20_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3824_ _2932_ _3211_ egd_top.BitStream_buffer.pc\[5\] vssd1 vssd1 vccd1 vccd1 _0338_
+ sky130_fd_sc_hd__and3_2
X_3755_ egd_top.BitStream_buffer.pc\[5\] _2932_ _3211_ vssd1 vssd1 vccd1 vccd1 _3289_
+ sky130_fd_sc_hd__or3_2
X_3686_ _3219_ vssd1 vssd1 vccd1 vccd1 _3220_ sky130_fd_sc_hd__clkbuf_4
X_6474_ _2835_ _2836_ vssd1 vssd1 vccd1 vccd1 _2837_ sky130_fd_sc_hd__nand2_1
X_5425_ _0591_ _3145_ _1928_ vssd1 vssd1 vccd1 vccd1 _1929_ sky130_fd_sc_hd__o21ai_1
X_5356_ _0865_ _0530_ _0940_ _0534_ vssd1 vssd1 vccd1 vccd1 _1860_ sky130_fd_sc_hd__o22a_1
XFILLER_58_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4307_ _3204_ _3156_ _0746_ _3160_ _0818_ vssd1 vssd1 vccd1 vccd1 _0819_ sky130_fd_sc_hd__a221oi_1
X_5287_ _1790_ _1791_ vssd1 vssd1 vccd1 vccd1 _1792_ sky130_fd_sc_hd__nor2_1
XFILLER_59_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4238_ egd_top.BitStream_buffer.BS_buffer\[65\] vssd1 vssd1 vccd1 vccd1 _0751_ sky130_fd_sc_hd__clkbuf_4
X_6683__55 clknet_1_1__leaf__2898_ vssd1 vssd1 vccd1 vccd1 net89 sky130_fd_sc_hd__inv_2
X_4169_ egd_top.BitStream_buffer.BS_buffer\[4\] vssd1 vssd1 vccd1 vccd1 _0682_ sky130_fd_sc_hd__inv_2
XFILLER_70_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_479 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3540_ _3073_ vssd1 vssd1 vccd1 vccd1 _3074_ sky130_fd_sc_hd__buf_4
X_5210_ _3047_ _3109_ vssd1 vssd1 vccd1 vccd1 _1715_ sky130_fd_sc_hd__nand2_1
X_3471_ _3008_ _2976_ _3002_ _3010_ vssd1 vssd1 vccd1 vccd1 _0303_ sky130_fd_sc_hd__o211a_1
XFILLER_89_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6190_ _2588_ vssd1 vssd1 vccd1 vccd1 _0183_ sky130_fd_sc_hd__inv_2
XFILLER_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5141_ _0401_ _0350_ _1646_ vssd1 vssd1 vccd1 vccd1 _1647_ sky130_fd_sc_hd__o21ai_1
X_5072_ _0771_ _3279_ _1578_ vssd1 vssd1 vccd1 vccd1 _1579_ sky130_fd_sc_hd__o21ai_1
X_4023_ egd_top.BitStream_buffer.BS_buffer\[30\] vssd1 vssd1 vccd1 vccd1 _0537_ sky130_fd_sc_hd__clkbuf_4
XFILLER_56_107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5974_ _2901_ vssd1 vssd1 vccd1 vccd1 _2458_ sky130_fd_sc_hd__buf_2
XFILLER_52_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4925_ _3235_ _3264_ vssd1 vssd1 vccd1 vccd1 _1433_ sky130_fd_sc_hd__nand2_1
XFILLER_40_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4856_ _1351_ _1355_ _1359_ _1363_ vssd1 vssd1 vccd1 vccd1 _1364_ sky130_fd_sc_hd__and4_1
XFILLER_20_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3807_ egd_top.BitStream_buffer.BS_buffer\[95\] vssd1 vssd1 vccd1 vccd1 _3341_ sky130_fd_sc_hd__clkbuf_4
X_4787_ _1294_ _1295_ vssd1 vssd1 vccd1 vccd1 _1296_ sky130_fd_sc_hd__nor2_1
X_3738_ egd_top.BitStream_buffer.BS_buffer\[77\] vssd1 vssd1 vccd1 vccd1 _3272_ sky130_fd_sc_hd__clkbuf_4
X_3669_ _3202_ vssd1 vssd1 vccd1 vccd1 _3203_ sky130_fd_sc_hd__buf_2
XFILLER_69_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6457_ _2818_ _2820_ _2701_ _2737_ vssd1 vssd1 vccd1 vccd1 _2821_ sky130_fd_sc_hd__a31o_1
X_6388_ _2713_ egd_top.BitStream_buffer.BitStream_buffer_output\[11\] vssd1 vssd1
+ vccd1 vccd1 _2758_ sky130_fd_sc_hd__nand2_1
X_5408_ _1902_ _1905_ _1908_ _1911_ vssd1 vssd1 vccd1 vccd1 _1912_ sky130_fd_sc_hd__and4_1
X_5339_ _0650_ _0425_ vssd1 vssd1 vccd1 vccd1 _1843_ sky130_fd_sc_hd__or2_1
XFILLER_85_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6647__22 clknet_1_0__leaf__2895_ vssd1 vssd1 vccd1 vccd1 net56 sky130_fd_sc_hd__inv_2
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6662__36 clknet_1_0__leaf__2896_ vssd1 vssd1 vccd1 vccd1 net70 sky130_fd_sc_hd__inv_2
XFILLER_74_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4710_ _0329_ _3040_ vssd1 vssd1 vccd1 vccd1 _1219_ sky130_fd_sc_hd__nand2_1
X_5690_ _0352_ _0416_ vssd1 vssd1 vccd1 vccd1 _2191_ sky130_fd_sc_hd__nand2_1
X_4641_ _1149_ _3260_ _1150_ vssd1 vssd1 vccd1 vccd1 _1151_ sky130_fd_sc_hd__o21ai_1
X_4572_ _0383_ _0349_ _1081_ vssd1 vssd1 vccd1 vccd1 _1082_ sky130_fd_sc_hd__o21ai_1
X_3523_ _2930_ vssd1 vssd1 vccd1 vccd1 _3057_ sky130_fd_sc_hd__inv_2
X_6311_ _2680_ _2681_ vssd1 vssd1 vccd1 vccd1 _2682_ sky130_fd_sc_hd__nand2_1
X_3454_ _2995_ _2975_ _2913_ _2997_ vssd1 vssd1 vccd1 vccd1 _0307_ sky130_fd_sc_hd__o211a_1
X_6242_ _3011_ _2603_ _2611_ _2617_ vssd1 vssd1 vccd1 vccd1 _0165_ sky130_fd_sc_hd__o211a_1
X_3385_ egd_top.BitStream_buffer.buffer_index\[4\] vssd1 vssd1 vccd1 vccd1 _2939_
+ sky130_fd_sc_hd__inv_2
X_6173_ _2553_ _1035_ vssd1 vssd1 vccd1 vccd1 _2574_ sky130_fd_sc_hd__nand2_1
XFILLER_69_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5124_ _3301_ _0780_ vssd1 vssd1 vccd1 vccd1 _1630_ sky130_fd_sc_hd__nand2_1
XFILLER_57_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5055_ _3340_ _0716_ vssd1 vssd1 vccd1 vccd1 _1562_ sky130_fd_sc_hd__nand2_1
X_4006_ _0519_ vssd1 vssd1 vccd1 vccd1 _0520_ sky130_fd_sc_hd__inv_2
X_5957_ _2441_ vssd1 vssd1 vccd1 vccd1 _2449_ sky130_fd_sc_hd__buf_2
X_4908_ _0804_ _3105_ vssd1 vssd1 vccd1 vccd1 _1416_ sky130_fd_sc_hd__or2_1
XFILLER_33_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5888_ _3244_ _0415_ _0751_ _0419_ _2387_ vssd1 vssd1 vccd1 vccd1 _2388_ sky130_fd_sc_hd__a221oi_1
X_4839_ _0412_ _0396_ _0399_ _0416_ _1346_ vssd1 vssd1 vccd1 vccd1 _1347_ sky130_fd_sc_hd__a221oi_1
X_6509_ _2868_ _2701_ _2870_ vssd1 vssd1 vccd1 vccd1 _2871_ sky130_fd_sc_hd__nand3_1
XFILLER_4_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6621__159 clknet_1_1__leaf__2892_ vssd1 vssd1 vccd1 vccd1 net193 sky130_fd_sc_hd__inv_2
XFILLER_24_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_6 _1111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_471 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6860_ net104 _0319_ vssd1 vssd1 vccd1 vccd1 net32 sky130_fd_sc_hd__dfxtp_2
XFILLER_19_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6791_ net195 _0250_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[29\]
+ sky130_fd_sc_hd__dfxtp_4
X_5811_ _3277_ _3240_ _2310_ vssd1 vssd1 vccd1 vccd1 _2311_ sky130_fd_sc_hd__o21ai_1
X_5742_ _0936_ _0545_ _2242_ vssd1 vssd1 vccd1 vccd1 _2243_ sky130_fd_sc_hd__o21ai_1
X_6596__136 clknet_1_0__leaf__2890_ vssd1 vssd1 vccd1 vccd1 net170 sky130_fd_sc_hd__inv_2
XFILLER_22_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5673_ _3093_ _3169_ vssd1 vssd1 vccd1 vccd1 _2175_ sky130_fd_sc_hd__nand2_1
XFILLER_30_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4624_ _0519_ _0504_ _0527_ _0508_ _1133_ vssd1 vssd1 vccd1 vccd1 _1134_ sky130_fd_sc_hd__a221oi_1
X_4555_ _3140_ _0741_ vssd1 vssd1 vccd1 vccd1 _1066_ sky130_fd_sc_hd__nand2_1
X_3506_ egd_top.BitStream_buffer.BS_buffer\[97\] vssd1 vssd1 vccd1 vccd1 _3040_ sky130_fd_sc_hd__clkbuf_4
X_4486_ _0995_ _0545_ _0996_ vssd1 vssd1 vccd1 vccd1 _0997_ sky130_fd_sc_hd__o21ai_1
X_3437_ _2982_ _2975_ _2913_ _2984_ vssd1 vssd1 vccd1 vccd1 _0311_ sky130_fd_sc_hd__o211a_1
X_6225_ _2601_ vssd1 vssd1 vccd1 vccd1 _2608_ sky130_fd_sc_hd__buf_2
XFILLER_85_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3368_ net18 vssd1 vssd1 vccd1 vccd1 _2922_ sky130_fd_sc_hd__inv_2
X_6156_ _2561_ _3085_ vssd1 vssd1 vccd1 vccd1 _2565_ sky130_fd_sc_hd__nand2_1
X_5107_ _3186_ _0553_ vssd1 vssd1 vccd1 vccd1 _1613_ sky130_fd_sc_hd__nand2_1
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6087_ _3008_ _2511_ _2516_ _2524_ vssd1 vssd1 vccd1 vccd1 _0221_ sky130_fd_sc_hd__o211a_1
X_5038_ _3015_ _3200_ _1544_ vssd1 vssd1 vccd1 vccd1 _1545_ sky130_fd_sc_hd__o21ai_1
XFILLER_72_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6641__17 clknet_1_1__leaf__2894_ vssd1 vssd1 vccd1 vccd1 net51 sky130_fd_sc_hd__inv_2
XFILLER_38_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput32 net32 vssd1 vssd1 vccd1 vccd1 la_data_out_30_27[1] sky130_fd_sc_hd__buf_12
Xoutput21 net21 vssd1 vssd1 vccd1 vccd1 la_data_out_23_16[1] sky130_fd_sc_hd__buf_12
XFILLER_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__2883_ clknet_0__2883_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__2883_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_76_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4340_ _0850_ _3330_ _0851_ vssd1 vssd1 vccd1 vccd1 _0852_ sky130_fd_sc_hd__o21ai_1
X_4271_ egd_top.BitStream_buffer.BS_buffer\[94\] vssd1 vssd1 vccd1 vccd1 _0784_ sky130_fd_sc_hd__clkinv_2
XFILLER_67_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6010_ _3008_ _2466_ _2474_ _2479_ vssd1 vssd1 vccd1 vccd1 _0253_ sky130_fd_sc_hd__o211a_1
XFILLER_79_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6843_ net87 _0302_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[123\]
+ sky130_fd_sc_hd__dfxtp_2
X_6604__143 clknet_1_0__leaf__2891_ vssd1 vssd1 vccd1 vccd1 net177 sky130_fd_sc_hd__inv_2
XFILLER_62_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3986_ _0492_ _0495_ _0499_ vssd1 vssd1 vccd1 vccd1 _0500_ sky130_fd_sc_hd__o21ai_1
X_6774_ net178 _0233_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[46\]
+ sky130_fd_sc_hd__dfxtp_2
X_5725_ _0520_ _0575_ _2223_ _2224_ _2225_ vssd1 vssd1 vccd1 vccd1 _2226_ sky130_fd_sc_hd__o2111a_1
XFILLER_22_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5656_ _0562_ _3137_ _3141_ _0553_ vssd1 vssd1 vccd1 vccd1 _2158_ sky130_fd_sc_hd__a22o_1
X_4607_ _0577_ egd_top.BitStream_buffer.BS_buffer\[12\] vssd1 vssd1 vccd1 vccd1 _1117_
+ sky130_fd_sc_hd__nand2_1
X_5587_ _0452_ _3210_ vssd1 vssd1 vccd1 vccd1 _2089_ sky130_fd_sc_hd__nand2_1
XFILLER_89_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4538_ _3254_ egd_top.BitStream_buffer.BS_buffer\[78\] vssd1 vssd1 vccd1 vccd1 _1049_
+ sky130_fd_sc_hd__nand2_1
X_4469_ _0569_ _0592_ _0682_ _0596_ _0979_ vssd1 vssd1 vccd1 vccd1 _0980_ sky130_fd_sc_hd__o221a_1
XFILLER_77_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6208_ _2925_ _2578_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.pc\[1\] sky130_fd_sc_hd__xor2_4
XFILLER_58_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6139_ _2553_ vssd1 vssd1 vccd1 vccd1 _2555_ sky130_fd_sc_hd__buf_2
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6689__61 clknet_1_1__leaf__2898_ vssd1 vssd1 vccd1 vccd1 net95 sky130_fd_sc_hd__inv_2
XFILLER_3_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3840_ egd_top.BitStream_buffer.BS_buffer\[38\] vssd1 vssd1 vccd1 vccd1 _0354_ sky130_fd_sc_hd__clkbuf_4
XFILLER_32_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3771_ _3288_ _3292_ _3293_ _3295_ _3304_ vssd1 vssd1 vccd1 vccd1 _3305_ sky130_fd_sc_hd__a221oi_1
X_5510_ _0659_ _0350_ _2012_ vssd1 vssd1 vccd1 vccd1 _2013_ sky130_fd_sc_hd__o21ai_1
XFILLER_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6490_ _2828_ _2823_ _2847_ vssd1 vssd1 vccd1 vccd1 _2852_ sky130_fd_sc_hd__nand3_1
X_5441_ egd_top.BitStream_buffer.BitStream_buffer_output\[5\] vssd1 vssd1 vccd1 vccd1
+ _1945_ sky130_fd_sc_hd__inv_2
X_5372_ _0986_ _0576_ _1873_ _1874_ _1875_ vssd1 vssd1 vccd1 vccd1 _1876_ sky130_fd_sc_hd__o2111a_1
X_4323_ _0833_ _3260_ _0834_ vssd1 vssd1 vccd1 vccd1 _0835_ sky130_fd_sc_hd__o21ai_1
XFILLER_86_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4254_ egd_top.BitStream_buffer.BS_buffer\[81\] vssd1 vssd1 vccd1 vccd1 _0767_ sky130_fd_sc_hd__clkinv_2
X_4185_ _0505_ _0504_ _0515_ _0508_ _0697_ vssd1 vssd1 vccd1 vccd1 _0698_ sky130_fd_sc_hd__a221oi_1
XFILLER_67_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_506 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__2885_ _2885_ vssd1 vssd1 vccd1 vccd1 clknet_0__2885_ sky130_fd_sc_hd__clkbuf_16
X_6826_ net70 _0285_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BitStream_buffer_output\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_23_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6757_ net161 _0216_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[63\]
+ sky130_fd_sc_hd__dfxtp_1
X_3969_ _0411_ _0482_ vssd1 vssd1 vccd1 vccd1 _0483_ sky130_fd_sc_hd__nand2_1
X_5708_ _3257_ _0449_ vssd1 vssd1 vccd1 vccd1 _2209_ sky130_fd_sc_hd__or2_1
XFILLER_50_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5639_ _0329_ _3128_ vssd1 vssd1 vccd1 vccd1 _2141_ sky130_fd_sc_hd__nand2_1
XFILLER_88_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5990_ _2979_ _2465_ _2458_ _2468_ vssd1 vssd1 vccd1 vccd1 _0262_ sky130_fd_sc_hd__o211a_1
X_4941_ _3159_ egd_top.BitStream_buffer.BS_buffer\[121\] vssd1 vssd1 vccd1 vccd1 _1449_
+ sky130_fd_sc_hd__nand2_1
X_4872_ _0486_ _0515_ vssd1 vssd1 vccd1 vccd1 _1380_ sky130_fd_sc_hd__nand2_1
XFILLER_17_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3823_ egd_top.BitStream_buffer.BS_buffer\[36\] vssd1 vssd1 vccd1 vccd1 _0337_ sky130_fd_sc_hd__clkbuf_4
XFILLER_20_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3754_ egd_top.BitStream_buffer.BS_buffer\[82\] vssd1 vssd1 vccd1 vccd1 _3288_ sky130_fd_sc_hd__clkbuf_4
XFILLER_9_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3685_ _3218_ vssd1 vssd1 vccd1 vccd1 _3219_ sky130_fd_sc_hd__inv_2
X_6473_ _2820_ _2818_ _2701_ vssd1 vssd1 vccd1 vccd1 _2836_ sky130_fd_sc_hd__o21ai_1
X_5424_ _3148_ _1076_ vssd1 vssd1 vccd1 vccd1 _1928_ sky130_fd_sc_hd__nand2_1
X_5355_ _0537_ _0504_ _0540_ _0508_ _1858_ vssd1 vssd1 vccd1 vccd1 _1859_ sky130_fd_sc_hd__a221oi_1
XFILLER_58_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4306_ _0816_ _0817_ vssd1 vssd1 vccd1 vccd1 _0818_ sky130_fd_sc_hd__nand2_1
X_5286_ _3087_ _0874_ _0339_ _0642_ _0352_ vssd1 vssd1 vccd1 vccd1 _1791_ sky130_fd_sc_hd__a32o_1
X_4237_ _0733_ _0749_ vssd1 vssd1 vccd1 vccd1 _0750_ sky130_fd_sc_hd__nand2_1
XFILLER_4_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4168_ _0676_ _0576_ _0677_ _0678_ _0680_ vssd1 vssd1 vccd1 vccd1 _0681_ sky130_fd_sc_hd__o2111a_1
XFILLER_74_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4099_ _0612_ vssd1 vssd1 vccd1 vccd1 _0613_ sky130_fd_sc_hd__clkbuf_2
XFILLER_43_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6809_ net53 _0268_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[11\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_23_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3470_ _2989_ _3009_ vssd1 vssd1 vccd1 vccd1 _3010_ sky130_fd_sc_hd__nand2_1
XFILLER_69_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5140_ _0353_ _0407_ vssd1 vssd1 vccd1 vccd1 _1646_ sky130_fd_sc_hd__nand2_1
XFILLER_69_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5071_ _3282_ _0774_ vssd1 vssd1 vccd1 vccd1 _1578_ sky130_fd_sc_hd__nand2_1
X_4022_ _0520_ _0523_ _0524_ _0526_ _0535_ vssd1 vssd1 vccd1 vccd1 _0536_ sky130_fd_sc_hd__o221a_1
XFILLER_84_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5973_ _3011_ _2443_ _2446_ _2457_ vssd1 vssd1 vccd1 vccd1 _0268_ sky130_fd_sc_hd__o211a_1
XFILLER_37_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4924_ _3232_ _3256_ vssd1 vssd1 vccd1 vccd1 _1432_ sky130_fd_sc_hd__nand2_1
XFILLER_40_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4855_ _3230_ _0470_ _3237_ _0473_ _1362_ vssd1 vssd1 vccd1 vccd1 _1363_ sky130_fd_sc_hd__a221oi_1
X_3806_ _3339_ vssd1 vssd1 vccd1 vccd1 _3340_ sky130_fd_sc_hd__clkbuf_4
XFILLER_20_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4786_ _3104_ _0459_ _2934_ _0461_ _0442_ vssd1 vssd1 vccd1 vccd1 _1295_ sky130_fd_sc_hd__a32o_1
X_3737_ _3270_ vssd1 vssd1 vccd1 vccd1 _3271_ sky130_fd_sc_hd__clkbuf_4
X_6525_ clknet_1_0__leaf__2883_ vssd1 vssd1 vccd1 vccd1 _2884_ sky130_fd_sc_hd__buf_1
X_3668_ _3201_ vssd1 vssd1 vccd1 vccd1 _3202_ sky130_fd_sc_hd__clkbuf_2
X_6456_ _2816_ vssd1 vssd1 vccd1 vccd1 _2820_ sky130_fd_sc_hd__inv_2
X_3599_ egd_top.BitStream_buffer.BS_buffer\[122\] vssd1 vssd1 vccd1 vccd1 _3133_ sky130_fd_sc_hd__buf_2
X_6387_ _2712_ _2631_ vssd1 vssd1 vccd1 vccd1 _2757_ sky130_fd_sc_hd__nand2_1
X_5407_ _3311_ _3271_ _0772_ _3275_ _1910_ vssd1 vssd1 vccd1 vccd1 _1911_ sky130_fd_sc_hd__a221oi_1
X_5338_ _1832_ _1835_ _1838_ _1841_ vssd1 vssd1 vccd1 vccd1 _1842_ sky130_fd_sc_hd__and4_1
XFILLER_87_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5269_ _0955_ _0439_ _1773_ vssd1 vssd1 vccd1 vccd1 _1774_ sky130_fd_sc_hd__o21ai_1
XFILLER_47_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_299 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4640_ _3263_ _3272_ vssd1 vssd1 vccd1 vccd1 _1150_ sky130_fd_sc_hd__nand2_1
X_4571_ _0352_ egd_top.BitStream_buffer.BS_buffer\[42\] vssd1 vssd1 vccd1 vccd1 _1081_
+ sky130_fd_sc_hd__nand2_1
X_6310_ _2677_ vssd1 vssd1 vccd1 vccd1 _2681_ sky130_fd_sc_hd__buf_6
X_3522_ _3055_ vssd1 vssd1 vccd1 vccd1 _3056_ sky130_fd_sc_hd__buf_2
X_3453_ _2989_ _2996_ vssd1 vssd1 vccd1 vccd1 _2997_ sky130_fd_sc_hd__nand2_1
X_6241_ _2608_ _0850_ vssd1 vssd1 vccd1 vccd1 _2617_ sky130_fd_sc_hd__nand2_1
X_6172_ _3020_ _2555_ _2570_ _2573_ vssd1 vssd1 vccd1 vccd1 _0185_ sky130_fd_sc_hd__o211a_1
X_3384_ egd_top.BitStream_buffer.buffer_index\[5\] vssd1 vssd1 vccd1 vccd1 _2938_
+ sky130_fd_sc_hd__inv_2
X_5123_ _1619_ _1622_ _1625_ _1628_ vssd1 vssd1 vccd1 vccd1 _1629_ sky130_fd_sc_hd__and4_1
X_5054_ _0329_ _3062_ vssd1 vssd1 vccd1 vccd1 _1561_ sky130_fd_sc_hd__nand2_1
XFILLER_72_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4005_ egd_top.BitStream_buffer.BS_buffer\[24\] vssd1 vssd1 vccd1 vccd1 _0519_ sky130_fd_sc_hd__clkbuf_4
X_6625__2 clknet_1_0__leaf__2893_ vssd1 vssd1 vccd1 vccd1 net36 sky130_fd_sc_hd__inv_2
XFILLER_65_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5956_ _2985_ _2442_ _2446_ _2448_ vssd1 vssd1 vccd1 vccd1 _0276_ sky130_fd_sc_hd__o211a_1
XFILLER_40_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4907_ _3098_ egd_top.BitStream_buffer.BS_buffer\[108\] vssd1 vssd1 vccd1 vccd1 _1415_
+ sky130_fd_sc_hd__nand2_1
X_5887_ _0474_ _0422_ _2386_ vssd1 vssd1 vccd1 vccd1 _2387_ sky130_fd_sc_hd__o21ai_1
X_4838_ _0437_ _0402_ _1345_ vssd1 vssd1 vccd1 vccd1 _1346_ sky130_fd_sc_hd__o21ai_1
X_6573__115 clknet_1_1__leaf__2888_ vssd1 vssd1 vccd1 vccd1 net149 sky130_fd_sc_hd__inv_2
X_4769_ _1276_ _0368_ _1277_ vssd1 vssd1 vccd1 vccd1 _1278_ sky130_fd_sc_hd__o21ai_1
X_6508_ _2819_ _2849_ _2869_ vssd1 vssd1 vccd1 vccd1 _2870_ sky130_fd_sc_hd__nand3_1
X_6439_ _2678_ _1705_ vssd1 vssd1 vccd1 vccd1 _2803_ sky130_fd_sc_hd__nand2_1
XFILLER_20_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_76 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_20 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_7 _1331_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6790_ net194 _0249_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[30\]
+ sky130_fd_sc_hd__dfxtp_1
X_5810_ _3243_ _3283_ vssd1 vssd1 vccd1 vccd1 _2310_ sky130_fd_sc_hd__nand2_1
X_5741_ _0547_ _0379_ vssd1 vssd1 vccd1 vccd1 _2242_ sky130_fd_sc_hd__nand2_1
XFILLER_15_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5672_ _3099_ _3153_ vssd1 vssd1 vccd1 vccd1 _2174_ sky130_fd_sc_hd__nand2_1
X_4623_ _0524_ _0512_ _1132_ vssd1 vssd1 vccd1 vccd1 _1133_ sky130_fd_sc_hd__o21ai_1
X_4554_ _1061_ _1062_ _1063_ _1064_ vssd1 vssd1 vccd1 vccd1 _1065_ sky130_fd_sc_hd__and4_1
X_3505_ _3038_ vssd1 vssd1 vccd1 vccd1 _3039_ sky130_fd_sc_hd__clkbuf_4
X_4485_ _0547_ _0540_ vssd1 vssd1 vccd1 vccd1 _0996_ sky130_fd_sc_hd__nand2_1
X_6224_ _2985_ _2602_ _2570_ _2607_ vssd1 vssd1 vccd1 vccd1 _0173_ sky130_fd_sc_hd__o211a_1
X_3436_ _2976_ _2983_ vssd1 vssd1 vccd1 vccd1 _2984_ sky130_fd_sc_hd__nand2_1
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3367_ egd_top.BitStream_buffer.pc\[1\] vssd1 vssd1 vccd1 vccd1 _2921_ sky130_fd_sc_hd__inv_2
X_6155_ _2995_ _2554_ _2558_ _2564_ vssd1 vssd1 vccd1 vccd1 _0193_ sky130_fd_sc_hd__o211a_1
X_5106_ _0741_ _3194_ _3197_ _3187_ _1611_ vssd1 vssd1 vccd1 vccd1 _1612_ sky130_fd_sc_hd__a221oi_1
XFILLER_85_534 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6086_ _2517_ _0650_ vssd1 vssd1 vccd1 vccd1 _2524_ sky130_fd_sc_hd__nand2_1
X_5037_ _3203_ _3138_ vssd1 vssd1 vccd1 vccd1 _1544_ sky130_fd_sc_hd__nand2_1
XFILLER_57_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5939_ _2436_ vssd1 vssd1 vccd1 vccd1 _0281_ sky130_fd_sc_hd__clkbuf_1
XFILLER_15_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput22 net22 vssd1 vssd1 vccd1 vccd1 la_data_out_23_16[2] sky130_fd_sc_hd__buf_12
Xoutput33 net33 vssd1 vssd1 vccd1 vccd1 la_data_out_30_27[2] sky130_fd_sc_hd__buf_12
XFILLER_88_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f__2882_ clknet_0__2882_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__2882_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_48_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4270_ _3327_ _3324_ _3326_ _0330_ _0782_ vssd1 vssd1 vccd1 vccd1 _0783_ sky130_fd_sc_hd__a221oi_1
XFILLER_86_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_504 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6842_ net86 _0301_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[124\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_50_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3985_ _0497_ _0498_ vssd1 vssd1 vccd1 vccd1 _0499_ sky130_fd_sc_hd__nand2_1
X_6773_ net177 _0232_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[47\]
+ sky130_fd_sc_hd__dfxtp_1
X_5724_ _1128_ _0587_ vssd1 vssd1 vccd1 vccd1 _2225_ sky130_fd_sc_hd__or2_1
XFILLER_10_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5655_ _2144_ _2156_ vssd1 vssd1 vccd1 vccd1 _2157_ sky130_fd_sc_hd__nand2_1
X_4606_ _0574_ _0558_ _1113_ _1114_ _1115_ vssd1 vssd1 vccd1 vccd1 _1116_ sky130_fd_sc_hd__o2111a_1
X_5586_ _0478_ _0414_ _0664_ _0418_ _2087_ vssd1 vssd1 vccd1 vccd1 _2088_ sky130_fd_sc_hd__a221oi_1
X_4537_ _3262_ egd_top.BitStream_buffer.BS_buffer\[76\] vssd1 vssd1 vccd1 vccd1 _1048_
+ sky130_fd_sc_hd__nand2_1
X_4468_ _0673_ _0598_ vssd1 vssd1 vccd1 vccd1 _0979_ sky130_fd_sc_hd__or2_1
XFILLER_89_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6207_ _2597_ vssd1 vssd1 vccd1 vccd1 _0179_ sky130_fd_sc_hd__inv_2
X_3419_ _2911_ _2968_ vssd1 vssd1 vccd1 vccd1 _2969_ sky130_fd_sc_hd__or2_1
X_4399_ _0900_ _0904_ _0906_ _0910_ vssd1 vssd1 vccd1 vccd1 _0911_ sky130_fd_sc_hd__and4_1
X_6138_ _2553_ vssd1 vssd1 vccd1 vccd1 _2554_ sky130_fd_sc_hd__buf_2
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6069_ _2982_ _2510_ _2501_ _2514_ vssd1 vssd1 vccd1 vccd1 _0229_ sky130_fd_sc_hd__o211a_1
XFILLER_26_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6579__121 clknet_1_0__leaf__2888_ vssd1 vssd1 vccd1 vccd1 net155 sky130_fd_sc_hd__inv_2
XFILLER_26_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_423 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3770_ _3296_ _3299_ _3303_ vssd1 vssd1 vccd1 vccd1 _3304_ sky130_fd_sc_hd__o21ai_1
XFILLER_12_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5440_ _1885_ _1942_ _1943_ vssd1 vssd1 vccd1 vccd1 _1944_ sky130_fd_sc_hd__nand3_1
XFILLER_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5371_ _0692_ _0588_ vssd1 vssd1 vccd1 vccd1 _1875_ sky130_fd_sc_hd__or2_1
X_6534__80 clknet_1_0__leaf__2884_ vssd1 vssd1 vccd1 vccd1 net114 sky130_fd_sc_hd__inv_2
X_4322_ _3263_ _3252_ vssd1 vssd1 vccd1 vccd1 _0834_ sky130_fd_sc_hd__nand2_1
X_4253_ _0754_ _0758_ _0762_ _0765_ vssd1 vssd1 vccd1 vccd1 _0766_ sky130_fd_sc_hd__and4_1
X_4184_ _0520_ _0512_ _0696_ vssd1 vssd1 vccd1 vccd1 _0697_ sky130_fd_sc_hd__o21ai_1
XFILLER_67_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_250 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6825_ net69 _0284_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BitStream_buffer_output\[2\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__2884_ _2884_ vssd1 vssd1 vccd1 vccd1 clknet_0__2884_ sky130_fd_sc_hd__clkbuf_16
XFILLER_23_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6756_ net160 _0215_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[64\]
+ sky130_fd_sc_hd__dfxtp_1
X_3968_ _0428_ _0446_ _0466_ _0481_ vssd1 vssd1 vccd1 vccd1 _0482_ sky130_fd_sc_hd__and4_1
XFILLER_50_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5707_ _0453_ _3217_ vssd1 vssd1 vccd1 vccd1 _2208_ sky130_fd_sc_hd__nand2_1
XFILLER_12_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3899_ _3052_ _2933_ vssd1 vssd1 vccd1 vccd1 _0413_ sky130_fd_sc_hd__and2_1
X_5638_ _3100_ _3324_ _3326_ _0714_ _2139_ vssd1 vssd1 vccd1 vccd1 _2140_ sky130_fd_sc_hd__a221oi_1
X_5569_ _1947_ _2071_ vssd1 vssd1 vccd1 vccd1 _0286_ sky130_fd_sc_hd__nor2_1
XFILLER_77_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4940_ _3162_ egd_top.BitStream_buffer.BS_buffer\[119\] vssd1 vssd1 vccd1 vccd1 _1448_
+ sky130_fd_sc_hd__nand2_1
XFILLER_64_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4871_ _1368_ _1372_ _1374_ _1378_ vssd1 vssd1 vccd1 vccd1 _1379_ sky130_fd_sc_hd__and4_1
X_3822_ _3209_ _0335_ vssd1 vssd1 vccd1 vccd1 _0336_ sky130_fd_sc_hd__nor2_1
XFILLER_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3753_ _3229_ _3247_ _3267_ _3286_ vssd1 vssd1 vccd1 vccd1 _3287_ sky130_fd_sc_hd__and4_1
X_3684_ _3104_ _3213_ vssd1 vssd1 vccd1 vccd1 _3218_ sky130_fd_sc_hd__nand2_1
X_6472_ _2827_ _2685_ vssd1 vssd1 vccd1 vccd1 _2835_ sky130_fd_sc_hd__nand2_1
X_5423_ _1916_ _1919_ _1923_ _1926_ vssd1 vssd1 vccd1 vccd1 _1927_ sky130_fd_sc_hd__and4_1
X_5354_ egd_top.BitStream_buffer.BS_buffer\[32\] _0514_ _0901_ _0365_ vssd1 vssd1
+ vccd1 vccd1 _1858_ sky130_fd_sc_hd__a22o_1
X_4305_ _3168_ _3153_ vssd1 vssd1 vccd1 vccd1 _0817_ sky130_fd_sc_hd__nand2_1
X_5285_ _0400_ _0341_ _0344_ egd_top.BitStream_buffer.BS_buffer\[46\] vssd1 vssd1
+ vccd1 vccd1 _1790_ sky130_fd_sc_hd__a22o_1
X_4236_ _0736_ _0740_ _0743_ _0748_ vssd1 vssd1 vccd1 vccd1 _0749_ sky130_fd_sc_hd__and4_1
X_4167_ _0679_ _0587_ vssd1 vssd1 vccd1 vccd1 _0680_ sky130_fd_sc_hd__or2_1
XFILLER_28_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4098_ _3071_ _0556_ vssd1 vssd1 vccd1 vccd1 _0612_ sky130_fd_sc_hd__nand2_1
XFILLER_82_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6808_ net52 _0267_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[12\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_11_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6739_ net143 _0198_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[97\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_2_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5070_ _3252_ _3216_ _3268_ _3220_ _1576_ vssd1 vssd1 vccd1 vccd1 _1577_ sky130_fd_sc_hd__a221oi_1
X_4021_ _0528_ _0530_ _0532_ _0534_ vssd1 vssd1 vccd1 vccd1 _0535_ sky130_fd_sc_hd__o22a_1
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5972_ _2449_ _0574_ vssd1 vssd1 vccd1 vccd1 _2457_ sky130_fd_sc_hd__nand2_1
XFILLER_64_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4923_ _3242_ egd_top.BitStream_buffer.BS_buffer\[70\] vssd1 vssd1 vccd1 vccd1 _1431_
+ sky130_fd_sc_hd__nand2_1
X_4854_ _1360_ _2935_ _1361_ vssd1 vssd1 vccd1 vccd1 _1362_ sky130_fd_sc_hd__o21ai_1
X_3805_ _3290_ _3077_ vssd1 vssd1 vccd1 vccd1 _3339_ sky130_fd_sc_hd__nor2_2
XFILLER_20_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4785_ _0447_ _0431_ _0435_ _0467_ vssd1 vssd1 vccd1 vccd1 _1294_ sky130_fd_sc_hd__a22o_1
X_3736_ _3269_ vssd1 vssd1 vccd1 vccd1 _3270_ sky130_fd_sc_hd__clkinv_2
X_6524_ clknet_1_1__leaf__2882_ vssd1 vssd1 vccd1 vccd1 _2883_ sky130_fd_sc_hd__buf_1
X_3667_ _3090_ _3134_ vssd1 vssd1 vccd1 vccd1 _3201_ sky130_fd_sc_hd__and2_1
X_6455_ _2817_ _2818_ vssd1 vssd1 vccd1 vccd1 _2819_ sky130_fd_sc_hd__nor2_1
X_3598_ _3065_ _3084_ _3108_ _3131_ vssd1 vssd1 vccd1 vccd1 _3132_ sky130_fd_sc_hd__and4_1
X_6386_ _2752_ _2755_ vssd1 vssd1 vccd1 vccd1 _2756_ sky130_fd_sc_hd__nand2_1
X_5406_ _3328_ _3279_ _1909_ vssd1 vssd1 vccd1 vccd1 _1910_ sky130_fd_sc_hd__o21ai_1
XFILLER_87_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5337_ _0454_ _0406_ _1839_ _1840_ vssd1 vssd1 vccd1 vccd1 _1841_ sky130_fd_sc_hd__a211oi_1
X_5268_ _0442_ _0471_ vssd1 vssd1 vccd1 vccd1 _1773_ sky130_fd_sc_hd__nand2_1
X_4219_ _3169_ _3081_ _3082_ _0726_ _0731_ vssd1 vssd1 vccd1 vccd1 _0732_ sky130_fd_sc_hd__a221oi_1
XFILLER_75_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5199_ egd_top.BitStream_buffer.BitStream_buffer_output\[7\] vssd1 vssd1 vccd1 vccd1
+ _1705_ sky130_fd_sc_hd__inv_2
XFILLER_18_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_507 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4570_ egd_top.BitStream_buffer.BitStream_buffer_output\[11\] _2965_ _0627_ vssd1
+ vssd1 vccd1 vccd1 _1080_ sky130_fd_sc_hd__o21ai_1
X_3521_ _3054_ vssd1 vssd1 vccd1 vccd1 _3055_ sky130_fd_sc_hd__inv_2
X_6240_ _3008_ _2603_ _2611_ _2616_ vssd1 vssd1 vccd1 vccd1 _0166_ sky130_fd_sc_hd__o211a_1
X_3452_ egd_top.BitStream_buffer.BS_buffer\[118\] vssd1 vssd1 vccd1 vccd1 _2996_ sky130_fd_sc_hd__inv_2
X_3383_ egd_top.BitStream_buffer.pc\[6\] _2936_ vssd1 vssd1 vccd1 vccd1 _2937_ sky130_fd_sc_hd__nor2_1
X_6171_ _2553_ _0808_ vssd1 vssd1 vccd1 vccd1 _2573_ sky130_fd_sc_hd__nand2_1
X_5122_ _3315_ _3271_ _0774_ _3275_ _1627_ vssd1 vssd1 vccd1 vccd1 _1628_ sky130_fd_sc_hd__a221oi_1
XFILLER_69_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5053_ _0323_ _3100_ vssd1 vssd1 vccd1 vccd1 _1560_ sky130_fd_sc_hd__nand2_1
X_4004_ _0502_ _0504_ _0505_ _0508_ _0517_ vssd1 vssd1 vccd1 vccd1 _0518_ sky130_fd_sc_hd__a221oi_1
XFILLER_37_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5955_ _2443_ _0597_ vssd1 vssd1 vccd1 vccd1 _2448_ sky130_fd_sc_hd__nand2_1
X_4906_ _3092_ _3109_ vssd1 vssd1 vccd1 vccd1 _1414_ sky130_fd_sc_hd__nand2_1
XFILLER_52_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5886_ _0955_ _0425_ vssd1 vssd1 vccd1 vccd1 _2386_ sky130_fd_sc_hd__or2_1
XFILLER_21_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4837_ _0405_ _0443_ vssd1 vssd1 vccd1 vccd1 _1345_ sky130_fd_sc_hd__nand2_1
X_4768_ _0371_ _0346_ vssd1 vssd1 vccd1 vccd1 _1277_ sky130_fd_sc_hd__nand2_1
X_3719_ _3114_ _3212_ vssd1 vssd1 vccd1 vccd1 _3253_ sky130_fd_sc_hd__and2_1
X_4699_ _3333_ _0785_ vssd1 vssd1 vccd1 vccd1 _1208_ sky130_fd_sc_hd__nand2_1
X_6507_ _2860_ vssd1 vssd1 vccd1 vccd1 _2869_ sky130_fd_sc_hd__inv_2
X_6438_ _2742_ _2801_ vssd1 vssd1 vccd1 vccd1 _2802_ sky130_fd_sc_hd__nor2_1
XFILLER_88_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6369_ _2739_ _2701_ vssd1 vssd1 vccd1 vccd1 _2740_ sky130_fd_sc_hd__nor2_1
XFILLER_48_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_88 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_8 _1581_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5740_ _0633_ _0506_ _2238_ _2239_ _2240_ vssd1 vssd1 vccd1 vccd1 _2241_ sky130_fd_sc_hd__o2111a_1
X_5671_ _3066_ _3039_ _3070_ _3048_ _2172_ vssd1 vssd1 vccd1 vccd1 _2173_ sky130_fd_sc_hd__a221oi_1
X_4622_ _0513_ _0531_ vssd1 vssd1 vccd1 vccd1 _1132_ sky130_fd_sc_hd__nand2_1
X_4553_ _3155_ egd_top.BitStream_buffer.BS_buffer\[117\] vssd1 vssd1 vccd1 vccd1 _1064_
+ sky130_fd_sc_hd__nand2_1
X_4484_ egd_top.BitStream_buffer.BS_buffer\[32\] vssd1 vssd1 vccd1 vccd1 _0995_ sky130_fd_sc_hd__inv_2
X_3504_ _3037_ vssd1 vssd1 vccd1 vccd1 _3038_ sky130_fd_sc_hd__clkbuf_2
X_3435_ egd_top.BitStream_buffer.BS_buffer\[114\] vssd1 vssd1 vccd1 vccd1 _2983_ sky130_fd_sc_hd__clkinv_2
X_6223_ _2603_ _1007_ vssd1 vssd1 vccd1 vccd1 _2607_ sky130_fd_sc_hd__nand2_1
XFILLER_85_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3366_ egd_top.BitStream_buffer.pc\[2\] egd_top.BitStream_buffer.pc\[3\] vssd1 vssd1
+ vccd1 vccd1 _2920_ sky130_fd_sc_hd__nand2_4
X_6154_ _2561_ _0713_ vssd1 vssd1 vccd1 vccd1 _2564_ sky130_fd_sc_hd__nand2_1
X_5105_ _3018_ _3200_ _1610_ vssd1 vssd1 vccd1 vccd1 _1611_ sky130_fd_sc_hd__o21ai_1
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6085_ _3005_ _2510_ _2516_ _2523_ vssd1 vssd1 vccd1 vccd1 _0222_ sky130_fd_sc_hd__o211a_1
X_5036_ _3149_ _3156_ _3133_ _3160_ _1542_ vssd1 vssd1 vccd1 vccd1 _1543_ sky130_fd_sc_hd__a221oi_1
XFILLER_85_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5938_ _2972_ _2901_ _2435_ vssd1 vssd1 vccd1 vccd1 _2436_ sky130_fd_sc_hd__and3_1
XFILLER_15_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5869_ _0676_ _3183_ _2368_ vssd1 vssd1 vccd1 vccd1 _2369_ sky130_fd_sc_hd__o21ai_1
XFILLER_5_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_89 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput23 net23 vssd1 vssd1 vccd1 vccd1 la_data_out_23_16[3] sky130_fd_sc_hd__buf_12
Xoutput34 net34 vssd1 vssd1 vccd1 vccd1 la_data_out_30_27[3] sky130_fd_sc_hd__buf_12
XFILLER_0_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6556__100 clknet_1_0__leaf__2886_ vssd1 vssd1 vccd1 vccd1 net134 sky130_fd_sc_hd__inv_2
XFILLER_12_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6841_ net85 _0300_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[125\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_35_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3984_ egd_top.BitStream_buffer.BS_buffer\[19\] vssd1 vssd1 vccd1 vccd1 _0498_ sky130_fd_sc_hd__clkbuf_4
XFILLER_22_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6772_ net176 _0231_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[48\]
+ sky130_fd_sc_hd__dfxtp_1
X_5723_ _0581_ _0509_ vssd1 vssd1 vccd1 vccd1 _2224_ sky130_fd_sc_hd__nand2_1
X_5654_ _2147_ _2150_ _2153_ _2155_ vssd1 vssd1 vccd1 vccd1 _2156_ sky130_fd_sc_hd__and4_1
XFILLER_30_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4605_ _0586_ _0570_ vssd1 vssd1 vccd1 vccd1 _1115_ sky130_fd_sc_hd__or2_1
X_5585_ _0887_ _0421_ _2086_ vssd1 vssd1 vccd1 vccd1 _2087_ sky130_fd_sc_hd__o21ai_1
X_4536_ _1043_ _3239_ _1044_ _1045_ _1046_ vssd1 vssd1 vccd1 vccd1 _1047_ sky130_fd_sc_hd__o2111a_1
X_4467_ _0688_ _0575_ _0975_ _0976_ _0977_ vssd1 vssd1 vccd1 vccd1 _0978_ sky130_fd_sc_hd__o2111a_1
X_4398_ egd_top.BitStream_buffer.BS_buffer\[32\] _0539_ _0365_ _0542_ _0909_ vssd1
+ vssd1 vccd1 vccd1 _0910_ sky130_fd_sc_hd__a221oi_1
XFILLER_77_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6206_ _2902_ egd_top.BitStream_buffer.pc\[2\] vssd1 vssd1 vccd1 vccd1 _2597_ sky130_fd_sc_hd__nand2_1
X_3418_ _2910_ _2903_ vssd1 vssd1 vccd1 vccd1 _2968_ sky130_fd_sc_hd__and2_1
X_6137_ _2552_ vssd1 vssd1 vccd1 vccd1 _2553_ sky130_fd_sc_hd__clkinv_2
X_3349_ net31 vssd1 vssd1 vccd1 vccd1 _2906_ sky130_fd_sc_hd__inv_2
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6068_ _2511_ _0659_ vssd1 vssd1 vccd1 vccd1 _2514_ sky130_fd_sc_hd__nand2_1
XFILLER_85_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5019_ _3093_ _3118_ vssd1 vssd1 vccd1 vccd1 _1526_ sky130_fd_sc_hd__nand2_1
XFILLER_26_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5370_ _0582_ _0502_ vssd1 vssd1 vccd1 vccd1 _1874_ sky130_fd_sc_hd__nand2_1
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4321_ egd_top.BitStream_buffer.BS_buffer\[74\] vssd1 vssd1 vccd1 vccd1 _0833_ sky130_fd_sc_hd__clkinv_2
X_6695__66 clknet_1_1__leaf__2899_ vssd1 vssd1 vccd1 vccd1 net100 sky130_fd_sc_hd__inv_2
X_4252_ _3272_ _3271_ _3283_ _3275_ _0764_ vssd1 vssd1 vccd1 vccd1 _0765_ sky130_fd_sc_hd__a221oi_1
XFILLER_86_107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4183_ _0514_ _0509_ vssd1 vssd1 vccd1 vccd1 _0696_ sky130_fd_sc_hd__nand2_1
XFILLER_67_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6824_ net68 _0283_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BitStream_buffer_output\[1\]
+ sky130_fd_sc_hd__dfxtp_2
Xclkbuf_0__2883_ _2883_ vssd1 vssd1 vccd1 vccd1 clknet_0__2883_ sky130_fd_sc_hd__clkbuf_16
X_6755_ net159 _0214_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[65\]
+ sky130_fd_sc_hd__dfxtp_1
X_3967_ _0467_ _0470_ _0471_ _0473_ _0480_ vssd1 vssd1 vccd1 vccd1 _0481_ sky130_fd_sc_hd__a221oi_1
X_5706_ _0457_ egd_top.BitStream_buffer.BS_buffer\[71\] vssd1 vssd1 vccd1 vccd1 _2207_
+ sky130_fd_sc_hd__nand2_1
X_3898_ egd_top.BitStream_buffer.BS_buffer\[50\] vssd1 vssd1 vccd1 vccd1 _0412_ sky130_fd_sc_hd__clkbuf_4
X_5637_ _3102_ _3330_ _2138_ vssd1 vssd1 vccd1 vccd1 _2139_ sky130_fd_sc_hd__o21ai_1
XFILLER_12_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5568_ _3026_ _2070_ vssd1 vssd1 vccd1 vccd1 _2071_ sky130_fd_sc_hd__nor2_1
XFILLER_88_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4519_ _3060_ egd_top.BitStream_buffer.BS_buffer\[102\] vssd1 vssd1 vccd1 vccd1 _1030_
+ sky130_fd_sc_hd__nand2_1
XFILLER_2_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5499_ _3147_ _0566_ vssd1 vssd1 vccd1 vccd1 _2002_ sky130_fd_sc_hd__nand2_1
XFILLER_58_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4870_ _0986_ _0603_ _1375_ _1376_ _1377_ vssd1 vssd1 vccd1 vccd1 _1378_ sky130_fd_sc_hd__o2111a_1
X_3821_ _3287_ _0334_ vssd1 vssd1 vccd1 vccd1 _0335_ sky130_fd_sc_hd__nand2_1
XFILLER_20_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3752_ _3268_ _3271_ _3272_ _3275_ _3285_ vssd1 vssd1 vccd1 vccd1 _3286_ sky130_fd_sc_hd__a221oi_1
XFILLER_9_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6471_ _2831_ _2834_ vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__nand2_1
X_3683_ egd_top.BitStream_buffer.BS_buffer\[69\] vssd1 vssd1 vccd1 vccd1 _3217_ sky130_fd_sc_hd__clkbuf_4
X_5422_ _0744_ _0726_ _3149_ _3081_ _1925_ vssd1 vssd1 vccd1 vccd1 _1926_ sky130_fd_sc_hd__a221oi_1
X_5353_ _1842_ _1856_ vssd1 vssd1 vccd1 vccd1 _1857_ sky130_fd_sc_hd__nand2_1
X_4304_ _3163_ _3157_ vssd1 vssd1 vccd1 vccd1 _0816_ sky130_fd_sc_hd__nand2_1
XFILLER_87_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5284_ _0948_ _0378_ _0412_ _0382_ _1788_ vssd1 vssd1 vccd1 vccd1 _1789_ sky130_fd_sc_hd__a221oi_1
XFILLER_87_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4235_ _0745_ _0747_ vssd1 vssd1 vccd1 vccd1 _0748_ sky130_fd_sc_hd__nor2_1
X_4166_ _0583_ vssd1 vssd1 vccd1 vccd1 _0679_ sky130_fd_sc_hd__inv_2
XFILLER_67_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4097_ egd_top.BitStream_buffer.BS_buffer\[13\] vssd1 vssd1 vccd1 vccd1 _0611_ sky130_fd_sc_hd__inv_2
XFILLER_82_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6807_ net51 _0266_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[13\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_23_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4999_ _0561_ egd_top.BitStream_buffer.BS_buffer\[13\] vssd1 vssd1 vccd1 vccd1 _1506_
+ sky130_fd_sc_hd__nand2_1
XFILLER_23_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6738_ net142 _0197_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[98\]
+ sky130_fd_sc_hd__dfxtp_1
X_6617__155 clknet_1_0__leaf__2892_ vssd1 vssd1 vccd1 vccd1 net189 sky130_fd_sc_hd__inv_2
XFILLER_2_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6659__33 clknet_1_0__leaf__2896_ vssd1 vssd1 vccd1 vccd1 net67 sky130_fd_sc_hd__inv_2
XFILLER_2_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6674__47 clknet_1_0__leaf__2897_ vssd1 vssd1 vccd1 vccd1 net81 sky130_fd_sc_hd__inv_2
XFILLER_19_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_493 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4020_ _0533_ vssd1 vssd1 vccd1 vccd1 _0534_ sky130_fd_sc_hd__buf_2
XFILLER_84_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5971_ _3008_ _2443_ _2446_ _2456_ vssd1 vssd1 vccd1 vccd1 _0269_ sky130_fd_sc_hd__o211a_1
X_4922_ egd_top.BitStream_buffer.BS_buffer\[71\] vssd1 vssd1 vccd1 vccd1 _1430_ sky130_fd_sc_hd__inv_2
XFILLER_45_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4853_ _0476_ egd_top.BitStream_buffer.BS_buffer\[68\] vssd1 vssd1 vccd1 vccd1 _1361_
+ sky130_fd_sc_hd__nand2_1
X_4784_ _0663_ _0450_ _1290_ _1291_ _1292_ vssd1 vssd1 vccd1 vccd1 _1293_ sky130_fd_sc_hd__o2111a_1
XFILLER_20_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3804_ egd_top.BitStream_buffer.BS_buffer\[94\] vssd1 vssd1 vccd1 vccd1 _3338_ sky130_fd_sc_hd__clkbuf_4
X_3735_ _3067_ _3213_ vssd1 vssd1 vccd1 vccd1 _3269_ sky130_fd_sc_hd__nand2_1
X_6523_ wb_clk_i vssd1 vssd1 vccd1 vccd1 _2882_ sky130_fd_sc_hd__buf_1
X_6454_ _2739_ _2788_ _2764_ vssd1 vssd1 vccd1 vccd1 _2818_ sky130_fd_sc_hd__nand3_1
X_3666_ _3199_ vssd1 vssd1 vccd1 vccd1 _3200_ sky130_fd_sc_hd__buf_2
X_5405_ _3282_ _3334_ vssd1 vssd1 vccd1 vccd1 _1909_ sky130_fd_sc_hd__nand2_1
X_3597_ _3109_ _3113_ _3117_ _3118_ _3130_ vssd1 vssd1 vccd1 vccd1 _3131_ sky130_fd_sc_hd__a221oi_1
X_6385_ _2753_ _2754_ _2670_ vssd1 vssd1 vccd1 vccd1 _2755_ sky130_fd_sc_hd__o21ai_1
X_5336_ _0429_ _0395_ _0398_ _0436_ vssd1 vssd1 vccd1 vccd1 _1840_ sky130_fd_sc_hd__a22o_1
X_5267_ _0447_ _0415_ _0467_ _0419_ _1771_ vssd1 vssd1 vccd1 vccd1 _1772_ sky130_fd_sc_hd__a221oi_1
XFILLER_87_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4218_ _0727_ _0729_ _0730_ vssd1 vssd1 vccd1 vccd1 _0731_ sky130_fd_sc_hd__o21ai_1
X_5198_ _1645_ _1702_ _1703_ vssd1 vssd1 vccd1 vccd1 _1704_ sky130_fd_sc_hd__nand3_1
X_4149_ _0660_ _0661_ vssd1 vssd1 vccd1 vccd1 _0662_ sky130_fd_sc_hd__nor2_1
XFILLER_70_102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_30 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3520_ _3035_ _3053_ vssd1 vssd1 vccd1 vccd1 _3054_ sky130_fd_sc_hd__nor2_1
XFILLER_6_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3451_ net16 vssd1 vssd1 vccd1 vccd1 _2995_ sky130_fd_sc_hd__clkbuf_4
X_3382_ _2935_ vssd1 vssd1 vccd1 vccd1 _2936_ sky130_fd_sc_hd__inv_2
X_6638__14 clknet_1_1__leaf__2894_ vssd1 vssd1 vccd1 vccd1 net48 sky130_fd_sc_hd__inv_2
X_6170_ _3017_ _2555_ _2570_ _2572_ vssd1 vssd1 vccd1 vccd1 _0186_ sky130_fd_sc_hd__o211a_1
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5121_ _3306_ _3279_ _1626_ vssd1 vssd1 vccd1 vccd1 _1627_ sky130_fd_sc_hd__o21ai_1
XFILLER_84_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6653__28 clknet_1_1__leaf__2895_ vssd1 vssd1 vccd1 vccd1 net62 sky130_fd_sc_hd__inv_2
X_5052_ _1554_ _1558_ vssd1 vssd1 vccd1 vccd1 _1559_ sky130_fd_sc_hd__nand2_1
X_4003_ _0510_ _0512_ _0516_ vssd1 vssd1 vccd1 vccd1 _0517_ sky130_fd_sc_hd__o21ai_1
XFILLER_84_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__2889_ clknet_0__2889_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__2889_
+ sky130_fd_sc_hd__clkbuf_16
X_5954_ _2982_ _2442_ _2446_ _2447_ vssd1 vssd1 vccd1 vccd1 _0277_ sky130_fd_sc_hd__o211a_1
X_4905_ _0718_ _3055_ _1410_ _1411_ _1412_ vssd1 vssd1 vccd1 vccd1 _1413_ sky130_fd_sc_hd__o2111a_1
XFILLER_40_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5885_ _2375_ _2378_ _2381_ _2384_ vssd1 vssd1 vccd1 vccd1 _2385_ sky130_fd_sc_hd__and4_1
X_4836_ _0874_ _0388_ _0948_ _0944_ _1343_ vssd1 vssd1 vccd1 vccd1 _1344_ sky130_fd_sc_hd__a221oi_1
XFILLER_33_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4767_ _0354_ vssd1 vssd1 vccd1 vccd1 _1276_ sky130_fd_sc_hd__inv_2
X_6506_ _2867_ _2860_ vssd1 vssd1 vccd1 vccd1 _2868_ sky130_fd_sc_hd__nand2_1
X_4698_ egd_top.BitStream_buffer.BitStream_buffer_output\[10\] _2965_ _0627_ vssd1
+ vssd1 vccd1 vccd1 _1207_ sky130_fd_sc_hd__o21ai_1
X_3718_ egd_top.BitStream_buffer.BS_buffer\[75\] vssd1 vssd1 vccd1 vccd1 _3252_ sky130_fd_sc_hd__clkbuf_4
X_3649_ _3182_ vssd1 vssd1 vccd1 vccd1 _3183_ sky130_fd_sc_hd__clkbuf_4
X_6437_ _2777_ _2745_ vssd1 vssd1 vccd1 vccd1 _2801_ sky130_fd_sc_hd__nand2_1
X_6368_ _2738_ vssd1 vssd1 vccd1 vccd1 _2739_ sky130_fd_sc_hd__inv_2
XFILLER_88_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5319_ _1813_ _1817_ _1819_ _1823_ vssd1 vssd1 vccd1 vccd1 _1824_ sky130_fd_sc_hd__and4_1
XFILLER_0_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6299_ _2669_ vssd1 vssd1 vccd1 vccd1 _2670_ sky130_fd_sc_hd__inv_2
XFILLER_29_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_9 _1977_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_282 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5670_ _0808_ _3056_ _2171_ vssd1 vssd1 vccd1 vccd1 _2172_ sky130_fd_sc_hd__o21ai_1
XFILLER_15_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4621_ _0502_ _0486_ _0505_ _0489_ _1130_ vssd1 vssd1 vccd1 vccd1 _1131_ sky130_fd_sc_hd__a221oi_1
X_4552_ _3167_ egd_top.BitStream_buffer.BS_buffer\[115\] vssd1 vssd1 vccd1 vccd1 _1063_
+ sky130_fd_sc_hd__nand2_1
X_4483_ _0532_ _0512_ _0991_ _0992_ _0993_ vssd1 vssd1 vccd1 vccd1 _0994_ sky130_fd_sc_hd__o2111a_1
X_3503_ _3033_ _3036_ vssd1 vssd1 vccd1 vccd1 _3037_ sky130_fd_sc_hd__and2_1
X_6222_ _2982_ _2602_ _2570_ _2606_ vssd1 vssd1 vccd1 vccd1 _0174_ sky130_fd_sc_hd__o211a_1
X_3434_ net5 vssd1 vssd1 vccd1 vccd1 _2982_ sky130_fd_sc_hd__buf_4
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3365_ net30 net29 vssd1 vssd1 vccd1 vccd1 _2919_ sky130_fd_sc_hd__nand2_1
X_6153_ _2992_ _2554_ _2558_ _2563_ vssd1 vssd1 vccd1 vccd1 _0194_ sky130_fd_sc_hd__o211a_1
X_5104_ _3203_ _3173_ vssd1 vssd1 vccd1 vccd1 _1610_ sky130_fd_sc_hd__nand2_1
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6084_ _2517_ _0462_ vssd1 vssd1 vccd1 vccd1 _2523_ sky130_fd_sc_hd__nand2_1
X_5035_ _1540_ _1541_ vssd1 vssd1 vccd1 vccd1 _1542_ sky130_fd_sc_hd__nand2_1
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5937_ _2971_ _2938_ vssd1 vssd1 vccd1 vccd1 _2435_ sky130_fd_sc_hd__nand2_1
XFILLER_13_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5868_ _3185_ egd_top.BitStream_buffer.BS_buffer\[13\] vssd1 vssd1 vccd1 vccd1 _2368_
+ sky130_fd_sc_hd__nand2_1
X_4819_ _0492_ _0613_ _1325_ _1326_ _1327_ vssd1 vssd1 vccd1 vccd1 _1328_ sky130_fd_sc_hd__o2111a_1
X_5799_ _0329_ _0722_ vssd1 vssd1 vccd1 vccd1 _2300_ sky130_fd_sc_hd__nand2_1
XFILLER_31_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput24 net24 vssd1 vssd1 vccd1 vccd1 la_data_out_23_16[4] sky130_fd_sc_hd__buf_12
XFILLER_0_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_474 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6840_ net84 _0299_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[126\]
+ sky130_fd_sc_hd__dfxtp_2
X_6771_ net175 _0230_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[49\]
+ sky130_fd_sc_hd__dfxtp_1
X_3983_ _0496_ vssd1 vssd1 vccd1 vccd1 _0497_ sky130_fd_sc_hd__buf_4
X_5722_ _0577_ _0505_ vssd1 vssd1 vccd1 vccd1 _2223_ sky130_fd_sc_hd__nand2_1
XFILLER_62_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5653_ _3334_ _3271_ _0780_ _3275_ _2154_ vssd1 vssd1 vccd1 vccd1 _2155_ sky130_fd_sc_hd__a221oi_1
X_4604_ _0560_ _0583_ vssd1 vssd1 vccd1 vccd1 _1114_ sky130_fd_sc_hd__nand2_1
X_5584_ _0647_ _0424_ vssd1 vssd1 vccd1 vccd1 _2086_ sky130_fd_sc_hd__or2_1
X_4535_ _3235_ _3221_ vssd1 vssd1 vccd1 vccd1 _1046_ sky130_fd_sc_hd__nand2_1
X_4466_ _0676_ _0587_ vssd1 vssd1 vccd1 vccd1 _0977_ sky130_fd_sc_hd__or2_1
X_4397_ _0907_ _0546_ _0908_ vssd1 vssd1 vccd1 vccd1 _0909_ sky130_fd_sc_hd__o21ai_1
X_3417_ egd_top.BitStream_buffer.buffer_index\[6\] vssd1 vssd1 vccd1 vccd1 _2967_
+ sky130_fd_sc_hd__inv_2
X_6205_ _2596_ _2579_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.pc\[2\] sky130_fd_sc_hd__xnor2_4
XFILLER_58_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6136_ _2970_ net198 net196 _2939_ vssd1 vssd1 vccd1 vccd1 _2552_ sky130_fd_sc_hd__and4_1
X_3348_ _2904_ vssd1 vssd1 vccd1 vccd1 _2905_ sky130_fd_sc_hd__clkinv_2
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6067_ _2979_ _2510_ _2501_ _2513_ vssd1 vssd1 vccd1 vccd1 _0230_ sky130_fd_sc_hd__o211a_1
XFILLER_45_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5018_ _0714_ _3039_ _3128_ _3048_ _1524_ vssd1 vssd1 vccd1 vccd1 _1525_ sky130_fd_sc_hd__a221oi_2
XFILLER_53_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6586__127 clknet_1_1__leaf__2889_ vssd1 vssd1 vccd1 vccd1 net161 sky130_fd_sc_hd__inv_2
XFILLER_76_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4320_ _3210_ _3233_ _3236_ _3217_ _0831_ vssd1 vssd1 vccd1 vccd1 _0832_ sky130_fd_sc_hd__a221oi_1
X_4251_ _3296_ _3279_ _0763_ vssd1 vssd1 vccd1 vccd1 _0764_ sky130_fd_sc_hd__o21ai_1
XFILLER_4_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4182_ egd_top.BitStream_buffer.BS_buffer\[17\] _0487_ _0491_ _0490_ _0694_ vssd1
+ vssd1 vccd1 vccd1 _0695_ sky130_fd_sc_hd__a221oi_1
XFILLER_35_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6823_ net67 _0282_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.buffer_index\[6\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__2882_ _2882_ vssd1 vssd1 vccd1 vccd1 clknet_0__2882_ sky130_fd_sc_hd__clkbuf_16
XFILLER_50_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6754_ net158 _0213_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[66\]
+ sky130_fd_sc_hd__dfxtp_1
X_3966_ _0474_ _2935_ _0479_ vssd1 vssd1 vccd1 vccd1 _0480_ sky130_fd_sc_hd__o21ai_1
XFILLER_50_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5705_ _0664_ _0414_ _3244_ _0418_ _2205_ vssd1 vssd1 vccd1 vccd1 _2206_ sky130_fd_sc_hd__a221oi_1
X_3897_ _0357_ _0374_ _0392_ _0410_ vssd1 vssd1 vccd1 vccd1 _0411_ sky130_fd_sc_hd__and4_1
X_5636_ _3333_ _3094_ vssd1 vssd1 vccd1 vccd1 _2138_ sky130_fd_sc_hd__nand2_1
X_5567_ _2011_ _2068_ _2069_ vssd1 vssd1 vccd1 vccd1 _2070_ sky130_fd_sc_hd__nand3_1
X_5498_ _1997_ _1998_ _1999_ _2000_ vssd1 vssd1 vccd1 vccd1 _2001_ sky130_fd_sc_hd__and4_1
X_4518_ _1025_ _3122_ _1026_ _1027_ _1028_ vssd1 vssd1 vccd1 vccd1 _1029_ sky130_fd_sc_hd__o2111a_1
X_4449_ _0443_ vssd1 vssd1 vccd1 vccd1 _0960_ sky130_fd_sc_hd__inv_2
X_6540__85 clknet_1_1__leaf__2885_ vssd1 vssd1 vccd1 vccd1 net119 sky130_fd_sc_hd__inv_2
XFILLER_85_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6119_ _2904_ vssd1 vssd1 vccd1 vccd1 _2543_ sky130_fd_sc_hd__clkbuf_4
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3820_ _3305_ _3321_ _3337_ _0333_ vssd1 vssd1 vccd1 vccd1 _0334_ sky130_fd_sc_hd__and4_1
XFILLER_32_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3751_ _3277_ _3279_ _3284_ vssd1 vssd1 vccd1 vccd1 _3285_ sky130_fd_sc_hd__o21ai_1
XFILLER_71_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3682_ _3215_ vssd1 vssd1 vccd1 vccd1 _3216_ sky130_fd_sc_hd__clkbuf_4
X_6470_ _2833_ _2788_ vssd1 vssd1 vccd1 vccd1 _2834_ sky130_fd_sc_hd__nand2_1
X_5421_ _2996_ _0729_ _1924_ vssd1 vssd1 vccd1 vccd1 _1925_ sky130_fd_sc_hd__o21ai_1
X_5352_ _1845_ _1848_ _1852_ _1855_ vssd1 vssd1 vccd1 vccd1 _1856_ sky130_fd_sc_hd__and4_1
X_4303_ _3173_ _3137_ _3177_ _3141_ _0814_ vssd1 vssd1 vccd1 vccd1 _0815_ sky130_fd_sc_hd__a221oi_1
XFILLER_87_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5283_ _0960_ _0385_ _1787_ vssd1 vssd1 vccd1 vccd1 _1788_ sky130_fd_sc_hd__o21ai_1
X_4234_ _3104_ egd_top.BitStream_buffer.BS_buffer\[118\] _3142_ _0746_ _3202_ vssd1
+ vssd1 vccd1 vccd1 _0747_ sky130_fd_sc_hd__a32o_1
X_4165_ _0582_ egd_top.BitStream_buffer.BS_buffer\[11\] vssd1 vssd1 vccd1 vccd1 _0678_
+ sky130_fd_sc_hd__nand2_1
XFILLER_82_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4096_ _0609_ egd_top.BitStream_buffer.BS_buffer\[14\] vssd1 vssd1 vccd1 vccd1 _0610_
+ sky130_fd_sc_hd__nand2_1
XFILLER_55_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6806_ net50 _0265_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[14\]
+ sky130_fd_sc_hd__dfxtp_4
X_4998_ _1496_ _1498_ _1501_ _1504_ vssd1 vssd1 vccd1 vccd1 _1505_ sky130_fd_sc_hd__and4_1
XFILLER_11_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6737_ net141 _0196_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[99\]
+ sky130_fd_sc_hd__dfxtp_1
X_3949_ _3121_ _2933_ vssd1 vssd1 vccd1 vccd1 _0463_ sky130_fd_sc_hd__nand2_2
X_6668_ clknet_1_0__leaf__2882_ vssd1 vssd1 vccd1 vccd1 _2897_ sky130_fd_sc_hd__buf_1
X_5619_ _0513_ egd_top.BitStream_buffer.BS_buffer\[34\] vssd1 vssd1 vccd1 vccd1 _2121_
+ sky130_fd_sc_hd__nand2_1
XFILLER_58_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5970_ _2449_ _0679_ vssd1 vssd1 vccd1 vccd1 _2456_ sky130_fd_sc_hd__nand2_1
X_4921_ _3248_ _3215_ _3252_ _3219_ _1428_ vssd1 vssd1 vccd1 vccd1 _1429_ sky130_fd_sc_hd__a221oi_1
XFILLER_60_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4852_ egd_top.BitStream_buffer.BS_buffer\[69\] vssd1 vssd1 vccd1 vccd1 _1360_ sky130_fd_sc_hd__clkinv_2
XFILLER_20_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3803_ _3322_ _3324_ _3326_ _3327_ _3336_ vssd1 vssd1 vccd1 vccd1 _3337_ sky130_fd_sc_hd__a221oi_1
X_4783_ _0955_ _0464_ vssd1 vssd1 vccd1 vccd1 _1292_ sky130_fd_sc_hd__or2_1
X_6522_ _2875_ _2832_ _2685_ _2878_ vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__a2bb2o_1
XFILLER_20_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3734_ egd_top.BitStream_buffer.BS_buffer\[76\] vssd1 vssd1 vccd1 vccd1 _3268_ sky130_fd_sc_hd__clkbuf_4
X_3665_ _3104_ _3142_ vssd1 vssd1 vccd1 vccd1 _3199_ sky130_fd_sc_hd__nand2_2
XFILLER_9_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6453_ _2816_ _2701_ vssd1 vssd1 vccd1 vccd1 _2817_ sky130_fd_sc_hd__nand2_1
X_5404_ _3283_ _3216_ _3276_ _3220_ _1907_ vssd1 vssd1 vccd1 vccd1 _1908_ sky130_fd_sc_hd__a221oi_1
X_3596_ _3119_ _3123_ _3129_ vssd1 vssd1 vccd1 vccd1 _3130_ sky130_fd_sc_hd__o21ai_1
X_6384_ _2635_ _2702_ vssd1 vssd1 vccd1 vccd1 _2754_ sky130_fd_sc_hd__nor2_1
X_5335_ _0462_ _0403_ vssd1 vssd1 vccd1 vccd1 _1839_ sky130_fd_sc_hd__nor2_1
XFILLER_87_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5266_ _0650_ _0422_ _1770_ vssd1 vssd1 vccd1 vccd1 _1771_ sky130_fd_sc_hd__o21ai_1
X_4217_ _3074_ _3075_ vssd1 vssd1 vccd1 vccd1 _0730_ sky130_fd_sc_hd__nand2_1
XFILLER_68_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5197_ _0622_ _0579_ vssd1 vssd1 vccd1 vccd1 _1703_ sky130_fd_sc_hd__nand2_1
X_4148_ _0416_ _0414_ _0418_ _0443_ vssd1 vssd1 vccd1 vccd1 _0661_ sky130_fd_sc_hd__a22o_1
XFILLER_83_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4079_ _0592_ vssd1 vssd1 vccd1 vccd1 _0593_ sky130_fd_sc_hd__buf_2
XFILLER_18_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3450_ _2992_ _2975_ _2913_ _2994_ vssd1 vssd1 vccd1 vccd1 _0308_ sky130_fd_sc_hd__o211a_1
X_3381_ _2931_ _2934_ vssd1 vssd1 vccd1 vccd1 _2935_ sky130_fd_sc_hd__nand2_4
XFILLER_69_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5120_ _3282_ _3311_ vssd1 vssd1 vccd1 vccd1 _1626_ sky130_fd_sc_hd__nand2_1
XFILLER_69_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5051_ _0784_ _3308_ _1555_ _1556_ _1557_ vssd1 vssd1 vccd1 vccd1 _1558_ sky130_fd_sc_hd__o2111a_1
X_4002_ _0514_ _0515_ vssd1 vssd1 vccd1 vccd1 _0516_ sky130_fd_sc_hd__nand2_1
XFILLER_84_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0__f__2888_ clknet_0__2888_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__2888_
+ sky130_fd_sc_hd__clkbuf_16
X_5953_ _2443_ _0591_ vssd1 vssd1 vccd1 vccd1 _2447_ sky130_fd_sc_hd__nand2_1
X_4904_ _3060_ _0722_ vssd1 vssd1 vccd1 vccd1 _1412_ sky130_fd_sc_hd__nand2_1
X_5884_ _0459_ _0396_ _0399_ _0447_ _2383_ vssd1 vssd1 vccd1 vccd1 _2384_ sky130_fd_sc_hd__a221oi_1
XFILLER_40_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4835_ _0401_ _0380_ _1342_ vssd1 vssd1 vccd1 vccd1 _1343_ sky130_fd_sc_hd__o21ai_1
X_4766_ _0379_ _0342_ _0345_ _0389_ _1274_ vssd1 vssd1 vccd1 vccd1 _1275_ sky130_fd_sc_hd__a221oi_1
X_3717_ _3250_ vssd1 vssd1 vccd1 vccd1 _3251_ sky130_fd_sc_hd__buf_6
X_6505_ _2819_ _2849_ vssd1 vssd1 vccd1 vccd1 _2867_ sky130_fd_sc_hd__nand2_1
X_4697_ _1080_ _1206_ vssd1 vssd1 vccd1 vccd1 _0293_ sky130_fd_sc_hd__nor2_1
X_3648_ _3181_ vssd1 vssd1 vccd1 vccd1 _3182_ sky130_fd_sc_hd__inv_2
X_6436_ _2800_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.exp_golomb_len\[3\]
+ sky130_fd_sc_hd__clkbuf_1
X_3579_ _3112_ vssd1 vssd1 vccd1 vccd1 _3113_ sky130_fd_sc_hd__buf_2
X_6367_ _2735_ _2684_ vssd1 vssd1 vccd1 vccd1 _2738_ sky130_fd_sc_hd__nand2_1
X_5318_ _0520_ _0604_ _1820_ _1821_ _1822_ vssd1 vssd1 vccd1 vccd1 _1823_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6298_ _2659_ _2668_ vssd1 vssd1 vccd1 vccd1 _2669_ sky130_fd_sc_hd__nand2_2
X_5249_ _0792_ _3144_ _3148_ _0930_ vssd1 vssd1 vccd1 vccd1 _1754_ sky130_fd_sc_hd__a22o_1
XFILLER_29_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4620_ _1128_ _0494_ _1129_ vssd1 vssd1 vccd1 vccd1 _1130_ sky130_fd_sc_hd__o21ai_1
X_4551_ _3159_ egd_top.BitStream_buffer.BS_buffer\[118\] vssd1 vssd1 vccd1 vccd1 _1062_
+ sky130_fd_sc_hd__nand2_1
X_4482_ _0507_ _0519_ vssd1 vssd1 vccd1 vccd1 _0993_ sky130_fd_sc_hd__nand2_1
X_3502_ _3035_ vssd1 vssd1 vccd1 vccd1 _3036_ sky130_fd_sc_hd__inv_2
X_6221_ _2603_ _0842_ vssd1 vssd1 vccd1 vccd1 _2606_ sky130_fd_sc_hd__nand2_1
X_3433_ _2979_ _2975_ _2913_ _2981_ vssd1 vssd1 vccd1 vccd1 _0312_ sky130_fd_sc_hd__o211a_1
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6152_ _2561_ _3102_ vssd1 vssd1 vccd1 vccd1 _2563_ sky130_fd_sc_hd__nand2_1
X_5103_ _3133_ _3156_ _3138_ _3160_ _1608_ vssd1 vssd1 vccd1 vccd1 _1609_ sky130_fd_sc_hd__a221oi_1
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3364_ _2917_ vssd1 vssd1 vccd1 vccd1 _2918_ sky130_fd_sc_hd__inv_2
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6083_ _3001_ _2510_ _2516_ _2522_ vssd1 vssd1 vccd1 vccd1 _0223_ sky130_fd_sc_hd__o211a_1
X_5034_ _3168_ _3198_ vssd1 vssd1 vccd1 vccd1 _1541_ sky130_fd_sc_hd__nand2_1
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5936_ _2434_ vssd1 vssd1 vccd1 vccd1 _0282_ sky130_fd_sc_hd__clkbuf_1
XFILLER_15_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5867_ _2363_ _2364_ _2365_ _2366_ vssd1 vssd1 vccd1 vccd1 _2367_ sky130_fd_sc_hd__and4_1
XFILLER_21_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4818_ _0897_ _0603_ vssd1 vssd1 vccd1 vccd1 _1327_ sky130_fd_sc_hd__or2_1
X_5798_ _0714_ _3324_ _3326_ _3128_ _2298_ vssd1 vssd1 vccd1 vccd1 _2299_ sky130_fd_sc_hd__a221oi_1
X_4749_ _3264_ _3215_ _3248_ _3220_ _1257_ vssd1 vssd1 vccd1 vccd1 _1258_ sky130_fd_sc_hd__a221oi_1
XFILLER_31_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6419_ _2779_ _2785_ vssd1 vssd1 vccd1 vccd1 _2788_ sky130_fd_sc_hd__nand2_1
Xoutput25 net25 vssd1 vssd1 vccd1 vccd1 la_data_out_23_16[5] sky130_fd_sc_hd__buf_12
XFILLER_0_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_504 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6546__91 clknet_1_0__leaf__2885_ vssd1 vssd1 vccd1 vccd1 net125 sky130_fd_sc_hd__inv_2
XFILLER_39_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6563__106 clknet_1_0__leaf__2887_ vssd1 vssd1 vccd1 vccd1 net140 sky130_fd_sc_hd__inv_2
XFILLER_39_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3982_ _0488_ _3059_ vssd1 vssd1 vccd1 vccd1 _0496_ sky130_fd_sc_hd__nor2_2
XFILLER_62_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6770_ net174 _0229_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[50\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_35_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_478 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5721_ _0897_ _0557_ _2219_ _2220_ _2221_ vssd1 vssd1 vccd1 vccd1 _2222_ sky130_fd_sc_hd__o2111a_1
XFILLER_15_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5652_ _3322_ _3281_ _1153_ egd_top.BitStream_buffer.BS_buffer\[91\] vssd1 vssd1
+ vccd1 vccd1 _2154_ sky130_fd_sc_hd__a22o_1
XFILLER_30_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4603_ _0564_ _0579_ vssd1 vssd1 vccd1 vccd1 _1113_ sky130_fd_sc_hd__nand2_1
X_5583_ _2075_ _2078_ _2081_ _2084_ vssd1 vssd1 vccd1 vccd1 _2085_ sky130_fd_sc_hd__and4_1
X_4534_ _3242_ _3237_ vssd1 vssd1 vccd1 vccd1 _1045_ sky130_fd_sc_hd__nand2_1
XFILLER_7_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4465_ _0581_ egd_top.BitStream_buffer.BS_buffer\[13\] vssd1 vssd1 vccd1 vccd1 _0976_
+ sky130_fd_sc_hd__nand2_1
X_4396_ _0548_ _0537_ vssd1 vssd1 vccd1 vccd1 _0908_ sky130_fd_sc_hd__nand2_1
X_6204_ _2580_ _2581_ vssd1 vssd1 vccd1 vccd1 _2596_ sky130_fd_sc_hd__nand2_2
X_3416_ net7 vssd1 vssd1 vccd1 vccd1 _2966_ sky130_fd_sc_hd__buf_4
X_3347_ net19 vssd1 vssd1 vccd1 vccd1 _2904_ sky130_fd_sc_hd__buf_4
X_6135_ _3023_ _2533_ _2543_ _2551_ vssd1 vssd1 vccd1 vccd1 _0200_ sky130_fd_sc_hd__o211a_1
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6066_ _2511_ _0420_ vssd1 vssd1 vccd1 vccd1 _2513_ sky130_fd_sc_hd__nand2_1
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5017_ _3119_ _3056_ _1523_ vssd1 vssd1 vccd1 vccd1 _1524_ sky130_fd_sc_hd__o21ai_1
XFILLER_85_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5919_ _0510_ _0588_ vssd1 vssd1 vccd1 vccd1 _2419_ sky130_fd_sc_hd__or2_1
XFILLER_1_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4250_ _3282_ _3276_ vssd1 vssd1 vccd1 vccd1 _0763_ sky130_fd_sc_hd__nand2_1
X_4181_ _0692_ _0495_ _0693_ vssd1 vssd1 vccd1 vccd1 _0694_ sky130_fd_sc_hd__o21ai_1
XFILLER_79_194 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6822_ net66 _0281_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.buffer_index\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_35_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6753_ net157 _0212_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[67\]
+ sky130_fd_sc_hd__dfxtp_1
X_3965_ _0477_ _0478_ vssd1 vssd1 vccd1 vccd1 _0479_ sky130_fd_sc_hd__nand2_1
X_5704_ _0955_ _0421_ _2204_ vssd1 vssd1 vccd1 vccd1 _2205_ sky130_fd_sc_hd__o21ai_1
X_3896_ _0393_ _0396_ _0399_ _0400_ _0409_ vssd1 vssd1 vccd1 vccd1 _0410_ sky130_fd_sc_hd__a221oi_1
XFILLER_50_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5635_ _0709_ _3308_ _2134_ _2135_ _2136_ vssd1 vssd1 vccd1 vccd1 _2137_ sky130_fd_sc_hd__o2111a_1
X_5566_ _0621_ egd_top.BitStream_buffer.BS_buffer\[11\] vssd1 vssd1 vccd1 vccd1 _2069_
+ sky130_fd_sc_hd__nand2_1
X_5497_ _3155_ egd_top.BitStream_buffer.BS_buffer\[125\] vssd1 vssd1 vccd1 vccd1 _2000_
+ sky130_fd_sc_hd__nand2_1
X_4517_ _3116_ _3075_ vssd1 vssd1 vccd1 vccd1 _1028_ sky130_fd_sc_hd__nand2_1
XFILLER_2_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4448_ _0955_ _0450_ _0956_ _0957_ _0958_ vssd1 vssd1 vccd1 vccd1 _0959_ sky130_fd_sc_hd__o2111a_1
X_4379_ _0887_ _0450_ _0888_ _0889_ _0890_ vssd1 vssd1 vccd1 vccd1 _0891_ sky130_fd_sc_hd__o2111a_1
X_6118_ _2998_ _2532_ _2528_ _2542_ vssd1 vssd1 vccd1 vccd1 _0208_ sky130_fd_sc_hd__o211a_1
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6049_ _3008_ _2489_ _2501_ _2502_ vssd1 vssd1 vccd1 vccd1 _0237_ sky130_fd_sc_hd__o211a_1
XFILLER_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6592__132 clknet_1_1__leaf__2890_ vssd1 vssd1 vccd1 vccd1 net166 sky130_fd_sc_hd__inv_2
XFILLER_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3750_ _3282_ _3283_ vssd1 vssd1 vccd1 vccd1 _3284_ sky130_fd_sc_hd__nand2_1
X_3681_ _3214_ vssd1 vssd1 vccd1 vccd1 _3215_ sky130_fd_sc_hd__clkbuf_2
XFILLER_9_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5420_ _3074_ _3198_ vssd1 vssd1 vccd1 vccd1 _1924_ sky130_fd_sc_hd__nand2_1
XFILLER_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5351_ _3221_ _0470_ _3227_ _0473_ _1854_ vssd1 vssd1 vccd1 vccd1 _1855_ sky130_fd_sc_hd__a221oi_1
X_4302_ _3009_ _3145_ _0813_ vssd1 vssd1 vccd1 vccd1 _0814_ sky130_fd_sc_hd__o21ai_1
X_5282_ _0388_ _0416_ vssd1 vssd1 vccd1 vccd1 _1787_ sky130_fd_sc_hd__nand2_1
X_4233_ egd_top.BitStream_buffer.BS_buffer\[117\] vssd1 vssd1 vccd1 vccd1 _0746_ sky130_fd_sc_hd__clkbuf_4
XFILLER_59_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6628__5 clknet_1_1__leaf__2893_ vssd1 vssd1 vccd1 vccd1 net39 sky130_fd_sc_hd__inv_2
XFILLER_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4164_ _0578_ _0585_ vssd1 vssd1 vccd1 vccd1 _0677_ sky130_fd_sc_hd__nand2_1
X_4095_ _0608_ vssd1 vssd1 vccd1 vccd1 _0609_ sky130_fd_sc_hd__buf_2
XFILLER_82_112 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6805_ net49 _0264_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[15\]
+ sky130_fd_sc_hd__dfxtp_4
X_4997_ _0346_ _0539_ _0354_ _0542_ _1503_ vssd1 vssd1 vccd1 vccd1 _1504_ sky130_fd_sc_hd__a221oi_1
XFILLER_11_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6736_ net140 _0195_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[100\]
+ sky130_fd_sc_hd__dfxtp_1
X_3948_ _0461_ vssd1 vssd1 vccd1 vccd1 _0462_ sky130_fd_sc_hd__clkinv_2
X_3879_ egd_top.BitStream_buffer.BS_buffer\[44\] vssd1 vssd1 vccd1 vccd1 _0393_ sky130_fd_sc_hd__clkbuf_4
X_5618_ _0503_ egd_top.BitStream_buffer.BS_buffer\[32\] vssd1 vssd1 vccd1 vccd1 _2120_
+ sky130_fd_sc_hd__nand2_1
X_5549_ _0561_ egd_top.BitStream_buffer.BS_buffer\[17\] vssd1 vssd1 vccd1 vccd1 _2052_
+ sky130_fd_sc_hd__nand2_1
XFILLER_78_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4920_ _1426_ _1145_ _1427_ vssd1 vssd1 vccd1 vccd1 _1428_ sky130_fd_sc_hd__o21ai_1
XFILLER_60_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4851_ _0448_ _0439_ _1356_ _1357_ _1358_ vssd1 vssd1 vccd1 vccd1 _1359_ sky130_fd_sc_hd__o2111a_1
X_3802_ _3328_ _3330_ _3335_ vssd1 vssd1 vccd1 vccd1 _3336_ sky130_fd_sc_hd__o21ai_1
X_4782_ _0458_ _0664_ vssd1 vssd1 vccd1 vccd1 _1291_ sky130_fd_sc_hd__nand2_1
X_6521_ _2832_ _2860_ _2881_ vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__o21ai_1
X_3733_ _3248_ _3251_ _3252_ _3255_ _3266_ vssd1 vssd1 vccd1 vccd1 _3267_ sky130_fd_sc_hd__a221oi_1
X_3664_ egd_top.BitStream_buffer.BS_buffer\[119\] vssd1 vssd1 vccd1 vccd1 _3198_ sky130_fd_sc_hd__clkbuf_4
X_6452_ _2810_ _2815_ vssd1 vssd1 vccd1 vccd1 _2816_ sky130_fd_sc_hd__nand2_1
X_5403_ _0767_ _1145_ _1906_ vssd1 vssd1 vccd1 vccd1 _1907_ sky130_fd_sc_hd__o21ai_1
X_3595_ _3127_ _3128_ vssd1 vssd1 vccd1 vccd1 _3129_ sky130_fd_sc_hd__nand2_1
X_6383_ egd_top.BitStream_buffer.BitStream_buffer_output\[9\] _2703_ vssd1 vssd1 vccd1
+ vccd1 _2753_ sky130_fd_sc_hd__nor2_1
X_5334_ _0443_ _0388_ _0655_ _0944_ _1837_ vssd1 vssd1 vccd1 vccd1 _1838_ sky130_fd_sc_hd__a221oi_1
X_5265_ _0462_ _0425_ vssd1 vssd1 vccd1 vccd1 _1770_ sky130_fd_sc_hd__or2_1
XFILLER_87_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4216_ _0728_ vssd1 vssd1 vccd1 vccd1 _0729_ sky130_fd_sc_hd__buf_2
X_5196_ _1673_ _1701_ vssd1 vssd1 vccd1 vccd1 _1702_ sky130_fd_sc_hd__nor2_1
XFILLER_68_451 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4147_ _0420_ _0425_ _0659_ _0421_ vssd1 vssd1 vccd1 vccd1 _0660_ sky130_fd_sc_hd__o22ai_1
XFILLER_83_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4078_ _3052_ _0556_ vssd1 vssd1 vccd1 vccd1 _0592_ sky130_fd_sc_hd__nand2_2
XFILLER_55_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6623__161 clknet_1_1__leaf__2892_ vssd1 vssd1 vccd1 vccd1 net195 sky130_fd_sc_hd__inv_2
XFILLER_43_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6719_ net123 _0178_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.pc_previous\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_50_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3380_ _2933_ vssd1 vssd1 vccd1 vccd1 _2934_ sky130_fd_sc_hd__clkbuf_4
X_5050_ _1003_ _3319_ vssd1 vssd1 vccd1 vccd1 _1557_ sky130_fd_sc_hd__or2_1
X_4001_ egd_top.BitStream_buffer.BS_buffer\[22\] vssd1 vssd1 vccd1 vccd1 _0515_ sky130_fd_sc_hd__clkbuf_4
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0__f__2887_ clknet_0__2887_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__2887_
+ sky130_fd_sc_hd__clkbuf_16
X_5952_ _2901_ vssd1 vssd1 vccd1 vccd1 _2446_ sky130_fd_sc_hd__buf_2
XFILLER_37_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4903_ _3047_ _0714_ vssd1 vssd1 vccd1 vccd1 _1411_ sky130_fd_sc_hd__nand2_1
X_5883_ _0887_ _0403_ _2382_ vssd1 vssd1 vccd1 vccd1 _2383_ sky130_fd_sc_hd__o21ai_1
XFILLER_60_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4834_ _0377_ _0407_ vssd1 vssd1 vccd1 vccd1 _1342_ sky130_fd_sc_hd__nand2_1
X_4765_ _0637_ _0350_ _1273_ vssd1 vssd1 vccd1 vccd1 _1274_ sky130_fd_sc_hd__o21ai_1
X_3716_ _3249_ vssd1 vssd1 vccd1 vccd1 _3250_ sky130_fd_sc_hd__buf_2
X_6504_ _2862_ _2685_ _2865_ vssd1 vssd1 vccd1 vccd1 _2866_ sky130_fd_sc_hd__nand3_1
X_4696_ _3026_ _1205_ vssd1 vssd1 vccd1 vccd1 _1206_ sky130_fd_sc_hd__nor2_1
X_3647_ _3076_ _3134_ vssd1 vssd1 vccd1 vccd1 _3181_ sky130_fd_sc_hd__and2_1
X_6435_ _2690_ _2684_ _2700_ vssd1 vssd1 vccd1 vccd1 _2800_ sky130_fd_sc_hd__and3_1
XFILLER_20_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3578_ _3041_ _3111_ vssd1 vssd1 vccd1 vccd1 _3112_ sky130_fd_sc_hd__nor2_2
X_6366_ _2736_ vssd1 vssd1 vccd1 vccd1 _2737_ sky130_fd_sc_hd__inv_2
XFILLER_88_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5317_ _1128_ _0613_ vssd1 vssd1 vccd1 vccd1 _1822_ sky130_fd_sc_hd__or2_1
X_6297_ _2642_ _2667_ vssd1 vssd1 vccd1 vccd1 _2668_ sky130_fd_sc_hd__nor2_1
X_5248_ _1741_ _1745_ _1749_ _1752_ vssd1 vssd1 vccd1 vccd1 _1753_ sky130_fd_sc_hd__and4_1
XFILLER_29_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5179_ _1676_ _1679_ _1681_ _1684_ vssd1 vssd1 vccd1 vccd1 _1685_ sky130_fd_sc_hd__and4_1
XFILLER_68_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4550_ _3162_ egd_top.BitStream_buffer.BS_buffer\[116\] vssd1 vssd1 vccd1 vccd1 _1061_
+ sky130_fd_sc_hd__nand2_1
X_4481_ _0503_ _0509_ vssd1 vssd1 vccd1 vccd1 _0992_ sky130_fd_sc_hd__nand2_1
X_3501_ egd_top.BitStream_buffer.pc\[4\] _2932_ _3034_ vssd1 vssd1 vccd1 vccd1 _3035_
+ sky130_fd_sc_hd__or3_2
X_6220_ _2979_ _2602_ _2570_ _2605_ vssd1 vssd1 vccd1 vccd1 _0175_ sky130_fd_sc_hd__o211a_1
X_3432_ _2976_ _2980_ vssd1 vssd1 vccd1 vccd1 _2981_ sky130_fd_sc_hd__nand2_1
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3363_ _2915_ _2916_ vssd1 vssd1 vccd1 vccd1 _2917_ sky130_fd_sc_hd__and2_1
X_6151_ _2988_ _2554_ _2558_ _2562_ vssd1 vssd1 vccd1 vccd1 _0195_ sky130_fd_sc_hd__o211a_1
X_5102_ _1606_ _1607_ vssd1 vssd1 vccd1 vccd1 _1608_ sky130_fd_sc_hd__nand2_1
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6082_ _2517_ _0965_ vssd1 vssd1 vccd1 vccd1 _2522_ sky130_fd_sc_hd__nand2_1
X_5033_ _3163_ _0744_ vssd1 vssd1 vccd1 vccd1 _1540_ sky130_fd_sc_hd__nand2_1
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5935_ _2974_ _2901_ _2433_ vssd1 vssd1 vccd1 vccd1 _2434_ sky130_fd_sc_hd__and3_1
X_5866_ _3144_ _0562_ vssd1 vssd1 vccd1 vccd1 _2366_ sky130_fd_sc_hd__nand2_1
XFILLER_33_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4817_ _0609_ _0498_ vssd1 vssd1 vccd1 vccd1 _1326_ sky130_fd_sc_hd__nand2_1
XFILLER_21_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5797_ _0713_ _3330_ _2297_ vssd1 vssd1 vccd1 vccd1 _2298_ sky130_fd_sc_hd__o21ai_1
X_4748_ _1149_ _1145_ _1256_ vssd1 vssd1 vccd1 vccd1 _1257_ sky130_fd_sc_hd__o21ai_1
X_4679_ _3015_ _3145_ _1188_ vssd1 vssd1 vccd1 vccd1 _1189_ sky130_fd_sc_hd__o21ai_1
X_6418_ _2770_ _2786_ vssd1 vssd1 vccd1 vccd1 _2787_ sky130_fd_sc_hd__nand2_1
Xoutput26 net26 vssd1 vssd1 vccd1 vccd1 la_data_out_23_16[6] sky130_fd_sc_hd__buf_12
XFILLER_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6349_ _2717_ _2719_ vssd1 vssd1 vccd1 vccd1 _2720_ sky130_fd_sc_hd__nand2_1
XFILLER_88_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_56 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3981_ _0494_ vssd1 vssd1 vccd1 vccd1 _0495_ sky130_fd_sc_hd__buf_2
XFILLER_62_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5720_ _0492_ _0570_ vssd1 vssd1 vccd1 vccd1 _2221_ sky130_fd_sc_hd__or2_1
XFILLER_62_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5651_ _0837_ _3216_ _3302_ _3220_ _2152_ vssd1 vssd1 vccd1 vccd1 _2153_ sky130_fd_sc_hd__a221oi_1
XFILLER_30_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4602_ _1096_ _1111_ vssd1 vssd1 vccd1 vccd1 _1112_ sky130_fd_sc_hd__and2_1
X_5582_ _0454_ _0395_ _0398_ _0461_ _2083_ vssd1 vssd1 vccd1 vccd1 _2084_ sky130_fd_sc_hd__a221oi_1
XFILLER_7_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4533_ _3232_ egd_top.BitStream_buffer.BS_buffer\[69\] vssd1 vssd1 vccd1 vccd1 _1044_
+ sky130_fd_sc_hd__nand2_1
X_4464_ _0577_ egd_top.BitStream_buffer.BS_buffer\[11\] vssd1 vssd1 vccd1 vccd1 _0975_
+ sky130_fd_sc_hd__nand2_1
X_6203_ _2595_ vssd1 vssd1 vccd1 vccd1 _0180_ sky130_fd_sc_hd__inv_2
X_4395_ _0540_ vssd1 vssd1 vccd1 vccd1 _0907_ sky130_fd_sc_hd__inv_2
X_3415_ _2965_ _2949_ _2902_ vssd1 vssd1 vccd1 vccd1 _0314_ sky130_fd_sc_hd__o21ai_1
X_3346_ net34 vssd1 vssd1 vccd1 vccd1 _2903_ sky130_fd_sc_hd__inv_2
X_6134_ _2531_ _3277_ vssd1 vssd1 vccd1 vccd1 _2551_ sky130_fd_sc_hd__nand2_1
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6065_ _2966_ _2510_ _2501_ _2512_ vssd1 vssd1 vccd1 vccd1 _0231_ sky130_fd_sc_hd__o211a_1
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5016_ _3061_ _3109_ vssd1 vssd1 vccd1 vccd1 _1523_ sky130_fd_sc_hd__nand2_1
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5918_ _0582_ _0519_ vssd1 vssd1 vccd1 vccd1 _2418_ sky130_fd_sc_hd__nand2_1
XFILLER_41_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5849_ _3291_ egd_top.BitStream_buffer.BS_buffer\[96\] vssd1 vssd1 vccd1 vccd1 _2349_
+ sky130_fd_sc_hd__nand2_1
XFILLER_1_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4180_ _0497_ _0502_ vssd1 vssd1 vccd1 vccd1 _0693_ sky130_fd_sc_hd__nand2_1
XFILLER_82_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6821_ net65 _0280_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.buffer_index\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_90_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3964_ egd_top.BitStream_buffer.BS_buffer\[62\] vssd1 vssd1 vccd1 vccd1 _0478_ sky130_fd_sc_hd__clkbuf_4
X_6752_ net156 _0211_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[68\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_23_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5703_ _0887_ _0424_ vssd1 vssd1 vccd1 vccd1 _2204_ sky130_fd_sc_hd__or2_1
X_3895_ _0401_ _0403_ _0408_ vssd1 vssd1 vccd1 vccd1 _0409_ sky130_fd_sc_hd__o21ai_1
X_5634_ _1169_ _3319_ vssd1 vssd1 vccd1 vccd1 _2136_ sky130_fd_sc_hd__or2_1
X_5565_ _2039_ _2067_ vssd1 vssd1 vccd1 vccd1 _2068_ sky130_fd_sc_hd__nor2_1
X_5496_ _3167_ egd_top.BitStream_buffer.BS_buffer\[123\] vssd1 vssd1 vccd1 vccd1 _1999_
+ sky130_fd_sc_hd__nand2_1
X_4516_ _3112_ _3070_ vssd1 vssd1 vccd1 vccd1 _1027_ sky130_fd_sc_hd__nand2_1
XFILLER_2_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4447_ _0647_ _0463_ vssd1 vssd1 vccd1 vccd1 _0958_ sky130_fd_sc_hd__or2_1
X_6686__58 clknet_1_0__leaf__2898_ vssd1 vssd1 vccd1 vccd1 net92 sky130_fd_sc_hd__inv_2
XFILLER_85_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6117_ _2538_ _1430_ vssd1 vssd1 vccd1 vccd1 _2542_ sky130_fd_sc_hd__nand2_1
X_4378_ _0448_ _0464_ vssd1 vssd1 vccd1 vccd1 _0890_ sky130_fd_sc_hd__or2_1
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6048_ _2494_ _0936_ vssd1 vssd1 vccd1 vccd1 _2502_ sky130_fd_sc_hd__nand2_1
XFILLER_37_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_24 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3680_ _3090_ _3213_ vssd1 vssd1 vccd1 vccd1 _3214_ sky130_fd_sc_hd__and2_1
XFILLER_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5350_ _0759_ _2935_ _1853_ vssd1 vssd1 vccd1 vccd1 _1854_ sky130_fd_sc_hd__o21ai_1
X_4301_ _3148_ _3138_ vssd1 vssd1 vccd1 vccd1 _0813_ sky130_fd_sc_hd__nand2_1
X_5281_ _0869_ _0360_ _0363_ _0393_ _1785_ vssd1 vssd1 vccd1 vccd1 _1786_ sky130_fd_sc_hd__a221oi_1
X_4232_ _3198_ _3193_ _3196_ _0744_ vssd1 vssd1 vccd1 vccd1 _0745_ sky130_fd_sc_hd__a22o_1
X_4163_ egd_top.BitStream_buffer.BS_buffer\[12\] vssd1 vssd1 vccd1 vccd1 _0676_ sky130_fd_sc_hd__inv_2
XFILLER_67_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4094_ _0559_ _3077_ vssd1 vssd1 vccd1 vccd1 _0608_ sky130_fd_sc_hd__nor2_2
XFILLER_82_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4996_ _0940_ _0546_ _1502_ vssd1 vssd1 vccd1 vccd1 _1503_ sky130_fd_sc_hd__o21ai_1
XFILLER_63_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6804_ net48 _0263_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[16\]
+ sky130_fd_sc_hd__dfxtp_4
X_3947_ egd_top.BitStream_buffer.BS_buffer\[57\] vssd1 vssd1 vccd1 vccd1 _0461_ sky130_fd_sc_hd__clkbuf_4
X_6735_ net139 _0194_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[101\]
+ sky130_fd_sc_hd__dfxtp_1
X_3878_ _0375_ _0378_ _0379_ _0382_ _0391_ vssd1 vssd1 vccd1 vccd1 _0392_ sky130_fd_sc_hd__a221oi_1
X_5617_ _0702_ _0494_ _2116_ _2117_ _2118_ vssd1 vssd1 vccd1 vccd1 _2119_ sky130_fd_sc_hd__o2111a_1
X_5548_ _2042_ _2045_ _2047_ _2050_ vssd1 vssd1 vccd1 vccd1 _2051_ sky130_fd_sc_hd__and4_1
XFILLER_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5479_ _3232_ _3272_ vssd1 vssd1 vccd1 vccd1 _1982_ sky130_fd_sc_hd__nand2_1
XFILLER_78_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_382 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6600__140 clknet_1_1__leaf__2890_ vssd1 vssd1 vccd1 vccd1 net174 sky130_fd_sc_hd__inv_2
XFILLER_6_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6665__39 clknet_1_1__leaf__2896_ vssd1 vssd1 vccd1 vccd1 net73 sky130_fd_sc_hd__inv_2
XFILLER_77_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6599__139 clknet_1_1__leaf__2890_ vssd1 vssd1 vccd1 vccd1 net173 sky130_fd_sc_hd__inv_2
XFILLER_33_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4850_ _0435_ _0471_ vssd1 vssd1 vccd1 vccd1 _1358_ sky130_fd_sc_hd__nand2_1
XFILLER_45_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3801_ _3333_ _3334_ vssd1 vssd1 vccd1 vccd1 _3335_ sky130_fd_sc_hd__nand2_1
X_4781_ _0453_ _0471_ vssd1 vssd1 vccd1 vccd1 _1290_ sky130_fd_sc_hd__nand2_1
X_6520_ _2877_ _2878_ _2880_ vssd1 vssd1 vccd1 vccd1 _2881_ sky130_fd_sc_hd__nand3_1
X_6630__7 clknet_1_0__leaf__2893_ vssd1 vssd1 vccd1 vccd1 net41 sky130_fd_sc_hd__inv_2
X_3732_ _3257_ _3260_ _3265_ vssd1 vssd1 vccd1 vccd1 _3266_ sky130_fd_sc_hd__o21ai_1
X_3663_ _3196_ vssd1 vssd1 vccd1 vccd1 _3197_ sky130_fd_sc_hd__buf_6
X_6451_ _2812_ _2813_ _2673_ _2669_ _2814_ vssd1 vssd1 vccd1 vccd1 _2815_ sky130_fd_sc_hd__o32a_1
X_5402_ _3224_ _0837_ vssd1 vssd1 vccd1 vccd1 _1906_ sky130_fd_sc_hd__nand2_1
X_6382_ _2688_ _2751_ _2717_ vssd1 vssd1 vccd1 vccd1 _2752_ sky130_fd_sc_hd__o21ai_1
X_3594_ egd_top.BitStream_buffer.BS_buffer\[104\] vssd1 vssd1 vccd1 vccd1 _3128_ sky130_fd_sc_hd__clkbuf_4
X_5333_ _0879_ _0380_ _1836_ vssd1 vssd1 vccd1 vccd1 _1837_ sky130_fd_sc_hd__o21ai_1
X_5264_ _1721_ _1737_ _1753_ _1768_ vssd1 vssd1 vccd1 vccd1 _1769_ sky130_fd_sc_hd__and4_1
XFILLER_87_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5195_ _1685_ _1700_ vssd1 vssd1 vccd1 vccd1 _1701_ sky130_fd_sc_hd__nand2_1
X_4215_ _3069_ vssd1 vssd1 vccd1 vccd1 _0728_ sky130_fd_sc_hd__inv_2
XFILLER_68_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4146_ egd_top.BitStream_buffer.BS_buffer\[50\] vssd1 vssd1 vccd1 vccd1 _0659_ sky130_fd_sc_hd__inv_2
XFILLER_55_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4077_ egd_top.BitStream_buffer.BS_buffer\[2\] vssd1 vssd1 vccd1 vccd1 _0591_ sky130_fd_sc_hd__inv_2
XFILLER_24_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4979_ _0453_ _0664_ vssd1 vssd1 vccd1 vccd1 _1486_ sky130_fd_sc_hd__nand2_1
X_6718_ net122 _0177_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.pc_previous\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_3_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4000_ _0513_ vssd1 vssd1 vccd1 vccd1 _0514_ sky130_fd_sc_hd__buf_4
XFILLER_37_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6607__146 clknet_1_1__leaf__2891_ vssd1 vssd1 vccd1 vccd1 net180 sky130_fd_sc_hd__inv_2
XFILLER_37_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0__f__2886_ clknet_0__2886_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__2886_
+ sky130_fd_sc_hd__clkbuf_16
X_5951_ _2979_ _2442_ _3002_ _2445_ vssd1 vssd1 vccd1 vccd1 _0278_ sky130_fd_sc_hd__o211a_1
X_4902_ _3038_ egd_top.BitStream_buffer.BS_buffer\[102\] vssd1 vssd1 vccd1 vccd1 _1410_
+ sky130_fd_sc_hd__nand2_1
X_5882_ _0406_ _0467_ vssd1 vssd1 vccd1 vccd1 _2382_ sky130_fd_sc_hd__nand2_1
X_4833_ _0375_ _0359_ _0362_ _0379_ _1340_ vssd1 vssd1 vccd1 vccd1 _1341_ sky130_fd_sc_hd__a221oi_1
XFILLER_21_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4764_ _0353_ _0869_ vssd1 vssd1 vccd1 vccd1 _1273_ sky130_fd_sc_hd__nand2_1
X_3715_ _3110_ _3212_ vssd1 vssd1 vccd1 vccd1 _3249_ sky130_fd_sc_hd__and2_1
X_6503_ _2864_ _2827_ vssd1 vssd1 vccd1 vccd1 _2865_ sky130_fd_sc_hd__nand2_1
X_4695_ _1141_ _1203_ _1204_ vssd1 vssd1 vccd1 vccd1 _1205_ sky130_fd_sc_hd__nand3_1
X_6434_ _2798_ _2643_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.exp_golomb_len\[2\]
+ sky130_fd_sc_hd__nor2_1
X_3646_ _3179_ vssd1 vssd1 vccd1 vccd1 _3180_ sky130_fd_sc_hd__buf_4
X_3577_ _3110_ vssd1 vssd1 vccd1 vccd1 _3111_ sky130_fd_sc_hd__clkinv_2
X_6365_ net17 _2922_ vssd1 vssd1 vccd1 vccd1 _2736_ sky130_fd_sc_hd__nor2_1
X_5316_ _0606_ _0505_ vssd1 vssd1 vccd1 vccd1 _1821_ sky130_fd_sc_hd__nand2_1
X_6296_ _2637_ _2625_ vssd1 vssd1 vccd1 vccd1 _2667_ sky130_fd_sc_hd__nand2_1
X_5247_ _0772_ _3282_ _3334_ _1153_ _1751_ vssd1 vssd1 vccd1 vccd1 _1752_ sky130_fd_sc_hd__a221oi_1
XFILLER_75_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5178_ _0354_ _0539_ _0347_ _0542_ _1683_ vssd1 vssd1 vccd1 vccd1 _1684_ sky130_fd_sc_hd__a221oi_1
XFILLER_56_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4129_ egd_top.BitStream_buffer.BS_buffer\[47\] vssd1 vssd1 vccd1 vccd1 _0642_ sky130_fd_sc_hd__clkbuf_4
XFILLER_83_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_499 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_94 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3500_ egd_top.BitStream_buffer.pc\[5\] vssd1 vssd1 vccd1 vccd1 _3034_ sky130_fd_sc_hd__inv_2
XFILLER_51_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4480_ _0513_ _0527_ vssd1 vssd1 vccd1 vccd1 _0991_ sky130_fd_sc_hd__nand2_1
X_3431_ egd_top.BitStream_buffer.BS_buffer\[113\] vssd1 vssd1 vccd1 vccd1 _2980_ sky130_fd_sc_hd__clkinv_2
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3362_ net30 vssd1 vssd1 vccd1 vccd1 _2916_ sky130_fd_sc_hd__inv_2
X_6150_ _2561_ _0796_ vssd1 vssd1 vccd1 vccd1 _2562_ sky130_fd_sc_hd__nand2_1
X_5101_ _3168_ _0744_ vssd1 vssd1 vccd1 vccd1 _1607_ sky130_fd_sc_hd__nand2_1
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6081_ _2998_ _2510_ _2516_ _2521_ vssd1 vssd1 vccd1 vccd1 _0224_ sky130_fd_sc_hd__o211a_1
XFILLER_85_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5032_ _0792_ _3137_ _0930_ _3141_ _1538_ vssd1 vssd1 vccd1 vccd1 _1539_ sky130_fd_sc_hd__a221oi_1
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5934_ _2972_ _2967_ vssd1 vssd1 vccd1 vccd1 _2433_ sky130_fd_sc_hd__nand2_1
X_5865_ _3136_ _0579_ vssd1 vssd1 vccd1 vccd1 _2365_ sky130_fd_sc_hd__nand2_1
X_4816_ _0606_ egd_top.BitStream_buffer.BS_buffer\[17\] vssd1 vssd1 vccd1 vccd1 _1325_
+ sky130_fd_sc_hd__nand2_1
XFILLER_21_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5796_ _3333_ _0716_ vssd1 vssd1 vccd1 vccd1 _2297_ sky130_fd_sc_hd__nand2_1
X_4747_ _3223_ _3252_ vssd1 vssd1 vccd1 vccd1 _1256_ sky130_fd_sc_hd__nand2_1
X_4678_ _3148_ _3177_ vssd1 vssd1 vccd1 vccd1 _1188_ sky130_fd_sc_hd__nand2_1
X_3629_ _3162_ vssd1 vssd1 vccd1 vccd1 _3163_ sky130_fd_sc_hd__buf_6
X_6417_ _2779_ _2785_ _2926_ vssd1 vssd1 vccd1 vccd1 _2786_ sky130_fd_sc_hd__a21oi_1
Xoutput27 net27 vssd1 vssd1 vccd1 vccd1 la_data_out_23_16[7] sky130_fd_sc_hd__buf_12
X_6348_ _2687_ _2718_ vssd1 vssd1 vccd1 vccd1 _2719_ sky130_fd_sc_hd__nand2_1
XFILLER_88_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6279_ _2648_ _2649_ vssd1 vssd1 vccd1 vccd1 _2650_ sky130_fd_sc_hd__nand2_1
XFILLER_88_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3980_ _0493_ vssd1 vssd1 vccd1 vccd1 _0494_ sky130_fd_sc_hd__clkinv_2
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5650_ _1007_ _1145_ _2151_ vssd1 vssd1 vccd1 vccd1 _2152_ sky130_fd_sc_hd__o21ai_1
XFILLER_87_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4601_ _1100_ _1104_ _1107_ _1110_ vssd1 vssd1 vccd1 vccd1 _1111_ sky130_fd_sc_hd__and4_1
XFILLER_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6537__82 clknet_1_1__leaf__2885_ vssd1 vssd1 vccd1 vccd1 net116 sky130_fd_sc_hd__inv_2
X_5581_ _0448_ _0402_ _2082_ vssd1 vssd1 vccd1 vccd1 _2083_ sky130_fd_sc_hd__o21ai_1
X_4532_ egd_top.BitStream_buffer.BS_buffer\[68\] vssd1 vssd1 vccd1 vccd1 _1043_ sky130_fd_sc_hd__clkinv_2
X_4463_ _0679_ _0557_ _0971_ _0972_ _0973_ vssd1 vssd1 vccd1 vccd1 _0974_ sky130_fd_sc_hd__o2111a_1
X_6202_ _2902_ egd_top.BitStream_buffer.pc\[3\] vssd1 vssd1 vccd1 vccd1 _2595_ sky130_fd_sc_hd__nand2_1
X_6552__96 clknet_1_1__leaf__2886_ vssd1 vssd1 vccd1 vccd1 net130 sky130_fd_sc_hd__inv_2
X_3414_ _2964_ vssd1 vssd1 vccd1 vccd1 _2965_ sky130_fd_sc_hd__buf_2
X_4394_ _0699_ _0534_ _0543_ _0526_ _0905_ vssd1 vssd1 vccd1 vccd1 _0906_ sky130_fd_sc_hd__o221a_1
X_6133_ _3020_ _2533_ _2543_ _2550_ vssd1 vssd1 vccd1 vccd1 _0201_ sky130_fd_sc_hd__o211a_1
X_3345_ net34 _2900_ _2902_ vssd1 vssd1 vccd1 vccd1 _0321_ sky130_fd_sc_hd__o21a_1
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6064_ _2511_ _0423_ vssd1 vssd1 vccd1 vccd1 _2512_ sky130_fd_sc_hd__nand2_1
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5015_ _1494_ _1521_ vssd1 vssd1 vccd1 vccd1 _1522_ sky130_fd_sc_hd__nor2_1
XFILLER_38_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5917_ _0578_ _0515_ vssd1 vssd1 vccd1 vccd1 _2417_ sky130_fd_sc_hd__nand2_1
XFILLER_13_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5848_ _0784_ _3298_ vssd1 vssd1 vccd1 vccd1 _2348_ sky130_fd_sc_hd__or2_1
X_5779_ _3243_ _3272_ vssd1 vssd1 vccd1 vccd1 _2280_ sky130_fd_sc_hd__nand2_1
XFILLER_5_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6700__71 clknet_1_1__leaf__2899_ vssd1 vssd1 vccd1 vccd1 net105 sky130_fd_sc_hd__inv_2
XFILLER_76_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_358 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6820_ net64 _0279_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[0\]
+ sky130_fd_sc_hd__dfxtp_2
X_6751_ net155 _0210_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[69\]
+ sky130_fd_sc_hd__dfxtp_1
X_3963_ _0476_ vssd1 vssd1 vccd1 vccd1 _0477_ sky130_fd_sc_hd__clkbuf_4
X_5702_ _2193_ _2196_ _2199_ _2202_ vssd1 vssd1 vccd1 vccd1 _2203_ sky130_fd_sc_hd__and4_1
X_3894_ _0406_ _0407_ vssd1 vssd1 vccd1 vccd1 _0408_ sky130_fd_sc_hd__nand2_1
XFILLER_31_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5633_ _3314_ _3028_ vssd1 vssd1 vccd1 vccd1 _2135_ sky130_fd_sc_hd__nand2_1
X_5564_ _2051_ _2066_ vssd1 vssd1 vccd1 vccd1 _2067_ sky130_fd_sc_hd__nand2_1
XFILLER_12_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4515_ _3126_ _3118_ vssd1 vssd1 vccd1 vccd1 _1026_ sky130_fd_sc_hd__nand2_1
X_5495_ _3159_ _0741_ vssd1 vssd1 vccd1 vccd1 _1998_ sky130_fd_sc_hd__nand2_1
X_4446_ _0458_ _0471_ vssd1 vssd1 vccd1 vccd1 _0957_ sky130_fd_sc_hd__nand2_1
X_4377_ _0458_ _0467_ vssd1 vssd1 vccd1 vccd1 _0889_ sky130_fd_sc_hd__nand2_1
X_6116_ _2995_ _2532_ _2528_ _2541_ vssd1 vssd1 vccd1 vccd1 _0209_ sky130_fd_sc_hd__o211a_1
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6047_ _2904_ vssd1 vssd1 vccd1 vccd1 _2501_ sky130_fd_sc_hd__buf_2
XFILLER_81_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6531__77 clknet_1_1__leaf__2884_ vssd1 vssd1 vccd1 vccd1 net111 sky130_fd_sc_hd__inv_2
XFILLER_78_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4300_ _0799_ _0803_ _0807_ _0811_ vssd1 vssd1 vccd1 vccd1 _0812_ sky130_fd_sc_hd__and4_1
X_5280_ _0936_ _0368_ _1784_ vssd1 vssd1 vccd1 vccd1 _1785_ sky130_fd_sc_hd__o21ai_1
XFILLER_87_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4231_ egd_top.BitStream_buffer.BS_buffer\[120\] vssd1 vssd1 vccd1 vccd1 _0744_ sky130_fd_sc_hd__clkbuf_4
XFILLER_67_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4162_ _0670_ _0558_ _0671_ _0672_ _0674_ vssd1 vssd1 vccd1 vccd1 _0675_ sky130_fd_sc_hd__o2111a_1
X_4093_ _0606_ egd_top.BitStream_buffer.BS_buffer\[12\] vssd1 vssd1 vccd1 vccd1 _0607_
+ sky130_fd_sc_hd__nand2_1
XFILLER_67_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6691__62 clknet_1_0__leaf__2899_ vssd1 vssd1 vccd1 vccd1 net96 sky130_fd_sc_hd__inv_2
XFILLER_67_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4995_ _0548_ _0364_ vssd1 vssd1 vccd1 vccd1 _1502_ sky130_fd_sc_hd__nand2_1
XFILLER_23_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6803_ net47 _0262_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[17\]
+ sky130_fd_sc_hd__dfxtp_4
X_3946_ _0458_ _0459_ vssd1 vssd1 vccd1 vccd1 _0460_ sky130_fd_sc_hd__nand2_1
X_6576__118 clknet_1_1__leaf__2888_ vssd1 vssd1 vccd1 vccd1 net152 sky130_fd_sc_hd__inv_2
X_6734_ net138 _0193_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[102\]
+ sky130_fd_sc_hd__dfxtp_2
X_3877_ _0383_ _0385_ _0390_ vssd1 vssd1 vccd1 vccd1 _0391_ sky130_fd_sc_hd__o21ai_1
X_5616_ _0489_ egd_top.BitStream_buffer.BS_buffer\[29\] vssd1 vssd1 vccd1 vccd1 _2118_
+ sky130_fd_sc_hd__nand2_1
X_5547_ _0379_ _0539_ _0389_ _0542_ _2049_ vssd1 vssd1 vccd1 vccd1 _2050_ sky130_fd_sc_hd__a221oi_1
XFILLER_2_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5478_ _3242_ egd_top.BitStream_buffer.BS_buffer\[75\] vssd1 vssd1 vccd1 vccd1 _1981_
+ sky130_fd_sc_hd__nand2_1
X_4429_ _0337_ vssd1 vssd1 vccd1 vccd1 _0940_ sky130_fd_sc_hd__inv_2
XFILLER_86_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_114 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4780_ _0436_ _0415_ _0454_ _0419_ _1288_ vssd1 vssd1 vccd1 vccd1 _1289_ sky130_fd_sc_hd__a221oi_1
X_3800_ egd_top.BitStream_buffer.BS_buffer\[88\] vssd1 vssd1 vccd1 vccd1 _3334_ sky130_fd_sc_hd__clkbuf_4
X_3731_ _3263_ _3264_ vssd1 vssd1 vccd1 vccd1 _3265_ sky130_fd_sc_hd__nand2_1
X_3662_ _3195_ vssd1 vssd1 vccd1 vccd1 _3196_ sky130_fd_sc_hd__clkbuf_2
XFILLER_9_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6450_ _2712_ _2702_ _2631_ vssd1 vssd1 vccd1 vccd1 _2814_ sky130_fd_sc_hd__a21o_1
X_3593_ _3126_ vssd1 vssd1 vccd1 vccd1 _3127_ sky130_fd_sc_hd__buf_2
X_6381_ _1705_ _2686_ vssd1 vssd1 vccd1 vccd1 _2751_ sky130_fd_sc_hd__nor2_1
X_5401_ _3268_ _3233_ _3236_ _3272_ _1904_ vssd1 vssd1 vccd1 vccd1 _1905_ sky130_fd_sc_hd__a221oi_2
X_5332_ _0378_ _0412_ vssd1 vssd1 vccd1 vccd1 _1836_ sky130_fd_sc_hd__nand2_1
XFILLER_87_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5263_ _1760_ _1764_ _1767_ vssd1 vssd1 vccd1 vccd1 _1768_ sky130_fd_sc_hd__and3_1
X_5194_ _1689_ _1693_ _1695_ _1699_ vssd1 vssd1 vccd1 vccd1 _1700_ sky130_fd_sc_hd__and4_1
X_4214_ egd_top.BitStream_buffer.BS_buffer\[109\] vssd1 vssd1 vccd1 vccd1 _0727_ sky130_fd_sc_hd__inv_2
X_4145_ _0653_ _0438_ _0654_ _0656_ _0657_ vssd1 vssd1 vccd1 vccd1 _0658_ sky130_fd_sc_hd__o2111a_1
XFILLER_83_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4076_ _0574_ _0576_ _0580_ _0584_ _0589_ vssd1 vssd1 vccd1 vccd1 _0590_ sky130_fd_sc_hd__o2111a_1
XFILLER_55_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4978_ _0471_ _0432_ _0435_ _0478_ _1484_ vssd1 vssd1 vccd1 vccd1 _1485_ sky130_fd_sc_hd__a221oi_1
X_6717_ net121 _0176_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[80\]
+ sky130_fd_sc_hd__dfxtp_1
X_3929_ egd_top.BitStream_buffer.BS_buffer\[52\] vssd1 vssd1 vccd1 vccd1 _0443_ sky130_fd_sc_hd__clkbuf_4
XFILLER_3_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6670__43 clknet_1_0__leaf__2897_ vssd1 vssd1 vccd1 vccd1 net77 sky130_fd_sc_hd__inv_2
XFILLER_46_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6559__102 clknet_1_1__leaf__2887_ vssd1 vssd1 vccd1 vccd1 net136 sky130_fd_sc_hd__inv_2
XFILLER_91_88 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0__f__2885_ clknet_0__2885_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__2885_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_1_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5950_ _2443_ _0594_ vssd1 vssd1 vccd1 vccd1 _2445_ sky130_fd_sc_hd__nand2_1
XFILLER_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4901_ _1397_ _1401_ _1405_ _1408_ vssd1 vssd1 vccd1 vccd1 _1409_ sky130_fd_sc_hd__and4_1
XFILLER_52_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5881_ _0874_ _0360_ _0363_ _0948_ _2380_ vssd1 vssd1 vccd1 vccd1 _2381_ sky130_fd_sc_hd__a221oi_2
XFILLER_33_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4832_ _0348_ _0367_ _1339_ vssd1 vssd1 vccd1 vccd1 _1340_ sky130_fd_sc_hd__o21ai_1
XFILLER_60_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4763_ _1222_ _1238_ _1255_ _1271_ vssd1 vssd1 vccd1 vccd1 _1272_ sky130_fd_sc_hd__and4_1
X_4694_ _0622_ _0566_ vssd1 vssd1 vccd1 vccd1 _1204_ sky130_fd_sc_hd__nand2_1
X_6502_ _2863_ _2849_ vssd1 vssd1 vccd1 vccd1 _2864_ sky130_fd_sc_hd__nor2_1
X_3714_ egd_top.BitStream_buffer.BS_buffer\[74\] vssd1 vssd1 vccd1 vccd1 _3248_ sky130_fd_sc_hd__clkbuf_4
X_6433_ _2799_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.exp_golomb_len\[1\]
+ sky130_fd_sc_hd__inv_2
X_3645_ _3178_ vssd1 vssd1 vccd1 vccd1 _3179_ sky130_fd_sc_hd__clkbuf_2
XFILLER_20_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3576_ _3051_ _3031_ egd_top.BitStream_buffer.pc\[3\] vssd1 vssd1 vccd1 vccd1 _3110_
+ sky130_fd_sc_hd__and3_2
X_6364_ _2722_ _2734_ vssd1 vssd1 vccd1 vccd1 _2735_ sky130_fd_sc_hd__nand2_1
X_5315_ _0609_ _0509_ vssd1 vssd1 vccd1 vccd1 _1820_ sky130_fd_sc_hd__nand2_1
X_6295_ _2665_ _2635_ vssd1 vssd1 vccd1 vccd1 _2666_ sky130_fd_sc_hd__nand2_1
X_5246_ _0771_ _3273_ _1750_ vssd1 vssd1 vccd1 vccd1 _1751_ sky130_fd_sc_hd__o21ai_1
X_5177_ _1084_ _0546_ _1682_ vssd1 vssd1 vccd1 vccd1 _1683_ sky130_fd_sc_hd__o21ai_1
XFILLER_68_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4128_ _0637_ _0384_ _0638_ _0639_ _0640_ vssd1 vssd1 vccd1 vccd1 _0641_ sky130_fd_sc_hd__o2111a_1
X_4059_ _0554_ _0558_ _0563_ _0567_ _0572_ vssd1 vssd1 vccd1 vccd1 _0573_ sky130_fd_sc_hd__o2111a_1
XFILLER_71_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3430_ net6 vssd1 vssd1 vccd1 vccd1 _2979_ sky130_fd_sc_hd__buf_4
X_3361_ net29 net28 vssd1 vssd1 vccd1 vccd1 _2915_ sky130_fd_sc_hd__nor2_1
X_5100_ _3163_ _3149_ vssd1 vssd1 vccd1 vccd1 _1606_ sky130_fd_sc_hd__nand2_1
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6080_ _2517_ _0883_ vssd1 vssd1 vccd1 vccd1 _2521_ sky130_fd_sc_hd__nand2_1
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5031_ _3024_ _3145_ _1537_ vssd1 vssd1 vccd1 vccd1 _1538_ sky130_fd_sc_hd__o21ai_1
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5933_ _2309_ _2432_ vssd1 vssd1 vccd1 vccd1 _0283_ sky130_fd_sc_hd__nor2_1
XFILLER_80_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5864_ _3140_ _0585_ vssd1 vssd1 vccd1 vccd1 _2364_ sky130_fd_sc_hd__nand2_1
X_4815_ _0554_ _0593_ _0673_ _0596_ _1323_ vssd1 vssd1 vccd1 vccd1 _1324_ sky130_fd_sc_hd__o221a_1
XFILLER_21_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5795_ _0796_ _3308_ _2293_ _2294_ _2295_ vssd1 vssd1 vccd1 vccd1 _2296_ sky130_fd_sc_hd__o2111a_1
X_4746_ _1247_ _1251_ _1254_ vssd1 vssd1 vccd1 vccd1 _1255_ sky130_fd_sc_hd__and3_1
X_4677_ _1176_ _1180_ _1183_ _1186_ vssd1 vssd1 vccd1 vccd1 _1187_ sky130_fd_sc_hd__and4_1
X_3628_ _3161_ vssd1 vssd1 vccd1 vccd1 _3162_ sky130_fd_sc_hd__buf_4
X_6416_ _2669_ _2780_ _2783_ _2784_ vssd1 vssd1 vccd1 vccd1 _2785_ sky130_fd_sc_hd__o211a_1
Xoutput28 net28 vssd1 vssd1 vccd1 vccd1 la_data_out_26_24[0] sky130_fd_sc_hd__buf_12
X_6347_ egd_top.BitStream_buffer.BitStream_buffer_output\[6\] egd_top.BitStream_buffer.BitStream_buffer_output\[5\]
+ vssd1 vssd1 vccd1 vccd1 _2718_ sky130_fd_sc_hd__nand2_1
X_3559_ _3092_ vssd1 vssd1 vccd1 vccd1 _3093_ sky130_fd_sc_hd__buf_4
X_6278_ egd_top.BitStream_buffer.BitStream_buffer_output\[6\] vssd1 vssd1 vccd1 vccd1
+ _2649_ sky130_fd_sc_hd__inv_2
X_5229_ _0328_ _0716_ vssd1 vssd1 vccd1 vccd1 _1734_ sky130_fd_sc_hd__nand2_1
XFILLER_56_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4600_ egd_top.BitStream_buffer.BS_buffer\[64\] _0469_ _0751_ _0473_ _1109_ vssd1
+ vssd1 vccd1 vccd1 _1110_ sky130_fd_sc_hd__a221oi_1
XFILLER_30_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5580_ _0405_ _0459_ vssd1 vssd1 vccd1 vccd1 _2082_ sky130_fd_sc_hd__nand2_1
X_4531_ _3264_ _3224_ _3248_ _3226_ _1041_ vssd1 vssd1 vccd1 vccd1 _1042_ sky130_fd_sc_hd__a221oi_1
XFILLER_7_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4462_ _0670_ _0570_ vssd1 vssd1 vccd1 vccd1 _0973_ sky130_fd_sc_hd__or2_1
XFILLER_7_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6201_ _2594_ _2582_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.pc\[3\] sky130_fd_sc_hd__xnor2_4
X_3413_ egd_top.BitStream_buffer.BitStream_buffer_valid_n vssd1 vssd1 vccd1 vccd1
+ _2964_ sky130_fd_sc_hd__inv_2
X_4393_ _0524_ _0530_ _0532_ _0523_ vssd1 vssd1 vccd1 vccd1 _0905_ sky130_fd_sc_hd__o22a_1
X_3344_ _2901_ vssd1 vssd1 vccd1 vccd1 _2902_ sky130_fd_sc_hd__clkbuf_4
X_6132_ _2531_ _1574_ vssd1 vssd1 vccd1 vccd1 _2550_ sky130_fd_sc_hd__nand2_1
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6063_ _2509_ vssd1 vssd1 vccd1 vccd1 _2511_ sky130_fd_sc_hd__buf_2
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5014_ _1505_ _1520_ vssd1 vssd1 vccd1 vccd1 _1521_ sky130_fd_sc_hd__nand2_1
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5916_ _0692_ _0571_ _2413_ _2414_ _2415_ vssd1 vssd1 vccd1 vccd1 _2416_ sky130_fd_sc_hd__o2111a_1
XFILLER_41_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5847_ _3300_ egd_top.BitStream_buffer.BS_buffer\[95\] vssd1 vssd1 vccd1 vccd1 _2347_
+ sky130_fd_sc_hd__nand2_1
X_5778_ _3293_ _3224_ _3315_ _3226_ _2278_ vssd1 vssd1 vccd1 vccd1 _2279_ sky130_fd_sc_hd__a221oi_1
X_4729_ _1226_ _1230_ _1234_ _1237_ vssd1 vssd1 vccd1 vccd1 _1238_ sky130_fd_sc_hd__and4_1
XFILLER_67_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6750_ net154 _0209_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[70\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_23_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3962_ _0475_ vssd1 vssd1 vccd1 vccd1 _0476_ sky130_fd_sc_hd__clkbuf_2
X_5701_ _0461_ _0395_ _0398_ _0459_ _2201_ vssd1 vssd1 vccd1 vccd1 _2202_ sky130_fd_sc_hd__a221oi_2
XFILLER_31_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3893_ egd_top.BitStream_buffer.BS_buffer\[46\] vssd1 vssd1 vccd1 vccd1 _0407_ sky130_fd_sc_hd__clkbuf_4
XFILLER_50_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5632_ _3310_ _0708_ vssd1 vssd1 vccd1 vccd1 _2134_ sky130_fd_sc_hd__nand2_1
X_5563_ _2055_ _2059_ _2061_ _2065_ vssd1 vssd1 vccd1 vccd1 _2066_ sky130_fd_sc_hd__and4_1
X_4514_ egd_top.BitStream_buffer.BS_buffer\[108\] vssd1 vssd1 vccd1 vccd1 _1025_ sky130_fd_sc_hd__clkinv_2
X_5494_ _3162_ egd_top.BitStream_buffer.BS_buffer\[124\] vssd1 vssd1 vccd1 vccd1 _1997_
+ sky130_fd_sc_hd__nand2_1
X_4445_ _0452_ _0447_ vssd1 vssd1 vccd1 vccd1 _0956_ sky130_fd_sc_hd__nand2_1
X_4376_ _0453_ _0459_ vssd1 vssd1 vccd1 vccd1 _0888_ sky130_fd_sc_hd__nand2_1
X_6115_ _2538_ _0755_ vssd1 vssd1 vccd1 vccd1 _2541_ sky130_fd_sc_hd__nand2_1
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6046_ _3005_ _2487_ _2488_ _2500_ vssd1 vssd1 vccd1 vccd1 _0238_ sky130_fd_sc_hd__o211a_1
XFILLER_66_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4230_ _0741_ _3180_ _0623_ _3186_ _0742_ vssd1 vssd1 vccd1 vccd1 _0743_ sky130_fd_sc_hd__a221oi_1
XFILLER_4_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4161_ _0673_ _0571_ vssd1 vssd1 vccd1 vccd1 _0674_ sky130_fd_sc_hd__or2_1
XFILLER_4_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4092_ _0605_ vssd1 vssd1 vccd1 vccd1 _0606_ sky130_fd_sc_hd__buf_2
XFILLER_67_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6802_ net46 _0261_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_23_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4994_ _0509_ _0487_ _0519_ _0490_ _1500_ vssd1 vssd1 vccd1 vccd1 _1501_ sky130_fd_sc_hd__a221oi_1
X_3945_ egd_top.BitStream_buffer.BS_buffer\[58\] vssd1 vssd1 vccd1 vccd1 _0459_ sky130_fd_sc_hd__clkbuf_4
X_6733_ net137 _0192_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[103\]
+ sky130_fd_sc_hd__dfxtp_1
X_5615_ _0496_ _0540_ vssd1 vssd1 vccd1 vccd1 _2117_ sky130_fd_sc_hd__nand2_1
X_3876_ _0388_ _0389_ vssd1 vssd1 vccd1 vccd1 _0390_ sky130_fd_sc_hd__nand2_1
XFILLER_31_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5546_ _0629_ _0546_ _2048_ vssd1 vssd1 vccd1 vccd1 _2049_ sky130_fd_sc_hd__o21ai_1
X_5477_ _3276_ _3216_ _0837_ _3220_ _1979_ vssd1 vssd1 vccd1 vccd1 _1980_ sky130_fd_sc_hd__a221oi_1
X_4428_ _0347_ _0342_ _0345_ _0375_ _0938_ vssd1 vssd1 vccd1 vccd1 _0939_ sky130_fd_sc_hd__a221oi_1
XFILLER_86_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4359_ _0388_ _0393_ vssd1 vssd1 vccd1 vccd1 _0871_ sky130_fd_sc_hd__nand2_1
XFILLER_48_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6029_ _2979_ _2487_ _2488_ _2491_ vssd1 vssd1 vccd1 vccd1 _0246_ sky130_fd_sc_hd__o211a_1
XFILLER_64_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3730_ egd_top.BitStream_buffer.BS_buffer\[73\] vssd1 vssd1 vccd1 vccd1 _3264_ sky130_fd_sc_hd__clkbuf_4
XFILLER_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3661_ _3087_ _3142_ vssd1 vssd1 vccd1 vccd1 _3195_ sky130_fd_sc_hd__and2_1
XFILLER_70_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3592_ _3041_ _3125_ vssd1 vssd1 vccd1 vccd1 _3126_ sky130_fd_sc_hd__nor2_2
XFILLER_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6380_ _2746_ _2749_ _2681_ vssd1 vssd1 vccd1 vccd1 _2750_ sky130_fd_sc_hd__nand3_1
X_5400_ _1144_ _3240_ _1903_ vssd1 vssd1 vccd1 vccd1 _1904_ sky130_fd_sc_hd__o21ai_1
X_5331_ _0407_ _0342_ _0345_ _0642_ _1834_ vssd1 vssd1 vccd1 vccd1 _1835_ sky130_fd_sc_hd__a221oi_1
XFILLER_5_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5262_ _3187_ _3193_ _3196_ _0623_ _1766_ vssd1 vssd1 vccd1 vccd1 _1767_ sky130_fd_sc_hd__a221oi_1
X_5193_ _0510_ _0604_ _1696_ _1697_ _1698_ vssd1 vssd1 vccd1 vccd1 _1699_ sky130_fd_sc_hd__o2111a_1
X_4213_ _3078_ vssd1 vssd1 vccd1 vccd1 _0726_ sky130_fd_sc_hd__clkbuf_4
XFILLER_68_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4144_ _0434_ _0454_ vssd1 vssd1 vccd1 vccd1 _0657_ sky130_fd_sc_hd__nand2_1
XFILLER_55_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6582__123 clknet_1_0__leaf__2889_ vssd1 vssd1 vccd1 vccd1 net157 sky130_fd_sc_hd__inv_2
XFILLER_18_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4075_ _0586_ _0588_ vssd1 vssd1 vccd1 vccd1 _0589_ sky130_fd_sc_hd__or2_1
XFILLER_83_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6716_ net120 _0175_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[81\]
+ sky130_fd_sc_hd__dfxtp_1
X_4977_ _0647_ _0439_ _1483_ vssd1 vssd1 vccd1 vccd1 _1484_ sky130_fd_sc_hd__o21ai_1
X_3928_ _0441_ vssd1 vssd1 vccd1 vccd1 _0442_ sky130_fd_sc_hd__buf_2
X_3859_ _0366_ _0368_ _0372_ vssd1 vssd1 vccd1 vccd1 _0373_ sky130_fd_sc_hd__o21ai_1
XFILLER_50_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5529_ _0458_ _3217_ vssd1 vssd1 vccd1 vccd1 _2032_ sky130_fd_sc_hd__nand2_1
XFILLER_78_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6655__30 clknet_1_1__leaf__2895_ vssd1 vssd1 vccd1 vccd1 net64 sky130_fd_sc_hd__inv_2
XFILLER_75_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f__2884_ clknet_0__2884_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__2884_
+ sky130_fd_sc_hd__clkbuf_16
X_5880_ _0401_ _0368_ _2379_ vssd1 vssd1 vccd1 vccd1 _2380_ sky130_fd_sc_hd__o21ai_1
X_4900_ _3094_ _3339_ _0716_ _0322_ _1407_ vssd1 vssd1 vccd1 vccd1 _1408_ sky130_fd_sc_hd__a221oi_1
X_4831_ _0370_ _0354_ vssd1 vssd1 vccd1 vccd1 _1339_ sky130_fd_sc_hd__nand2_1
XFILLER_21_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4762_ _1258_ _1262_ _1267_ _1270_ vssd1 vssd1 vccd1 vccd1 _1271_ sky130_fd_sc_hd__and4_1
X_4693_ _1174_ _1202_ vssd1 vssd1 vccd1 vccd1 _1203_ sky130_fd_sc_hd__nor2_1
X_6501_ _2926_ _2860_ vssd1 vssd1 vccd1 vccd1 _2863_ sky130_fd_sc_hd__nor2_1
X_3713_ _3230_ _3233_ _3236_ _3237_ _3246_ vssd1 vssd1 vccd1 vccd1 _3247_ sky130_fd_sc_hd__a221oi_1
X_3644_ _3071_ _3142_ vssd1 vssd1 vccd1 vccd1 _3178_ sky130_fd_sc_hd__and2_1
X_6432_ _2798_ _2659_ vssd1 vssd1 vccd1 vccd1 _2799_ sky130_fd_sc_hd__or2_1
X_6363_ _2726_ _2733_ _2681_ vssd1 vssd1 vccd1 vccd1 _2734_ sky130_fd_sc_hd__nand3_1
X_3575_ egd_top.BitStream_buffer.BS_buffer\[106\] vssd1 vssd1 vccd1 vccd1 _3109_ sky130_fd_sc_hd__clkbuf_4
X_5314_ _0574_ _0593_ _0679_ _0596_ _1818_ vssd1 vssd1 vccd1 vccd1 _1819_ sky130_fd_sc_hd__o221a_1
X_6294_ _2664_ vssd1 vssd1 vccd1 vccd1 _2665_ sky130_fd_sc_hd__inv_2
XFILLER_88_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5245_ _3270_ _0774_ vssd1 vssd1 vccd1 vccd1 _1750_ sky130_fd_sc_hd__nand2_1
X_5176_ _0548_ _0337_ vssd1 vssd1 vccd1 vccd1 _1682_ sky130_fd_sc_hd__nand2_1
X_4127_ _0382_ egd_top.BitStream_buffer.BS_buffer\[42\] vssd1 vssd1 vccd1 vccd1 _0640_
+ sky130_fd_sc_hd__nand2_1
X_4058_ _0569_ _0571_ vssd1 vssd1 vccd1 vccd1 _0572_ sky130_fd_sc_hd__or2_1
XFILLER_83_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3360_ _2912_ _2914_ vssd1 vssd1 vccd1 vccd1 _0318_ sky130_fd_sc_hd__nor2_1
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5030_ _3148_ _0623_ vssd1 vssd1 vccd1 vccd1 _1537_ sky130_fd_sc_hd__nand2_1
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6634__11 clknet_1_0__leaf__2893_ vssd1 vssd1 vccd1 vccd1 net45 sky130_fd_sc_hd__inv_2
XFILLER_65_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_224 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5932_ _3026_ _2431_ vssd1 vssd1 vccd1 vccd1 _2432_ sky130_fd_sc_hd__nor2_1
XFILLER_53_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5863_ _3147_ _0553_ vssd1 vssd1 vccd1 vccd1 _2363_ sky130_fd_sc_hd__nand2_1
X_4814_ _0670_ _0599_ vssd1 vssd1 vccd1 vccd1 _1323_ sky130_fd_sc_hd__or2_1
XFILLER_61_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5794_ _3049_ _3319_ vssd1 vssd1 vccd1 vccd1 _2295_ sky130_fd_sc_hd__or2_1
X_4745_ egd_top.BitStream_buffer.BS_buffer\[123\] _3194_ _3197_ _3173_ _1253_ vssd1
+ vssd1 vccd1 vccd1 _1254_ sky130_fd_sc_hd__a221oi_1
XFILLER_31_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4676_ _3153_ _0726_ _3157_ _3081_ _1185_ vssd1 vssd1 vccd1 vccd1 _1186_ sky130_fd_sc_hd__a221oi_1
X_3627_ _3045_ _3142_ vssd1 vssd1 vccd1 vccd1 _3161_ sky130_fd_sc_hd__and2_1
X_6415_ _2665_ egd_top.BitStream_buffer.BitStream_buffer_output\[12\] _2757_ vssd1
+ vssd1 vccd1 vccd1 _2784_ sky130_fd_sc_hd__nand3_1
X_3558_ _3041_ _3091_ vssd1 vssd1 vccd1 vccd1 _3092_ sky130_fd_sc_hd__nor2_2
Xoutput29 net29 vssd1 vssd1 vccd1 vccd1 la_data_out_26_24[1] sky130_fd_sc_hd__buf_12
X_6346_ _2673_ vssd1 vssd1 vccd1 vccd1 _2717_ sky130_fd_sc_hd__inv_2
XFILLER_88_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3489_ egd_top.BitStream_buffer.BS_buffer\[127\] vssd1 vssd1 vccd1 vccd1 _3024_ sky130_fd_sc_hd__clkinv_2
X_6277_ _2647_ _1945_ vssd1 vssd1 vccd1 vccd1 _2648_ sky130_fd_sc_hd__nand2_1
X_5228_ _3049_ _3329_ _1730_ _1731_ _1732_ vssd1 vssd1 vccd1 vccd1 _1733_ sky130_fd_sc_hd__o2111a_1
X_5159_ _0458_ _3230_ vssd1 vssd1 vccd1 vccd1 _1665_ sky130_fd_sc_hd__nand2_1
XFILLER_29_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_390 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_427 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4530_ _3257_ _3218_ _1040_ vssd1 vssd1 vccd1 vccd1 _1041_ sky130_fd_sc_hd__o21ai_1
XFILLER_11_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4461_ _0560_ _0585_ vssd1 vssd1 vccd1 vccd1 _0972_ sky130_fd_sc_hd__nand2_1
XFILLER_7_75 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3412_ net28 _2951_ _2913_ _2963_ vssd1 vssd1 vccd1 vccd1 _0315_ sky130_fd_sc_hd__o211a_1
X_6200_ _2583_ _2584_ vssd1 vssd1 vccd1 vccd1 _2594_ sky130_fd_sc_hd__nand2_2
X_6698__69 clknet_1_1__leaf__2899_ vssd1 vssd1 vccd1 vccd1 net103 sky130_fd_sc_hd__inv_2
X_4392_ _0519_ _0514_ _0527_ _0901_ _0903_ vssd1 vssd1 vccd1 vccd1 _0904_ sky130_fd_sc_hd__a221oi_1
X_6131_ _3017_ _2533_ _2543_ _2549_ vssd1 vssd1 vccd1 vccd1 _0202_ sky130_fd_sc_hd__o211a_1
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3343_ net19 vssd1 vssd1 vccd1 vccd1 _2901_ sky130_fd_sc_hd__clkbuf_4
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6062_ _2509_ vssd1 vssd1 vccd1 vccd1 _2510_ sky130_fd_sc_hd__buf_2
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5013_ _1509_ _1513_ _1515_ _1519_ vssd1 vssd1 vccd1 vccd1 _1520_ sky130_fd_sc_hd__and4_1
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5915_ _0986_ _0557_ vssd1 vssd1 vccd1 vccd1 _2415_ sky130_fd_sc_hd__or2_1
XFILLER_53_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5846_ _3294_ egd_top.BitStream_buffer.BS_buffer\[97\] vssd1 vssd1 vccd1 vccd1 _2346_
+ sky130_fd_sc_hd__nand2_1
X_5777_ _3302_ _3215_ _3219_ _3288_ vssd1 vssd1 vccd1 vccd1 _2278_ sky130_fd_sc_hd__a22o_1
X_4728_ _3157_ _0726_ _3204_ _3081_ _1236_ vssd1 vssd1 vccd1 vccd1 _1237_ sky130_fd_sc_hd__a221oi_2
X_4659_ egd_top.BitStream_buffer.BS_buffer\[97\] vssd1 vssd1 vccd1 vccd1 _1169_ sky130_fd_sc_hd__clkinv_2
X_6329_ _2699_ vssd1 vssd1 vccd1 vccd1 _2700_ sky130_fd_sc_hd__inv_2
XFILLER_88_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3961_ _3076_ _2933_ vssd1 vssd1 vccd1 vccd1 _0475_ sky130_fd_sc_hd__and2_1
XFILLER_50_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5700_ _0647_ _0402_ _2200_ vssd1 vssd1 vccd1 vccd1 _2201_ sky130_fd_sc_hd__o21ai_1
XFILLER_92_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3892_ _0405_ vssd1 vssd1 vccd1 vccd1 _0406_ sky130_fd_sc_hd__buf_2
XFILLER_31_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5631_ _3338_ _3292_ _3341_ _3295_ _2132_ vssd1 vssd1 vccd1 vccd1 _2133_ sky130_fd_sc_hd__a221oi_1
X_5562_ _0532_ _0604_ _2062_ _2063_ _2064_ vssd1 vssd1 vccd1 vccd1 _2065_ sky130_fd_sc_hd__o2111a_1
X_4513_ _0718_ _3106_ _1021_ _1022_ _1023_ vssd1 vssd1 vccd1 vccd1 _1024_ sky130_fd_sc_hd__o2111a_1
X_5493_ _0792_ _3194_ _3197_ _0930_ _1995_ vssd1 vssd1 vccd1 vccd1 _1996_ sky130_fd_sc_hd__a221oi_1
X_4444_ egd_top.BitStream_buffer.BS_buffer\[62\] vssd1 vssd1 vccd1 vccd1 _0955_ sky130_fd_sc_hd__clkinv_2
X_4375_ _0471_ vssd1 vssd1 vccd1 vccd1 _0887_ sky130_fd_sc_hd__inv_2
X_6114_ _2992_ _2532_ _2528_ _2540_ vssd1 vssd1 vccd1 vccd1 _0210_ sky130_fd_sc_hd__o211a_1
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6045_ _2494_ _0861_ vssd1 vssd1 vccd1 vccd1 _2500_ sky130_fd_sc_hd__nand2_1
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5829_ _2986_ _3105_ vssd1 vssd1 vccd1 vccd1 _2329_ sky130_fd_sc_hd__or2_1
XFILLER_78_46 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4160_ egd_top.BitStream_buffer.BS_buffer\[6\] vssd1 vssd1 vccd1 vccd1 _0673_ sky130_fd_sc_hd__inv_2
XFILLER_67_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4091_ _0559_ _3068_ vssd1 vssd1 vccd1 vccd1 _0605_ sky130_fd_sc_hd__nor2_2
XFILLER_67_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6801_ net45 _0260_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_51_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4993_ _0528_ _0495_ _1499_ vssd1 vssd1 vccd1 vccd1 _1500_ sky130_fd_sc_hd__o21ai_1
XFILLER_63_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3944_ _0457_ vssd1 vssd1 vccd1 vccd1 _0458_ sky130_fd_sc_hd__buf_2
XFILLER_23_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6732_ net136 _0191_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[104\]
+ sky130_fd_sc_hd__dfxtp_2
X_3875_ egd_top.BitStream_buffer.BS_buffer\[42\] vssd1 vssd1 vccd1 vccd1 _0389_ sky130_fd_sc_hd__clkbuf_4
X_5614_ _0486_ egd_top.BitStream_buffer.BS_buffer\[28\] vssd1 vssd1 vccd1 vccd1 _2116_
+ sky130_fd_sc_hd__nand2_1
X_5545_ _0548_ _0347_ vssd1 vssd1 vccd1 vccd1 _2048_ sky130_fd_sc_hd__nand2_1
X_5476_ _0842_ _1145_ _1978_ vssd1 vssd1 vccd1 vccd1 _1979_ sky130_fd_sc_hd__o21ai_1
X_4427_ _0936_ _0350_ _0937_ vssd1 vssd1 vccd1 vccd1 _0938_ sky130_fd_sc_hd__o21ai_1
XFILLER_86_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4358_ egd_top.BitStream_buffer.BS_buffer\[45\] vssd1 vssd1 vccd1 vccd1 _0870_ sky130_fd_sc_hd__clkinv_2
X_4289_ _3099_ _3128_ vssd1 vssd1 vccd1 vccd1 _0801_ sky130_fd_sc_hd__nand2_1
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6028_ _2489_ _0366_ vssd1 vssd1 vccd1 vccd1 _2491_ sky130_fd_sc_hd__nand2_1
XFILLER_27_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_48 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3660_ _3193_ vssd1 vssd1 vccd1 vccd1 _3194_ sky130_fd_sc_hd__buf_2
X_3591_ _3124_ vssd1 vssd1 vccd1 vccd1 _3125_ sky130_fd_sc_hd__inv_2
XFILLER_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5330_ _0420_ _0350_ _1833_ vssd1 vssd1 vccd1 vccd1 _1834_ sky130_fd_sc_hd__o21ai_1
X_5261_ _3021_ _3199_ _1765_ vssd1 vssd1 vccd1 vccd1 _1766_ sky130_fd_sc_hd__o21ai_1
XFILLER_5_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4212_ _3118_ _3113_ _3117_ _3066_ _0724_ vssd1 vssd1 vccd1 vccd1 _0725_ sky130_fd_sc_hd__a221oi_1
X_5192_ _0986_ _0613_ vssd1 vssd1 vccd1 vccd1 _1698_ sky130_fd_sc_hd__or2_1
XFILLER_68_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4143_ _0441_ _0655_ vssd1 vssd1 vccd1 vccd1 _0656_ sky130_fd_sc_hd__nand2_1
X_4074_ _0587_ vssd1 vssd1 vccd1 vccd1 _0588_ sky130_fd_sc_hd__buf_2
XFILLER_68_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_311 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6715_ net119 _0174_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[82\]
+ sky130_fd_sc_hd__dfxtp_1
X_4976_ _0442_ _0447_ vssd1 vssd1 vccd1 vccd1 _1483_ sky130_fd_sc_hd__nand2_1
XFILLER_51_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3927_ _0440_ vssd1 vssd1 vccd1 vccd1 _0441_ sky130_fd_sc_hd__clkbuf_2
X_3858_ _0371_ egd_top.BitStream_buffer.BS_buffer\[32\] vssd1 vssd1 vccd1 vccd1 _0372_
+ sky130_fd_sc_hd__nand2_1
X_6646_ clknet_1_0__leaf__2882_ vssd1 vssd1 vccd1 vccd1 _2895_ sky130_fd_sc_hd__buf_1
X_3789_ _3290_ _3111_ vssd1 vssd1 vccd1 vccd1 _3323_ sky130_fd_sc_hd__nor2_2
X_5528_ _0453_ _3237_ vssd1 vssd1 vccd1 vccd1 _2031_ sky130_fd_sc_hd__nand2_1
X_5459_ _1950_ _1954_ _1958_ _1961_ vssd1 vssd1 vccd1 vccd1 _1962_ sky130_fd_sc_hd__and4_1
XFILLER_86_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_171 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__2883_ clknet_0__2883_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__2883_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_92_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4830_ _0389_ _0342_ _0345_ _0869_ _1337_ vssd1 vssd1 vccd1 vccd1 _1338_ sky130_fd_sc_hd__a221oi_1
XFILLER_33_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4761_ _3302_ _3270_ _3288_ _3274_ _1269_ vssd1 vssd1 vccd1 vccd1 _1270_ sky130_fd_sc_hd__a221oi_1
X_4692_ _1187_ _1201_ vssd1 vssd1 vccd1 vccd1 _1202_ sky130_fd_sc_hd__nand2_1
X_6500_ _2852_ _2861_ vssd1 vssd1 vccd1 vccd1 _2862_ sky130_fd_sc_hd__nand2_1
X_3712_ _3238_ _3240_ _3245_ vssd1 vssd1 vccd1 vccd1 _3246_ sky130_fd_sc_hd__o21ai_1
X_3643_ egd_top.BitStream_buffer.BS_buffer\[125\] vssd1 vssd1 vccd1 vccd1 _3177_ sky130_fd_sc_hd__clkbuf_4
X_6431_ _2700_ _2684_ vssd1 vssd1 vccd1 vccd1 _2798_ sky130_fd_sc_hd__nand2_1
X_6362_ _2729_ _2732_ vssd1 vssd1 vccd1 vccd1 _2733_ sky130_fd_sc_hd__nand2_1
X_5313_ _0676_ _0599_ vssd1 vssd1 vccd1 vccd1 _1818_ sky130_fd_sc_hd__or2_1
X_3574_ _3085_ _3089_ _3095_ _3101_ _3107_ vssd1 vssd1 vccd1 vccd1 _3108_ sky130_fd_sc_hd__o2111a_1
X_6293_ _2663_ _2644_ vssd1 vssd1 vccd1 vccd1 _2664_ sky130_fd_sc_hd__nand2_1
X_5244_ _3296_ _1145_ _1746_ _1747_ _1748_ vssd1 vssd1 vccd1 vccd1 _1749_ sky130_fd_sc_hd__o2111a_1
X_5175_ _0995_ _0523_ _0865_ _0526_ _1680_ vssd1 vssd1 vccd1 vccd1 _1681_ sky130_fd_sc_hd__o221a_1
XFILLER_68_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4126_ _0387_ egd_top.BitStream_buffer.BS_buffer\[43\] vssd1 vssd1 vccd1 vccd1 _0639_
+ sky130_fd_sc_hd__nand2_1
XFILLER_83_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4057_ _0570_ vssd1 vssd1 vccd1 vccd1 _0571_ sky130_fd_sc_hd__clkbuf_2
XFILLER_51_130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4959_ egd_top.BitStream_buffer.BS_buffer\[46\] vssd1 vssd1 vccd1 vccd1 _1466_ sky130_fd_sc_hd__inv_2
XFILLER_3_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_494 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6549__93 clknet_1_1__leaf__2886_ vssd1 vssd1 vccd1 vccd1 net127 sky130_fd_sc_hd__inv_2
XFILLER_51_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5931_ _2372_ _2429_ _2430_ vssd1 vssd1 vccd1 vccd1 _2431_ sky130_fd_sc_hd__nand3_1
XFILLER_53_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5862_ _2358_ _2359_ _2360_ _2361_ vssd1 vssd1 vccd1 vccd1 _2362_ sky130_fd_sc_hd__and4_1
XFILLER_33_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4813_ _0688_ _0588_ _1319_ _1320_ _1321_ vssd1 vssd1 vccd1 vccd1 _1322_ sky130_fd_sc_hd__o2111a_1
X_5793_ _3310_ _3062_ vssd1 vssd1 vccd1 vccd1 _2294_ sky130_fd_sc_hd__nand2_1
X_4744_ _3009_ _3200_ _1252_ vssd1 vssd1 vccd1 vccd1 _1253_ sky130_fd_sc_hd__o21ai_1
X_4675_ _2977_ _0729_ _1184_ vssd1 vssd1 vccd1 vccd1 _1185_ sky130_fd_sc_hd__o21ai_1
X_3626_ _3159_ vssd1 vssd1 vccd1 vccd1 _3160_ sky130_fd_sc_hd__buf_4
X_6414_ _2781_ _2782_ _2717_ vssd1 vssd1 vccd1 vccd1 _2783_ sky130_fd_sc_hd__o21ai_1
X_3557_ _3090_ vssd1 vssd1 vccd1 vccd1 _3091_ sky130_fd_sc_hd__inv_2
X_6345_ _2665_ _2715_ vssd1 vssd1 vccd1 vccd1 _2716_ sky130_fd_sc_hd__nand2_1
X_6276_ _2646_ _2629_ vssd1 vssd1 vccd1 vccd1 _2647_ sky130_fd_sc_hd__nand2_1
X_5227_ _3325_ _3094_ vssd1 vssd1 vccd1 vccd1 _1732_ sky130_fd_sc_hd__nand2_1
X_3488_ net1 vssd1 vssd1 vccd1 vccd1 _3023_ sky130_fd_sc_hd__clkbuf_4
XFILLER_84_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5158_ _0478_ _0432_ _0435_ _0664_ _1663_ vssd1 vssd1 vccd1 vccd1 _1664_ sky130_fd_sc_hd__a221oi_1
XFILLER_29_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4109_ egd_top.BitStream_buffer.BS_buffer\[0\] vssd1 vssd1 vccd1 vccd1 _0623_ sky130_fd_sc_hd__buf_2
X_5089_ _3127_ _3169_ vssd1 vssd1 vccd1 vccd1 _1595_ sky130_fd_sc_hd__nand2_1
XFILLER_56_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4460_ _0564_ _0553_ vssd1 vssd1 vccd1 vccd1 _0971_ sky130_fd_sc_hd__nand2_1
XFILLER_7_87 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4391_ _0510_ _0506_ _0902_ vssd1 vssd1 vccd1 vccd1 _0903_ sky130_fd_sc_hd__o21ai_1
X_3411_ _2951_ _2962_ vssd1 vssd1 vccd1 vccd1 _2963_ sky130_fd_sc_hd__nand2_1
X_6130_ _2538_ _1426_ vssd1 vssd1 vccd1 vccd1 _2549_ sky130_fd_sc_hd__nand2_1
X_3342_ net33 net32 net31 vssd1 vssd1 vccd1 vccd1 _2900_ sky130_fd_sc_hd__and3_1
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6061_ _2508_ vssd1 vssd1 vccd1 vccd1 _2509_ sky130_fd_sc_hd__inv_2
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5012_ _1128_ _0604_ _1516_ _1517_ _1518_ vssd1 vssd1 vccd1 vccd1 _1519_ sky130_fd_sc_hd__o2111a_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5914_ _0565_ _0491_ vssd1 vssd1 vccd1 vccd1 _2414_ sky130_fd_sc_hd__nand2_1
X_5845_ _3102_ _3307_ _2342_ _2343_ _2344_ vssd1 vssd1 vccd1 vccd1 _2345_ sky130_fd_sc_hd__o2111a_1
XFILLER_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5776_ _2262_ _2276_ vssd1 vssd1 vccd1 vccd1 _2277_ sky130_fd_sc_hd__nand2_1
XFILLER_21_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4727_ _2980_ _0729_ _1235_ vssd1 vssd1 vccd1 vccd1 _1236_ sky130_fd_sc_hd__o21ai_1
X_6528__74 clknet_1_0__leaf__2884_ vssd1 vssd1 vccd1 vccd1 net108 sky130_fd_sc_hd__inv_2
X_4658_ _3338_ _3324_ _3326_ _3341_ _1167_ vssd1 vssd1 vccd1 vccd1 _1168_ sky130_fd_sc_hd__a221oi_1
X_3609_ _3124_ _3142_ vssd1 vssd1 vccd1 vccd1 _3143_ sky130_fd_sc_hd__and2_1
X_6543__88 clknet_1_0__leaf__2885_ vssd1 vssd1 vccd1 vccd1 net122 sky130_fd_sc_hd__inv_2
XFILLER_1_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4589_ _0887_ _0463_ vssd1 vssd1 vccd1 vccd1 _1099_ sky130_fd_sc_hd__or2_1
XFILLER_88_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6328_ _2696_ _2698_ vssd1 vssd1 vccd1 vccd1 _2699_ sky130_fd_sc_hd__and2_1
X_6259_ _2628_ _1945_ _2629_ egd_top.BitStream_buffer.BitStream_buffer_output\[7\]
+ egd_top.BitStream_buffer.BitStream_buffer_output\[6\] vssd1 vssd1 vccd1 vccd1 _2630_
+ sky130_fd_sc_hd__a311oi_2
XFILLER_49_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3960_ egd_top.BitStream_buffer.BS_buffer\[63\] vssd1 vssd1 vccd1 vccd1 _0474_ sky130_fd_sc_hd__clkinv_2
XFILLER_16_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3891_ _0404_ vssd1 vssd1 vccd1 vccd1 _0405_ sky130_fd_sc_hd__inv_2
XFILLER_85_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5630_ _1003_ _3299_ _2131_ vssd1 vssd1 vccd1 vccd1 _2132_ sky130_fd_sc_hd__o21ai_1
X_5561_ _0520_ _0613_ vssd1 vssd1 vccd1 vccd1 _2064_ sky130_fd_sc_hd__or2_1
XFILLER_31_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5492_ _1602_ _3200_ _1994_ vssd1 vssd1 vccd1 vccd1 _1995_ sky130_fd_sc_hd__o21ai_1
X_4512_ _0721_ _3088_ vssd1 vssd1 vccd1 vccd1 _1023_ sky130_fd_sc_hd__or2_1
XFILLER_7_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4443_ _0664_ _0470_ _3244_ _0473_ _0953_ vssd1 vssd1 vccd1 vccd1 _0954_ sky130_fd_sc_hd__a221oi_1
X_4374_ _0454_ _0432_ _0435_ _0461_ _0885_ vssd1 vssd1 vccd1 vccd1 _0886_ sky130_fd_sc_hd__a221oi_1
X_6113_ _2538_ _1360_ vssd1 vssd1 vccd1 vccd1 _2540_ sky130_fd_sc_hd__nand2_1
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6044_ _3001_ _2487_ _2488_ _2499_ vssd1 vssd1 vccd1 vccd1 _0239_ sky130_fd_sc_hd__o211a_1
XFILLER_85_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5828_ _3099_ egd_top.BitStream_buffer.BS_buffer\[116\] vssd1 vssd1 vccd1 vccd1 _2328_
+ sky130_fd_sc_hd__nand2_1
XFILLER_22_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5759_ _3006_ _0729_ _2259_ vssd1 vssd1 vccd1 vccd1 _2260_ sky130_fd_sc_hd__o21ai_1
XFILLER_1_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_504 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_386 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4090_ _0603_ vssd1 vssd1 vccd1 vccd1 _0604_ sky130_fd_sc_hd__buf_2
XFILLER_67_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6800_ net44 _0259_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_4992_ _0497_ _0531_ vssd1 vssd1 vccd1 vccd1 _1499_ sky130_fd_sc_hd__nand2_1
XFILLER_90_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6731_ net135 _0190_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[105\]
+ sky130_fd_sc_hd__dfxtp_1
X_3943_ _0456_ vssd1 vssd1 vccd1 vccd1 _0457_ sky130_fd_sc_hd__clkinv_2
XFILLER_51_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3874_ _0387_ vssd1 vssd1 vccd1 vccd1 _0388_ sky130_fd_sc_hd__buf_2
X_5613_ _2104_ _2108_ _2110_ _2114_ vssd1 vssd1 vccd1 vccd1 _2115_ sky130_fd_sc_hd__and4_1
X_5544_ _0865_ _0523_ _1276_ _0526_ _2046_ vssd1 vssd1 vccd1 vccd1 _2047_ sky130_fd_sc_hd__o221a_1
XFILLER_8_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5475_ _3223_ _3302_ vssd1 vssd1 vccd1 vccd1 _1978_ sky130_fd_sc_hd__nand2_1
X_4426_ _0353_ _0379_ vssd1 vssd1 vccd1 vccd1 _0937_ sky130_fd_sc_hd__nand2_1
X_4357_ egd_top.BitStream_buffer.BS_buffer\[43\] vssd1 vssd1 vccd1 vccd1 _0869_ sky130_fd_sc_hd__clkbuf_4
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4288_ _3093_ _3100_ vssd1 vssd1 vccd1 vccd1 _0800_ sky130_fd_sc_hd__nand2_1
XFILLER_58_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6682__54 clknet_1_1__leaf__2898_ vssd1 vssd1 vccd1 vccd1 net88 sky130_fd_sc_hd__inv_2
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6027_ _2966_ _2487_ _2488_ _2490_ vssd1 vssd1 vccd1 vccd1 _0247_ sky130_fd_sc_hd__o211a_1
XFILLER_46_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3590_ _3030_ _3031_ egd_top.BitStream_buffer.pc\[3\] vssd1 vssd1 vccd1 vccd1 _3124_
+ sky130_fd_sc_hd__and3_2
X_5260_ _3202_ _3177_ vssd1 vssd1 vccd1 vccd1 _1765_ sky130_fd_sc_hd__nand2_1
X_4211_ _0721_ _3123_ _0723_ vssd1 vssd1 vccd1 vccd1 _0724_ sky130_fd_sc_hd__o21ai_1
XFILLER_48_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5191_ _0609_ _0515_ vssd1 vssd1 vccd1 vccd1 _1697_ sky130_fd_sc_hd__nand2_1
X_4142_ egd_top.BitStream_buffer.BS_buffer\[53\] vssd1 vssd1 vccd1 vccd1 _0655_ sky130_fd_sc_hd__clkbuf_4
X_4073_ _3121_ _0556_ vssd1 vssd1 vccd1 vccd1 _0587_ sky130_fd_sc_hd__nand2_1
XFILLER_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4975_ _0461_ _0415_ _0459_ _0419_ _1481_ vssd1 vssd1 vccd1 vccd1 _1482_ sky130_fd_sc_hd__a221oi_1
XFILLER_51_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6714_ net118 _0173_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[83\]
+ sky130_fd_sc_hd__dfxtp_1
X_3926_ _3090_ _2933_ vssd1 vssd1 vccd1 vccd1 _0440_ sky130_fd_sc_hd__and2_1
XFILLER_51_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3857_ _0370_ vssd1 vssd1 vccd1 vccd1 _0371_ sky130_fd_sc_hd__buf_2
XFILLER_50_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3788_ egd_top.BitStream_buffer.BS_buffer\[90\] vssd1 vssd1 vccd1 vccd1 _3322_ sky130_fd_sc_hd__clkbuf_4
X_5527_ _0751_ _0432_ _0435_ _3230_ _2029_ vssd1 vssd1 vccd1 vccd1 _2030_ sky130_fd_sc_hd__a221oi_1
XFILLER_3_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5458_ _0722_ _3339_ _3109_ _0322_ _1960_ vssd1 vssd1 vccd1 vccd1 _1961_ sky130_fd_sc_hd__a221oi_1
X_4409_ _0682_ _0593_ _0569_ _0599_ _0920_ vssd1 vssd1 vccd1 vccd1 _0921_ sky130_fd_sc_hd__o221a_1
XFILLER_59_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5389_ _3310_ _3028_ vssd1 vssd1 vccd1 vccd1 _1893_ sky130_fd_sc_hd__nand2_1
XFILLER_86_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6566__109 clknet_1_0__leaf__2887_ vssd1 vssd1 vccd1 vccd1 net143 sky130_fd_sc_hd__inv_2
XFILLER_77_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6661__35 clknet_1_1__leaf__2896_ vssd1 vssd1 vccd1 vccd1 net69 sky130_fd_sc_hd__inv_2
XFILLER_37_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__2882_ clknet_0__2882_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__2882_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_73_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4760_ _1158_ _3279_ _1268_ vssd1 vssd1 vccd1 vccd1 _1269_ sky130_fd_sc_hd__o21ai_1
X_4691_ _1190_ _1194_ _1197_ _1200_ vssd1 vssd1 vccd1 vccd1 _1201_ sky130_fd_sc_hd__and4_1
X_3711_ _3243_ _3244_ vssd1 vssd1 vccd1 vccd1 _3245_ sky130_fd_sc_hd__nand2_1
X_3642_ _3175_ vssd1 vssd1 vccd1 vccd1 _3176_ sky130_fd_sc_hd__buf_2
X_6430_ _2797_ vssd1 vssd1 vccd1 vccd1 egd_top.exp_golomb_decoding.te_range\[2\] sky130_fd_sc_hd__inv_2
X_6361_ _2730_ _2731_ vssd1 vssd1 vccd1 vccd1 _2732_ sky130_fd_sc_hd__nand2_1
X_5312_ _0897_ _0576_ _1814_ _1815_ _1816_ vssd1 vssd1 vccd1 vccd1 _1817_ sky130_fd_sc_hd__o2111a_1
X_3573_ _3102_ _3106_ vssd1 vssd1 vccd1 vccd1 _3107_ sky130_fd_sc_hd__or2_1
X_6292_ _2657_ _2624_ _2662_ vssd1 vssd1 vccd1 vccd1 _2663_ sky130_fd_sc_hd__a21oi_4
X_5243_ _3219_ _3283_ vssd1 vssd1 vccd1 vccd1 _1748_ sky130_fd_sc_hd__nand2_1
X_5174_ _0366_ _0530_ _0633_ _0534_ vssd1 vssd1 vccd1 vccd1 _1680_ sky130_fd_sc_hd__o22a_1
XFILLER_68_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4125_ _0377_ egd_top.BitStream_buffer.BS_buffer\[41\] vssd1 vssd1 vccd1 vccd1 _0638_
+ sky130_fd_sc_hd__nand2_1
X_4056_ _3104_ _0556_ vssd1 vssd1 vccd1 vccd1 _0570_ sky130_fd_sc_hd__nand2_1
XFILLER_71_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_142 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4958_ _1335_ _1465_ vssd1 vssd1 vccd1 vccd1 _0291_ sky130_fd_sc_hd__nor2_1
XFILLER_51_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4889_ _3028_ _3323_ _3325_ _3040_ _1396_ vssd1 vssd1 vccd1 vccd1 _1397_ sky130_fd_sc_hd__a221oi_1
X_3909_ egd_top.BitStream_buffer.BS_buffer\[48\] vssd1 vssd1 vccd1 vccd1 _0423_ sky130_fd_sc_hd__clkinv_2
XFILLER_3_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5930_ _0621_ egd_top.BitStream_buffer.BS_buffer\[14\] vssd1 vssd1 vccd1 vccd1 _2430_
+ sky130_fd_sc_hd__nand2_1
XFILLER_53_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5861_ _3155_ egd_top.BitStream_buffer.BS_buffer\[0\] vssd1 vssd1 vccd1 vccd1 _2361_
+ sky130_fd_sc_hd__nand2_1
X_6620__158 clknet_1_0__leaf__2892_ vssd1 vssd1 vccd1 vccd1 net192 sky130_fd_sc_hd__inv_2
X_4812_ _0685_ _0575_ vssd1 vssd1 vccd1 vccd1 _1321_ sky130_fd_sc_hd__or2_1
XFILLER_61_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5792_ _3314_ _3040_ vssd1 vssd1 vccd1 vccd1 _2293_ sky130_fd_sc_hd__nand2_1
X_4743_ _3203_ _3149_ vssd1 vssd1 vccd1 vccd1 _1252_ sky130_fd_sc_hd__nand2_1
X_4674_ _3074_ _3164_ vssd1 vssd1 vccd1 vccd1 _1184_ sky130_fd_sc_hd__nand2_1
X_6413_ _1586_ _2688_ vssd1 vssd1 vccd1 vccd1 _2782_ sky130_fd_sc_hd__nor2_1
X_3625_ _3158_ vssd1 vssd1 vccd1 vccd1 _3159_ sky130_fd_sc_hd__buf_2
X_3556_ _3030_ egd_top.BitStream_buffer.pc\[2\] _3032_ vssd1 vssd1 vccd1 vccd1 _3090_
+ sky130_fd_sc_hd__and3_2
X_6344_ _2713_ _2714_ vssd1 vssd1 vccd1 vccd1 _2715_ sky130_fd_sc_hd__nand2_1
X_6275_ _2645_ _2626_ vssd1 vssd1 vccd1 vccd1 _2646_ sky130_fd_sc_hd__nand2_1
XFILLER_88_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5226_ _3323_ _3062_ vssd1 vssd1 vccd1 vccd1 _1731_ sky130_fd_sc_hd__nand2_1
X_3487_ _3020_ _2976_ _3002_ _3022_ vssd1 vssd1 vccd1 vccd1 _0299_ sky130_fd_sc_hd__o211a_1
XFILLER_56_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5157_ _0887_ _0439_ _1662_ vssd1 vssd1 vccd1 vccd1 _1663_ sky130_fd_sc_hd__o21ai_1
X_5088_ _1035_ _3089_ _1591_ _1592_ _1593_ vssd1 vssd1 vccd1 vccd1 _1594_ sky130_fd_sc_hd__o2111a_1
X_4108_ _0621_ vssd1 vssd1 vccd1 vccd1 _0622_ sky130_fd_sc_hd__clkbuf_4
XFILLER_56_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6640__16 clknet_1_0__leaf__2894_ vssd1 vssd1 vccd1 vccd1 net50 sky130_fd_sc_hd__inv_2
XFILLER_44_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4039_ egd_top.BitStream_buffer.BS_buffer\[7\] vssd1 vssd1 vccd1 vccd1 _0553_ sky130_fd_sc_hd__clkbuf_4
XFILLER_71_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6595__135 clknet_1_0__leaf__2890_ vssd1 vssd1 vccd1 vccd1 net169 sky130_fd_sc_hd__inv_2
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4390_ _0504_ _0515_ vssd1 vssd1 vccd1 vccd1 _0902_ sky130_fd_sc_hd__nand2_1
XFILLER_7_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3410_ net28 _2961_ _2947_ vssd1 vssd1 vccd1 vccd1 _2962_ sky130_fd_sc_hd__o21ba_1
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6060_ net198 _2972_ vssd1 vssd1 vccd1 vccd1 _2508_ sky130_fd_sc_hd__nor2_1
XFILLER_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5011_ _0897_ _0613_ vssd1 vssd1 vccd1 vccd1 _1518_ sky130_fd_sc_hd__or2_1
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5913_ _0561_ _0502_ vssd1 vssd1 vccd1 vccd1 _2413_ sky130_fd_sc_hd__nand2_1
X_5844_ _0709_ _3318_ vssd1 vssd1 vccd1 vccd1 _2344_ sky130_fd_sc_hd__or2_1
XFILLER_34_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5775_ _2265_ _2269_ _2272_ _2275_ vssd1 vssd1 vccd1 vccd1 _2276_ sky130_fd_sc_hd__and4_1
X_4726_ _3073_ egd_top.BitStream_buffer.BS_buffer\[114\] vssd1 vssd1 vccd1 vccd1 _1235_
+ sky130_fd_sc_hd__nand2_1
X_4657_ _0324_ _3330_ _1166_ vssd1 vssd1 vccd1 vccd1 _1167_ sky130_fd_sc_hd__o21ai_1
X_3608_ _3134_ vssd1 vssd1 vccd1 vccd1 _3142_ sky130_fd_sc_hd__buf_2
X_6327_ _2697_ vssd1 vssd1 vccd1 vccd1 _2698_ sky130_fd_sc_hd__inv_2
XFILLER_1_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4588_ _0452_ _0467_ vssd1 vssd1 vccd1 vccd1 _1098_ sky130_fd_sc_hd__nand2_1
X_3539_ _3041_ _3072_ vssd1 vssd1 vccd1 vccd1 _3073_ sky130_fd_sc_hd__nor2_2
XFILLER_1_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6258_ egd_top.BitStream_buffer.BitStream_buffer_output\[4\] vssd1 vssd1 vccd1 vccd1
+ _2629_ sky130_fd_sc_hd__clkinv_2
XFILLER_88_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5209_ _3060_ _3066_ vssd1 vssd1 vccd1 vccd1 _1714_ sky130_fd_sc_hd__nand2_1
X_6189_ _2902_ egd_top.BitStream_buffer.pc\[6\] vssd1 vssd1 vccd1 vccd1 _2588_ sky130_fd_sc_hd__nand2_1
XFILLER_84_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6603__142 clknet_1_0__leaf__2891_ vssd1 vssd1 vccd1 vccd1 net176 sky130_fd_sc_hd__inv_2
XFILLER_16_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6688__60 clknet_1_0__leaf__2898_ vssd1 vssd1 vccd1 vccd1 net94 sky130_fd_sc_hd__inv_2
XFILLER_4_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3890_ _3076_ _0339_ vssd1 vssd1 vccd1 vccd1 _0404_ sky130_fd_sc_hd__nand2_1
XFILLER_43_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5560_ _0609_ _0527_ vssd1 vssd1 vccd1 vccd1 _2063_ sky130_fd_sc_hd__nand2_1
XFILLER_78_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5491_ _3203_ _3187_ vssd1 vssd1 vccd1 vccd1 _1994_ sky130_fd_sc_hd__nand2_1
X_4511_ _3093_ _0714_ vssd1 vssd1 vccd1 vccd1 _1022_ sky130_fd_sc_hd__nand2_1
X_4442_ _0751_ _0476_ _2936_ _3230_ vssd1 vssd1 vccd1 vccd1 _0953_ sky130_fd_sc_hd__a22o_1
X_4373_ _0883_ _0439_ _0884_ vssd1 vssd1 vccd1 vccd1 _0885_ sky130_fd_sc_hd__o21ai_1
X_6112_ _2988_ _2532_ _2528_ _2539_ vssd1 vssd1 vccd1 vccd1 _0211_ sky130_fd_sc_hd__o211a_1
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6043_ _2494_ _0629_ vssd1 vssd1 vccd1 vccd1 _2499_ sky130_fd_sc_hd__nand2_1
XFILLER_85_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5827_ _3092_ _3153_ vssd1 vssd1 vccd1 vccd1 _2327_ sky130_fd_sc_hd__nand2_1
X_5758_ _3074_ _3133_ vssd1 vssd1 vccd1 vccd1 _2259_ sky130_fd_sc_hd__nand2_1
XFILLER_22_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4709_ _1003_ _3308_ _1215_ _1216_ _1217_ vssd1 vssd1 vccd1 vccd1 _1218_ sky130_fd_sc_hd__o2111a_1
X_5689_ egd_top.BitStream_buffer.BitStream_buffer_output\[2\] _2965_ _0627_ vssd1
+ vssd1 vccd1 vccd1 _2190_ sky130_fd_sc_hd__o21ai_1
XFILLER_78_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1__f__2899_ clknet_0__2899_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__2899_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_48_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4991_ _0907_ _0523_ _0633_ _0526_ _1497_ vssd1 vssd1 vccd1 vccd1 _1498_ sky130_fd_sc_hd__o221a_1
XFILLER_63_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6730_ net134 _0189_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[106\]
+ sky130_fd_sc_hd__dfxtp_1
X_3942_ _3110_ _2934_ vssd1 vssd1 vccd1 vccd1 _0456_ sky130_fd_sc_hd__nand2_1
X_3873_ _0386_ vssd1 vssd1 vccd1 vccd1 _0387_ sky130_fd_sc_hd__clkbuf_2
X_5612_ _0524_ _0603_ _2111_ _2112_ _2113_ vssd1 vssd1 vccd1 vccd1 _2114_ sky130_fd_sc_hd__o2111a_1
X_5543_ _0940_ _0530_ _1084_ _0534_ vssd1 vssd1 vccd1 vccd1 _2046_ sky130_fd_sc_hd__o22a_1
X_5474_ _1965_ _1969_ _1973_ _1976_ vssd1 vssd1 vccd1 vccd1 _1977_ sky130_fd_sc_hd__and4_1
X_4425_ egd_top.BitStream_buffer.BS_buffer\[42\] vssd1 vssd1 vccd1 vccd1 _0936_ sky130_fd_sc_hd__inv_2
X_4356_ _0337_ _0360_ _0363_ _0346_ _0867_ vssd1 vssd1 vccd1 vccd1 _0868_ sky130_fd_sc_hd__a221oi_1
X_6667__41 clknet_1_0__leaf__2896_ vssd1 vssd1 vccd1 vccd1 net75 sky130_fd_sc_hd__inv_2
XFILLER_86_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4287_ _0708_ _3039_ _3062_ _3048_ _0798_ vssd1 vssd1 vccd1 vccd1 _0799_ sky130_fd_sc_hd__a221oi_2
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6026_ _2489_ _0995_ vssd1 vssd1 vccd1 vccd1 _2490_ sky130_fd_sc_hd__nand2_1
XFILLER_73_129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6859_ net103 _0318_ vssd1 vssd1 vccd1 vccd1 net31 sky130_fd_sc_hd__dfxtp_1
XFILLER_13_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4210_ _3127_ _0722_ vssd1 vssd1 vccd1 vccd1 _0723_ sky130_fd_sc_hd__nand2_1
X_5190_ _0606_ _0502_ vssd1 vssd1 vccd1 vccd1 _1696_ sky130_fd_sc_hd__nand2_1
X_4141_ _0431_ _0436_ vssd1 vssd1 vccd1 vccd1 _0654_ sky130_fd_sc_hd__nand2_1
X_4072_ _0585_ vssd1 vssd1 vccd1 vccd1 _0586_ sky130_fd_sc_hd__inv_2
XFILLER_83_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_140 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4974_ _0965_ _0422_ _1480_ vssd1 vssd1 vccd1 vccd1 _1481_ sky130_fd_sc_hd__o21ai_1
XFILLER_51_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6713_ net117 _0172_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[84\]
+ sky130_fd_sc_hd__dfxtp_1
X_3925_ _0438_ vssd1 vssd1 vccd1 vccd1 _0439_ sky130_fd_sc_hd__buf_2
X_3856_ _0369_ vssd1 vssd1 vccd1 vccd1 _0370_ sky130_fd_sc_hd__clkbuf_2
X_3787_ _3306_ _3308_ _3312_ _3316_ _3320_ vssd1 vssd1 vccd1 vccd1 _3321_ sky130_fd_sc_hd__o2111a_1
X_5526_ _0663_ _0439_ _2028_ vssd1 vssd1 vccd1 vccd1 _2029_ sky130_fd_sc_hd__o21ai_1
X_5457_ _0718_ _0326_ _1959_ vssd1 vssd1 vccd1 vccd1 _1960_ sky130_fd_sc_hd__o21ai_1
X_4408_ _0597_ _0595_ vssd1 vssd1 vccd1 vccd1 _0920_ sky130_fd_sc_hd__or2_1
XFILLER_59_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5388_ _3314_ _3338_ vssd1 vssd1 vccd1 vccd1 _1892_ sky130_fd_sc_hd__nand2_1
XFILLER_86_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_424 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4339_ _3333_ _3322_ vssd1 vssd1 vccd1 vccd1 _0851_ sky130_fd_sc_hd__nand2_1
X_6009_ _2471_ _0532_ vssd1 vssd1 vccd1 vccd1 _2479_ sky130_fd_sc_hd__nand2_1
XFILLER_91_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_471 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_398 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3710_ egd_top.BitStream_buffer.BS_buffer\[64\] vssd1 vssd1 vccd1 vccd1 _3244_ sky130_fd_sc_hd__clkbuf_4
X_4690_ _0623_ _3176_ _0792_ _3180_ _1199_ vssd1 vssd1 vccd1 vccd1 _1200_ sky130_fd_sc_hd__a221oi_1
X_3641_ _3174_ vssd1 vssd1 vccd1 vccd1 _3175_ sky130_fd_sc_hd__clkbuf_2
XFILLER_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3572_ _3105_ vssd1 vssd1 vccd1 vccd1 _3106_ sky130_fd_sc_hd__buf_2
X_6360_ _2678_ _2629_ vssd1 vssd1 vccd1 vccd1 _2731_ sky130_fd_sc_hd__nand2_1
X_5311_ _0492_ _0588_ vssd1 vssd1 vccd1 vccd1 _1816_ sky130_fd_sc_hd__or2_1
X_6291_ _2623_ vssd1 vssd1 vccd1 vccd1 _2662_ sky130_fd_sc_hd__inv_2
X_5242_ _3223_ _3276_ vssd1 vssd1 vccd1 vccd1 _1747_ sky130_fd_sc_hd__nand2_1
X_5173_ egd_top.BitStream_buffer.BS_buffer\[28\] _0504_ egd_top.BitStream_buffer.BS_buffer\[29\]
+ _0508_ _1678_ vssd1 vssd1 vccd1 vccd1 _1679_ sky130_fd_sc_hd__a221oi_1
X_4124_ egd_top.BitStream_buffer.BS_buffer\[44\] vssd1 vssd1 vccd1 vccd1 _0637_ sky130_fd_sc_hd__clkinv_2
Xinput1 la_data_in_58_43[0] vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__clkbuf_1
X_4055_ _0568_ vssd1 vssd1 vccd1 vccd1 _0569_ sky130_fd_sc_hd__inv_2
XFILLER_91_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4957_ _3026_ _1464_ vssd1 vssd1 vccd1 vccd1 _1465_ sky130_fd_sc_hd__nor2_1
XFILLER_20_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3908_ _0421_ vssd1 vssd1 vccd1 vccd1 _0422_ sky130_fd_sc_hd__buf_2
X_4888_ _0854_ _3329_ _1395_ vssd1 vssd1 vccd1 vccd1 _1396_ sky130_fd_sc_hd__o21ai_1
X_3839_ _0352_ vssd1 vssd1 vccd1 vccd1 _0353_ sky130_fd_sc_hd__buf_2
X_6558_ clknet_1_0__leaf__2883_ vssd1 vssd1 vccd1 vccd1 _2887_ sky130_fd_sc_hd__buf_1
XFILLER_3_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6489_ _2820_ _2832_ _2851_ vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__o21ai_1
X_5509_ _0353_ _0948_ vssd1 vssd1 vccd1 vccd1 _2012_ sky130_fd_sc_hd__nand2_1
XFILLER_10_66 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_452 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6572__114 clknet_1_1__leaf__2888_ vssd1 vssd1 vccd1 vccd1 net148 sky130_fd_sc_hd__inv_2
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5860_ _3167_ egd_top.BitStream_buffer.BS_buffer\[126\] vssd1 vssd1 vccd1 vccd1 _2360_
+ sky130_fd_sc_hd__nand2_1
X_4811_ _0578_ egd_top.BitStream_buffer.BS_buffer\[13\] vssd1 vssd1 vccd1 vccd1 _1320_
+ sky130_fd_sc_hd__nand2_1
XFILLER_61_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5791_ _3028_ _3295_ _3341_ _3292_ _2291_ vssd1 vssd1 vccd1 vccd1 _2292_ sky130_fd_sc_hd__a221oi_1
X_4742_ _3198_ _3156_ _0744_ _3160_ _1250_ vssd1 vssd1 vccd1 vccd1 _1251_ sky130_fd_sc_hd__a221oi_1
XFILLER_33_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4673_ _3075_ _3113_ _3117_ _3082_ _1182_ vssd1 vssd1 vccd1 vccd1 _1183_ sky130_fd_sc_hd__a221oi_1
X_3624_ _3058_ _3142_ vssd1 vssd1 vccd1 vccd1 _3158_ sky130_fd_sc_hd__and2_1
X_6412_ _2687_ _2703_ vssd1 vssd1 vccd1 vccd1 _2781_ sky130_fd_sc_hd__nor2_1
X_3555_ _3088_ vssd1 vssd1 vccd1 vccd1 _3089_ sky130_fd_sc_hd__clkbuf_4
X_6343_ egd_top.BitStream_buffer.BitStream_buffer_output\[10\] egd_top.BitStream_buffer.BitStream_buffer_output\[9\]
+ vssd1 vssd1 vccd1 vccd1 _2714_ sky130_fd_sc_hd__nand2_1
XFILLER_88_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6274_ _2627_ egd_top.BitStream_buffer.BitStream_buffer_output\[1\] vssd1 vssd1 vccd1
+ vccd1 _2645_ sky130_fd_sc_hd__nand2_1
X_3486_ _2974_ _3021_ vssd1 vssd1 vccd1 vccd1 _3022_ sky130_fd_sc_hd__nand2_1
X_5225_ _3332_ _3040_ vssd1 vssd1 vccd1 vccd1 _1730_ sky130_fd_sc_hd__nand2_1
XFILLER_56_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5156_ _0442_ _0467_ vssd1 vssd1 vccd1 vccd1 _1662_ sky130_fd_sc_hd__nand2_1
XFILLER_84_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4107_ _0620_ vssd1 vssd1 vccd1 vccd1 _0621_ sky130_fd_sc_hd__clkbuf_2
X_5087_ _0727_ _3106_ vssd1 vssd1 vccd1 vccd1 _1593_ sky130_fd_sc_hd__or2_1
XFILLER_29_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4038_ _0501_ _0518_ _0536_ _0551_ vssd1 vssd1 vccd1 vccd1 _0552_ sky130_fd_sc_hd__and4_1
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5989_ _2466_ _0922_ vssd1 vssd1 vccd1 vccd1 _2468_ sky130_fd_sc_hd__nand2_1
XFILLER_12_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5010_ _0609_ _0505_ vssd1 vssd1 vccd1 vccd1 _1517_ sky130_fd_sc_hd__nand2_1
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5912_ _2403_ _2406_ _2408_ _2411_ vssd1 vssd1 vccd1 vccd1 _2412_ sky130_fd_sc_hd__and4_1
X_5843_ _3309_ _3094_ vssd1 vssd1 vccd1 vccd1 _2343_ sky130_fd_sc_hd__nand2_1
XFILLER_21_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5774_ _0585_ _3176_ _0583_ _3180_ _2274_ vssd1 vssd1 vccd1 vccd1 _2275_ sky130_fd_sc_hd__a221oi_1
X_4725_ _0808_ _3122_ _1231_ _1232_ _1233_ vssd1 vssd1 vccd1 vccd1 _1234_ sky130_fd_sc_hd__o2111a_1
X_4656_ _3332_ _0330_ vssd1 vssd1 vccd1 vccd1 _1166_ sky130_fd_sc_hd__nand2_1
X_3607_ _3140_ vssd1 vssd1 vccd1 vccd1 _3141_ sky130_fd_sc_hd__buf_6
X_4587_ _0457_ _0478_ vssd1 vssd1 vccd1 vccd1 _1097_ sky130_fd_sc_hd__nand2_1
X_3538_ _3071_ vssd1 vssd1 vccd1 vccd1 _3072_ sky130_fd_sc_hd__clkinv_2
X_6326_ net18 net17 vssd1 vssd1 vccd1 vccd1 _2697_ sky130_fd_sc_hd__nand2_1
X_6257_ _2626_ _2627_ vssd1 vssd1 vccd1 vccd1 _2628_ sky130_fd_sc_hd__nand2_1
X_3469_ egd_top.BitStream_buffer.BS_buffer\[122\] vssd1 vssd1 vccd1 vccd1 _3009_ sky130_fd_sc_hd__clkinv_2
X_5208_ _3038_ _0722_ vssd1 vssd1 vccd1 vccd1 _1713_ sky130_fd_sc_hd__nand2_1
X_6188_ egd_top.BitStream_buffer.pc_previous\[6\] _2587_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.pc\[6\]
+ sky130_fd_sc_hd__xor2_4
XFILLER_29_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5139_ _1617_ _1644_ vssd1 vssd1 vccd1 vccd1 _1645_ sky130_fd_sc_hd__nor2_1
XFILLER_72_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_525 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6578__120 clknet_1_0__leaf__2888_ vssd1 vssd1 vccd1 vccd1 net154 sky130_fd_sc_hd__inv_2
X_4510_ _3098_ _0722_ vssd1 vssd1 vccd1 vccd1 _1021_ sky130_fd_sc_hd__nand2_1
XFILLER_7_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5490_ _1980_ _1984_ _1989_ _1992_ vssd1 vssd1 vccd1 vccd1 _1993_ sky130_fd_sc_hd__and4_1
X_4441_ _0939_ _0943_ _0947_ _0951_ vssd1 vssd1 vccd1 vccd1 _0952_ sky130_fd_sc_hd__and4_1
XFILLER_7_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6111_ _2538_ _1043_ vssd1 vssd1 vccd1 vccd1 _2539_ sky130_fd_sc_hd__nand2_1
X_4372_ _0442_ _0429_ vssd1 vssd1 vccd1 vccd1 _0884_ sky130_fd_sc_hd__nand2_1
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6042_ _2998_ _2487_ _2488_ _2498_ vssd1 vssd1 vccd1 vccd1 _0240_ sky130_fd_sc_hd__o211a_1
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5826_ _2977_ _3056_ _2323_ _2324_ _2325_ vssd1 vssd1 vccd1 vccd1 _2326_ sky130_fd_sc_hd__o2111a_1
XFILLER_22_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5757_ _3198_ _3113_ _3117_ _0744_ _2257_ vssd1 vssd1 vccd1 vccd1 _2258_ sky130_fd_sc_hd__a221oi_1
X_4708_ _0779_ _3318_ vssd1 vssd1 vccd1 vccd1 _1217_ sky130_fd_sc_hd__or2_1
X_5688_ _2072_ _2189_ vssd1 vssd1 vccd1 vccd1 _0285_ sky130_fd_sc_hd__nor2_1
X_4639_ egd_top.BitStream_buffer.BS_buffer\[76\] vssd1 vssd1 vccd1 vccd1 _1149_ sky130_fd_sc_hd__clkinv_2
XFILLER_89_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6309_ egd_top.BitStream_buffer.BitStream_buffer_output\[1\] _2678_ _2679_ vssd1
+ vssd1 vccd1 vccd1 _2680_ sky130_fd_sc_hd__o21ai_2
XFILLER_1_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__2898_ clknet_0__2898_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__2898_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_63_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4990_ _0995_ _0530_ _0366_ _0534_ vssd1 vssd1 vccd1 vccd1 _1497_ sky130_fd_sc_hd__o22a_1
X_3941_ _0453_ _0454_ vssd1 vssd1 vccd1 vccd1 _0455_ sky130_fd_sc_hd__nand2_1
XFILLER_90_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3872_ _3110_ _0338_ vssd1 vssd1 vccd1 vccd1 _0386_ sky130_fd_sc_hd__and2_1
X_5611_ _0528_ _0612_ vssd1 vssd1 vccd1 vccd1 _2113_ sky130_fd_sc_hd__or2_1
X_6591_ clknet_1_1__leaf__2883_ vssd1 vssd1 vccd1 vccd1 _2890_ sky130_fd_sc_hd__buf_1
X_5542_ _0540_ _0504_ egd_top.BitStream_buffer.BS_buffer\[32\] _0508_ _2044_ vssd1
+ vssd1 vccd1 vccd1 _2045_ sky130_fd_sc_hd__a221oi_1
X_5473_ _3149_ _0726_ _3133_ _3080_ _1975_ vssd1 vssd1 vccd1 vccd1 _1976_ sky130_fd_sc_hd__a221oi_1
X_4424_ egd_top.BitStream_buffer.BitStream_buffer_output\[12\] _2965_ _0627_ vssd1
+ vssd1 vccd1 vccd1 _0935_ sky130_fd_sc_hd__o21ai_1
X_4355_ _0865_ _0368_ _0866_ vssd1 vssd1 vccd1 vccd1 _0867_ sky130_fd_sc_hd__o21ai_1
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_447 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4286_ _0796_ _3056_ _0797_ vssd1 vssd1 vccd1 vccd1 _0798_ sky130_fd_sc_hd__o21ai_1
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6025_ _2486_ vssd1 vssd1 vccd1 vccd1 _2489_ sky130_fd_sc_hd__buf_2
XFILLER_27_514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6858_ net102 _0317_ vssd1 vssd1 vccd1 vccd1 net30 sky130_fd_sc_hd__dfxtp_2
XFILLER_22_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5809_ egd_top.BitStream_buffer.BitStream_buffer_output\[1\] _2964_ _0627_ vssd1
+ vssd1 vccd1 vccd1 _2309_ sky130_fd_sc_hd__o21ai_1
X_6789_ net193 _0248_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_89_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4140_ egd_top.BitStream_buffer.BS_buffer\[54\] vssd1 vssd1 vccd1 vccd1 _0653_ sky130_fd_sc_hd__clkinv_2
XFILLER_68_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4071_ egd_top.BitStream_buffer.BS_buffer\[9\] vssd1 vssd1 vccd1 vccd1 _0585_ sky130_fd_sc_hd__clkbuf_4
XFILLER_63_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4973_ _0883_ _0425_ vssd1 vssd1 vccd1 vccd1 _1480_ sky130_fd_sc_hd__or2_1
X_6712_ net116 _0171_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[85\]
+ sky130_fd_sc_hd__dfxtp_1
X_3924_ _3104_ _2934_ vssd1 vssd1 vccd1 vccd1 _0438_ sky130_fd_sc_hd__nand2_2
X_3855_ _3033_ _0338_ vssd1 vssd1 vccd1 vccd1 _0369_ sky130_fd_sc_hd__and2_1
X_3786_ _3317_ _3319_ vssd1 vssd1 vccd1 vccd1 _3320_ sky130_fd_sc_hd__or2_1
X_5525_ _0442_ _0664_ vssd1 vssd1 vccd1 vccd1 _2028_ sky130_fd_sc_hd__nand2_1
X_5456_ _0328_ _0714_ vssd1 vssd1 vccd1 vccd1 _1959_ sky130_fd_sc_hd__nand2_1
X_4407_ _0611_ _0576_ _0916_ _0917_ _0918_ vssd1 vssd1 vccd1 vccd1 _0919_ sky130_fd_sc_hd__o2111a_1
X_5387_ _0330_ _3292_ _0785_ _3295_ _1890_ vssd1 vssd1 vccd1 vccd1 _1891_ sky130_fd_sc_hd__a221oi_1
XFILLER_59_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4338_ egd_top.BitStream_buffer.BS_buffer\[91\] vssd1 vssd1 vccd1 vccd1 _0850_ sky130_fd_sc_hd__clkinv_2
X_4269_ _0779_ _3330_ _0781_ vssd1 vssd1 vccd1 vccd1 _0782_ sky130_fd_sc_hd__o21ai_1
XFILLER_86_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6008_ _3005_ _2465_ _2474_ _2478_ vssd1 vssd1 vccd1 vccd1 _0254_ sky130_fd_sc_hd__o211a_1
XFILLER_82_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3640_ _3067_ _3134_ vssd1 vssd1 vccd1 vccd1 _3174_ sky130_fd_sc_hd__and2_1
X_3571_ _3104_ _3036_ vssd1 vssd1 vccd1 vccd1 _3105_ sky130_fd_sc_hd__nand2_2
X_5310_ _0582_ _0498_ vssd1 vssd1 vccd1 vccd1 _1815_ sky130_fd_sc_hd__nand2_1
XFILLER_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6290_ egd_top.BitStream_buffer.BitStream_buffer_output\[11\] _2660_ vssd1 vssd1
+ vccd1 vccd1 _2661_ sky130_fd_sc_hd__or2_1
XFILLER_5_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5241_ _3215_ _3272_ vssd1 vssd1 vccd1 vccd1 _1746_ sky130_fd_sc_hd__nand2_1
X_5172_ _0907_ _0512_ _1677_ vssd1 vssd1 vccd1 vccd1 _1678_ sky130_fd_sc_hd__o21ai_1
X_4123_ _0364_ _0359_ _0362_ _0337_ _0635_ vssd1 vssd1 vccd1 vccd1 _0636_ sky130_fd_sc_hd__a221oi_1
XFILLER_83_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput2 la_data_in_58_43[10] vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__clkbuf_1
X_4054_ egd_top.BitStream_buffer.BS_buffer\[5\] vssd1 vssd1 vccd1 vccd1 _0568_ sky130_fd_sc_hd__buf_4
XFILLER_83_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4956_ _1394_ _1462_ _1463_ vssd1 vssd1 vccd1 vccd1 _1464_ sky130_fd_sc_hd__nand3_1
XFILLER_61_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3907_ _3045_ _2934_ vssd1 vssd1 vccd1 vccd1 _0421_ sky130_fd_sc_hd__nand2_2
X_4887_ _3332_ _3338_ vssd1 vssd1 vccd1 vccd1 _1395_ sky130_fd_sc_hd__nand2_1
X_3838_ _0351_ vssd1 vssd1 vccd1 vccd1 _0352_ sky130_fd_sc_hd__inv_2
X_5508_ _1962_ _1977_ _1993_ _2010_ vssd1 vssd1 vccd1 vccd1 _2011_ sky130_fd_sc_hd__and4_1
X_3769_ _3301_ _3302_ vssd1 vssd1 vccd1 vccd1 _3303_ sky130_fd_sc_hd__nand2_1
X_6488_ _2848_ _2923_ _2850_ vssd1 vssd1 vccd1 vccd1 _2851_ sky130_fd_sc_hd__nand3_1
XFILLER_10_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5439_ _0622_ _0583_ vssd1 vssd1 vccd1 vccd1 _1943_ sky130_fd_sc_hd__nand2_1
XFILLER_87_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4810_ _0582_ egd_top.BitStream_buffer.BS_buffer\[15\] vssd1 vssd1 vccd1 vccd1 _1319_
+ sky130_fd_sc_hd__nand2_1
XFILLER_33_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5790_ _0324_ _3299_ _2290_ vssd1 vssd1 vccd1 vccd1 _2291_ sky130_fd_sc_hd__o21ai_1
X_4741_ _1248_ _1249_ vssd1 vssd1 vccd1 vccd1 _1250_ sky130_fd_sc_hd__nand2_1
X_4672_ _0727_ _3123_ _1181_ vssd1 vssd1 vccd1 vccd1 _1182_ sky130_fd_sc_hd__o21ai_1
X_3623_ egd_top.BitStream_buffer.BS_buffer\[115\] vssd1 vssd1 vccd1 vccd1 _3157_ sky130_fd_sc_hd__clkbuf_4
X_6411_ egd_top.BitStream_buffer.BitStream_buffer_output\[10\] _2753_ vssd1 vssd1
+ vccd1 vccd1 _2780_ sky130_fd_sc_hd__xnor2_1
X_6555__99 clknet_1_0__leaf__2886_ vssd1 vssd1 vccd1 vccd1 net133 sky130_fd_sc_hd__inv_2
X_3554_ _3087_ _3036_ vssd1 vssd1 vccd1 vccd1 _3088_ sky130_fd_sc_hd__nand2_2
X_6342_ _2712_ vssd1 vssd1 vccd1 vccd1 _2713_ sky130_fd_sc_hd__inv_2
X_3485_ egd_top.BitStream_buffer.BS_buffer\[126\] vssd1 vssd1 vccd1 vccd1 _3021_ sky130_fd_sc_hd__inv_2
X_6273_ _2625_ _2643_ vssd1 vssd1 vccd1 vccd1 _2644_ sky130_fd_sc_hd__nor2_1
X_5224_ _0784_ _3319_ _1726_ _1727_ _1728_ vssd1 vssd1 vccd1 vccd1 _1729_ sky130_fd_sc_hd__o2111a_1
XFILLER_84_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5155_ _0459_ _0415_ _0447_ _0419_ _1660_ vssd1 vssd1 vccd1 vccd1 _1661_ sky130_fd_sc_hd__a221oi_1
X_4106_ _0619_ _2932_ _3211_ _3034_ vssd1 vssd1 vccd1 vccd1 _0620_ sky130_fd_sc_hd__and4_1
X_5086_ _3099_ _3075_ vssd1 vssd1 vccd1 vccd1 _1592_ sky130_fd_sc_hd__nand2_1
XFILLER_56_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4037_ _0537_ _0539_ _0540_ _0542_ _0550_ vssd1 vssd1 vccd1 vccd1 _0551_ sky130_fd_sc_hd__a221oi_1
XFILLER_71_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5988_ _2966_ _2465_ _2458_ _2467_ vssd1 vssd1 vccd1 vccd1 _0263_ sky130_fd_sc_hd__o211a_1
X_4939_ _3012_ _3199_ _1444_ _1445_ _1446_ vssd1 vssd1 vccd1 vccd1 _1447_ sky130_fd_sc_hd__o2111a_1
XFILLER_52_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_534 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5911_ _0393_ _0539_ _0400_ _0542_ _2410_ vssd1 vssd1 vccd1 vccd1 _2411_ sky130_fd_sc_hd__a221oi_1
XFILLER_19_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5842_ _3313_ _0708_ vssd1 vssd1 vccd1 vccd1 _2342_ sky130_fd_sc_hd__nand2_1
XFILLER_34_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5773_ _0574_ _3183_ _2273_ vssd1 vssd1 vccd1 vccd1 _2274_ sky130_fd_sc_hd__o21ai_1
X_4724_ _3116_ _3169_ vssd1 vssd1 vccd1 vccd1 _1233_ sky130_fd_sc_hd__nand2_1
XFILLER_21_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4655_ _0850_ _3308_ _1162_ _1163_ _1164_ vssd1 vssd1 vccd1 vccd1 _1165_ sky130_fd_sc_hd__o2111a_1
X_3606_ _3139_ vssd1 vssd1 vccd1 vccd1 _3140_ sky130_fd_sc_hd__clkbuf_2
X_4586_ _1083_ _1088_ _1092_ _1095_ vssd1 vssd1 vccd1 vccd1 _1096_ sky130_fd_sc_hd__and4_1
X_3537_ _2920_ _3042_ vssd1 vssd1 vccd1 vccd1 _3071_ sky130_fd_sc_hd__nor2_4
X_6325_ net21 egd_top.exp_golomb_decoding.te_range\[2\] net20 vssd1 vssd1 vccd1 vccd1
+ _2696_ sky130_fd_sc_hd__nor3b_1
X_6256_ egd_top.BitStream_buffer.BitStream_buffer_output\[2\] vssd1 vssd1 vccd1 vccd1
+ _2627_ sky130_fd_sc_hd__inv_2
X_3468_ net12 vssd1 vssd1 vccd1 vccd1 _3008_ sky130_fd_sc_hd__clkbuf_4
XFILLER_76_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5207_ _3157_ _3113_ _3117_ _3204_ _1711_ vssd1 vssd1 vccd1 vccd1 _1712_ sky130_fd_sc_hd__a221oi_1
XFILLER_69_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3399_ _2916_ _2915_ vssd1 vssd1 vccd1 vccd1 _2953_ sky130_fd_sc_hd__nor2_1
X_6187_ _2575_ _2586_ vssd1 vssd1 vccd1 vccd1 _2587_ sky130_fd_sc_hd__nor2_2
XFILLER_57_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5138_ _1629_ _1643_ vssd1 vssd1 vccd1 vccd1 _1644_ sky130_fd_sc_hd__nand2_1
X_5069_ _1574_ _1145_ _1575_ vssd1 vssd1 vccd1 vccd1 _1576_ sky130_fd_sc_hd__o21ai_1
XFILLER_25_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4440_ _0642_ _0396_ _0399_ _0874_ _0950_ vssd1 vssd1 vccd1 vccd1 _0951_ sky130_fd_sc_hd__a221oi_2
X_6110_ _2531_ vssd1 vssd1 vccd1 vccd1 _2538_ sky130_fd_sc_hd__buf_2
X_4371_ _0436_ vssd1 vssd1 vccd1 vccd1 _0883_ sky130_fd_sc_hd__clkinv_2
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6694__65 clknet_1_1__leaf__2899_ vssd1 vssd1 vccd1 vccd1 net99 sky130_fd_sc_hd__inv_2
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6041_ _2494_ _0348_ vssd1 vssd1 vccd1 vccd1 _2498_ sky130_fd_sc_hd__nand2_1
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5825_ _3061_ _3164_ vssd1 vssd1 vccd1 vccd1 _2325_ sky130_fd_sc_hd__nand2_1
X_5756_ _2996_ _3123_ _2256_ vssd1 vssd1 vccd1 vccd1 _2257_ sky130_fd_sc_hd__o21ai_1
X_5687_ _3026_ _2188_ vssd1 vssd1 vccd1 vccd1 _2189_ sky130_fd_sc_hd__nor2_1
X_4707_ _3310_ _3327_ vssd1 vssd1 vccd1 vccd1 _1216_ sky130_fd_sc_hd__nand2_1
X_4638_ _3256_ _3216_ _3264_ _3220_ _1147_ vssd1 vssd1 vccd1 vccd1 _1148_ sky130_fd_sc_hd__a221oi_1
X_4569_ _0935_ _1079_ vssd1 vssd1 vccd1 vccd1 _0294_ sky130_fd_sc_hd__nor2_1
X_6308_ _2678_ _2626_ vssd1 vssd1 vccd1 vccd1 _2679_ sky130_fd_sc_hd__nand2_1
XFILLER_89_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6239_ _2608_ _0779_ vssd1 vssd1 vccd1 vccd1 _2616_ sky130_fd_sc_hd__nand2_1
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f__2897_ clknet_0__2897_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__2897_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_48_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3940_ egd_top.BitStream_buffer.BS_buffer\[56\] vssd1 vssd1 vccd1 vccd1 _0454_ sky130_fd_sc_hd__buf_2
XFILLER_16_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3871_ _0384_ vssd1 vssd1 vccd1 vccd1 _0385_ sky130_fd_sc_hd__clkbuf_4
XFILLER_83_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5610_ _0605_ _0519_ vssd1 vssd1 vccd1 vccd1 _2112_ sky130_fd_sc_hd__nand2_1
X_5541_ _0633_ _0512_ _2043_ vssd1 vssd1 vccd1 vccd1 _2044_ sky130_fd_sc_hd__o21ai_1
XFILLER_8_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5472_ _2999_ _0729_ _1974_ vssd1 vssd1 vccd1 vccd1 _1975_ sky130_fd_sc_hd__o21ai_1
X_4423_ _3027_ _0932_ _0934_ vssd1 vssd1 vccd1 vccd1 _0295_ sky130_fd_sc_hd__o21a_1
X_4354_ _0371_ egd_top.BitStream_buffer.BS_buffer\[34\] vssd1 vssd1 vccd1 vccd1 _0866_
+ sky130_fd_sc_hd__nand2_1
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4285_ _3061_ _0716_ vssd1 vssd1 vccd1 vccd1 _0797_ sky130_fd_sc_hd__nand2_1
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6024_ _2904_ vssd1 vssd1 vccd1 vccd1 _2488_ sky130_fd_sc_hd__buf_2
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6857_ net101 _0316_ vssd1 vssd1 vccd1 vccd1 net29 sky130_fd_sc_hd__dfxtp_2
XFILLER_10_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6788_ net192 _0247_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[32\]
+ sky130_fd_sc_hd__dfxtp_4
X_5808_ _2190_ _2308_ vssd1 vssd1 vccd1 vccd1 _0284_ sky130_fd_sc_hd__nor2_1
X_5739_ _0901_ _0337_ vssd1 vssd1 vccd1 vccd1 _2240_ sky130_fd_sc_hd__nand2_1
XFILLER_13_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6658__32 clknet_1_0__leaf__2896_ vssd1 vssd1 vccd1 vccd1 net66 sky130_fd_sc_hd__inv_2
XFILLER_38_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6673__46 clknet_1_0__leaf__2897_ vssd1 vssd1 vccd1 vccd1 net80 sky130_fd_sc_hd__inv_2
XFILLER_57_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6616__154 clknet_1_0__leaf__2892_ vssd1 vssd1 vccd1 vccd1 net188 sky130_fd_sc_hd__inv_2
XFILLER_68_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4070_ _0582_ _0583_ vssd1 vssd1 vccd1 vccd1 _0584_ sky130_fd_sc_hd__nand2_1
XFILLER_83_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4972_ _1469_ _1472_ _1475_ _1478_ vssd1 vssd1 vccd1 vccd1 _1479_ sky130_fd_sc_hd__and4_1
XFILLER_24_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3923_ egd_top.BitStream_buffer.BS_buffer\[53\] vssd1 vssd1 vccd1 vccd1 _0437_ sky130_fd_sc_hd__inv_2
X_6711_ net115 _0170_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[86\]
+ sky130_fd_sc_hd__dfxtp_1
X_3854_ _0367_ vssd1 vssd1 vccd1 vccd1 _0368_ sky130_fd_sc_hd__buf_2
X_3785_ _3318_ vssd1 vssd1 vccd1 vccd1 _3319_ sky130_fd_sc_hd__buf_2
X_5524_ _0471_ _0415_ _0478_ _0419_ _2026_ vssd1 vssd1 vccd1 vccd1 _2027_ sky130_fd_sc_hd__a221oi_1
X_5455_ _3049_ _3308_ _1955_ _1956_ _1957_ vssd1 vssd1 vccd1 vccd1 _1958_ sky130_fd_sc_hd__o2111a_1
X_4406_ _0574_ _0588_ vssd1 vssd1 vccd1 vccd1 _0918_ sky130_fd_sc_hd__or2_1
X_5386_ _0779_ _3299_ _1889_ vssd1 vssd1 vccd1 vccd1 _1890_ sky130_fd_sc_hd__o21ai_1
X_4337_ _3328_ _3308_ _0846_ _0847_ _0848_ vssd1 vssd1 vccd1 vccd1 _0849_ sky130_fd_sc_hd__o2111a_1
XFILLER_75_18 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4268_ _3333_ _0780_ vssd1 vssd1 vccd1 vccd1 _0781_ sky130_fd_sc_hd__nand2_1
XFILLER_67_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6007_ _2471_ _0528_ vssd1 vssd1 vccd1 vccd1 _2478_ sky130_fd_sc_hd__nand2_1
X_4199_ _3040_ _3039_ _0708_ _3048_ _0711_ vssd1 vssd1 vccd1 vccd1 _0712_ sky130_fd_sc_hd__a221oi_1
XFILLER_27_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_0__2899_ _2899_ vssd1 vssd1 vccd1 vccd1 clknet_0__2899_ sky130_fd_sc_hd__clkbuf_16
XFILLER_24_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3570_ _3103_ vssd1 vssd1 vccd1 vccd1 _3104_ sky130_fd_sc_hd__buf_6
XFILLER_5_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5240_ _0833_ _3240_ _1742_ _1743_ _1744_ vssd1 vssd1 vccd1 vccd1 _1745_ sky130_fd_sc_hd__o2111a_1
XFILLER_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5171_ _0514_ _0537_ vssd1 vssd1 vccd1 vccd1 _1677_ sky130_fd_sc_hd__nand2_1
XFILLER_68_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6637__13 clknet_1_1__leaf__2894_ vssd1 vssd1 vccd1 vccd1 net47 sky130_fd_sc_hd__inv_2
X_4122_ _0633_ _0367_ _0634_ vssd1 vssd1 vccd1 vccd1 _0635_ sky130_fd_sc_hd__o21ai_1
X_4053_ _0565_ _0566_ vssd1 vssd1 vccd1 vccd1 _0567_ sky130_fd_sc_hd__nand2_1
XFILLER_56_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6652__27 clknet_1_1__leaf__2895_ vssd1 vssd1 vccd1 vccd1 net61 sky130_fd_sc_hd__inv_2
XFILLER_83_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput3 la_data_in_58_43[11] vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__clkbuf_1
XFILLER_64_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4955_ _0622_ _0562_ vssd1 vssd1 vccd1 vccd1 _1463_ sky130_fd_sc_hd__nand2_1
XFILLER_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3906_ egd_top.BitStream_buffer.BS_buffer\[49\] vssd1 vssd1 vccd1 vccd1 _0420_ sky130_fd_sc_hd__clkinv_2
XFILLER_51_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4886_ _1348_ _1364_ _1379_ _1393_ vssd1 vssd1 vccd1 vccd1 _1394_ sky130_fd_sc_hd__and4_1
X_3837_ _3096_ _0339_ vssd1 vssd1 vccd1 vccd1 _0351_ sky130_fd_sc_hd__nand2_1
X_3768_ egd_top.BitStream_buffer.BS_buffer\[81\] vssd1 vssd1 vccd1 vccd1 _3302_ sky130_fd_sc_hd__clkbuf_4
X_5507_ _1996_ _2001_ _2006_ _2009_ vssd1 vssd1 vccd1 vccd1 _2010_ sky130_fd_sc_hd__and4_1
X_6487_ _2835_ _2849_ _2836_ vssd1 vssd1 vccd1 vccd1 _2850_ sky130_fd_sc_hd__nand3_1
X_3699_ _3232_ vssd1 vssd1 vccd1 vccd1 _3233_ sky130_fd_sc_hd__clkbuf_4
X_5438_ _1913_ _1941_ vssd1 vssd1 vccd1 vccd1 _1942_ sky130_fd_sc_hd__nor2_1
X_5369_ _0578_ _0491_ vssd1 vssd1 vccd1 vccd1 _1873_ sky130_fd_sc_hd__nand2_1
XFILLER_59_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_167 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4740_ _3168_ egd_top.BitStream_buffer.BS_buffer\[117\] vssd1 vssd1 vccd1 vccd1 _1249_
+ sky130_fd_sc_hd__nand2_1
X_4671_ _3127_ _3066_ vssd1 vssd1 vccd1 vccd1 _1181_ sky130_fd_sc_hd__nand2_1
X_3622_ _3155_ vssd1 vssd1 vccd1 vccd1 _3156_ sky130_fd_sc_hd__buf_2
X_6410_ _2774_ _2778_ _2681_ vssd1 vssd1 vccd1 vccd1 _2779_ sky130_fd_sc_hd__nand3_1
X_6341_ egd_top.BitStream_buffer.BitStream_buffer_output\[10\] egd_top.BitStream_buffer.BitStream_buffer_output\[9\]
+ vssd1 vssd1 vccd1 vccd1 _2712_ sky130_fd_sc_hd__nor2_1
X_3553_ _3086_ vssd1 vssd1 vccd1 vccd1 _3087_ sky130_fd_sc_hd__buf_6
X_6272_ _2630_ _2637_ _2642_ vssd1 vssd1 vccd1 vccd1 _2643_ sky130_fd_sc_hd__o21ai_2
X_3484_ net8 vssd1 vssd1 vccd1 vccd1 _3020_ sky130_fd_sc_hd__buf_4
X_5223_ _1016_ _3307_ vssd1 vssd1 vccd1 vccd1 _1728_ sky130_fd_sc_hd__or2_1
X_5154_ _0462_ _0422_ _1659_ vssd1 vssd1 vccd1 vccd1 _1660_ sky130_fd_sc_hd__o21ai_1
X_4105_ _2929_ _3031_ _3032_ _2921_ _0559_ vssd1 vssd1 vccd1 vccd1 _0619_ sky130_fd_sc_hd__a41o_1
X_5085_ _3093_ _3066_ vssd1 vssd1 vccd1 vccd1 _1591_ sky130_fd_sc_hd__nand2_1
X_4036_ _0543_ _0546_ _0549_ vssd1 vssd1 vccd1 vccd1 _0550_ sky130_fd_sc_hd__o21ai_1
XFILLER_56_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5987_ _2466_ _0685_ vssd1 vssd1 vccd1 vccd1 _2467_ sky130_fd_sc_hd__nand2_1
X_4938_ _3196_ _3177_ vssd1 vssd1 vccd1 vccd1 _1446_ sky130_fd_sc_hd__nand2_1
X_4869_ _0692_ _0612_ vssd1 vssd1 vccd1 vccd1 _1377_ sky130_fd_sc_hd__or2_1
XFILLER_20_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5910_ _0383_ _0546_ _2409_ vssd1 vssd1 vccd1 vccd1 _2410_ sky130_fd_sc_hd__o21ai_1
XFILLER_34_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5841_ _3128_ _3323_ _3325_ _0722_ _2340_ vssd1 vssd1 vccd1 vccd1 _2341_ sky130_fd_sc_hd__a221oi_1
X_5772_ _3186_ egd_top.BitStream_buffer.BS_buffer\[12\] vssd1 vssd1 vccd1 vccd1 _2273_
+ sky130_fd_sc_hd__nand2_1
X_4723_ _3112_ _3082_ vssd1 vssd1 vccd1 vccd1 _1232_ sky130_fd_sc_hd__nand2_1
XFILLER_21_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4654_ _3328_ _3318_ vssd1 vssd1 vccd1 vccd1 _1164_ sky130_fd_sc_hd__or2_1
X_3605_ _3114_ _3134_ vssd1 vssd1 vccd1 vccd1 _3139_ sky130_fd_sc_hd__and2_1
X_4585_ egd_top.BitStream_buffer.BS_buffer\[48\] _0395_ _0398_ egd_top.BitStream_buffer.BS_buffer\[49\]
+ _1094_ vssd1 vssd1 vccd1 vccd1 _1095_ sky130_fd_sc_hd__a221oi_1
X_3536_ egd_top.BitStream_buffer.BS_buffer\[109\] vssd1 vssd1 vccd1 vccd1 _3070_ sky130_fd_sc_hd__clkbuf_4
X_6324_ _2694_ _2684_ vssd1 vssd1 vccd1 vccd1 _2695_ sky130_fd_sc_hd__nand2_2
XFILLER_88_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6255_ egd_top.BitStream_buffer.BitStream_buffer_output\[3\] vssd1 vssd1 vccd1 vccd1
+ _2626_ sky130_fd_sc_hd__inv_2
XFILLER_88_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5206_ _2983_ _3123_ _1710_ vssd1 vssd1 vccd1 vccd1 _1711_ sky130_fd_sc_hd__o21ai_1
X_3467_ _3005_ _2975_ _3002_ _3007_ vssd1 vssd1 vccd1 vccd1 _0304_ sky130_fd_sc_hd__o211a_1
X_3398_ net30 net28 vssd1 vssd1 vccd1 vccd1 _2952_ sky130_fd_sc_hd__nor2_1
X_6186_ _2585_ egd_top.BitStream_buffer.pc_previous\[4\] vssd1 vssd1 vccd1 vccd1 _2586_
+ sky130_fd_sc_hd__nand2_1
X_5137_ _1632_ _1636_ _1639_ _1642_ vssd1 vssd1 vccd1 vccd1 _1643_ sky130_fd_sc_hd__and4_1
X_5068_ _3224_ _3272_ vssd1 vssd1 vccd1 vccd1 _1575_ sky130_fd_sc_hd__nand2_1
XFILLER_84_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4019_ _0521_ _3051_ vssd1 vssd1 vccd1 vccd1 _0533_ sky130_fd_sc_hd__nand2_2
XFILLER_16_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6610__149 clknet_1_1__leaf__2891_ vssd1 vssd1 vccd1 vccd1 net183 sky130_fd_sc_hd__inv_2
XFILLER_87_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4370_ _0443_ _0415_ _0655_ _0419_ _0881_ vssd1 vssd1 vccd1 vccd1 _0882_ sky130_fd_sc_hd__a221oi_1
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6585__126 clknet_1_0__leaf__2889_ vssd1 vssd1 vccd1 vccd1 net160 sky130_fd_sc_hd__inv_2
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6040_ _2995_ _2487_ _2488_ _2497_ vssd1 vssd1 vccd1 vccd1 _0241_ sky130_fd_sc_hd__o211a_1
XFILLER_85_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5824_ _3047_ _3082_ vssd1 vssd1 vccd1 vccd1 _2324_ sky130_fd_sc_hd__nand2_1
XFILLER_22_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5755_ _3127_ _0746_ vssd1 vssd1 vccd1 vccd1 _2256_ sky130_fd_sc_hd__nand2_1
X_5686_ _2130_ _2186_ _2187_ vssd1 vssd1 vccd1 vccd1 _2188_ sky130_fd_sc_hd__nand3_1
X_4706_ _3314_ _0780_ vssd1 vssd1 vccd1 vccd1 _1215_ sky130_fd_sc_hd__nand2_1
XFILLER_8_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4637_ _1144_ _1145_ _1146_ vssd1 vssd1 vccd1 vccd1 _1147_ sky130_fd_sc_hd__o21ai_1
XFILLER_89_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4568_ _3026_ _1078_ vssd1 vssd1 vccd1 vccd1 _1079_ sky130_fd_sc_hd__nor2_1
X_3519_ _3052_ vssd1 vssd1 vccd1 vccd1 _3053_ sky130_fd_sc_hd__inv_2
X_6307_ _2658_ _2677_ _2623_ vssd1 vssd1 vccd1 vccd1 _2678_ sky130_fd_sc_hd__nand3_4
X_4499_ _3300_ _3315_ vssd1 vssd1 vccd1 vccd1 _1010_ sky130_fd_sc_hd__nand2_1
X_6238_ _3005_ _2602_ _2611_ _2615_ vssd1 vssd1 vccd1 vccd1 _0167_ sky130_fd_sc_hd__o211a_1
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6169_ _2561_ _0727_ vssd1 vssd1 vccd1 vccd1 _2572_ sky130_fd_sc_hd__nand2_1
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__2896_ clknet_0__2896_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__2896_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_48_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_398 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3870_ _3114_ _0339_ vssd1 vssd1 vccd1 vccd1 _0384_ sky130_fd_sc_hd__nand2_1
X_5540_ _0514_ _0365_ vssd1 vssd1 vccd1 vccd1 _2043_ sky130_fd_sc_hd__nand2_1
XFILLER_76_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5471_ _3073_ _0744_ vssd1 vssd1 vccd1 vccd1 _1974_ sky130_fd_sc_hd__nand2_1
XFILLER_8_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4422_ _0933_ _3027_ _2905_ vssd1 vssd1 vccd1 vccd1 _0934_ sky130_fd_sc_hd__a21oi_1
X_4353_ _0364_ vssd1 vssd1 vccd1 vccd1 _0865_ sky130_fd_sc_hd__inv_2
XFILLER_86_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4284_ egd_top.BitStream_buffer.BS_buffer\[100\] vssd1 vssd1 vccd1 vccd1 _0796_ sky130_fd_sc_hd__clkinv_2
XTAP_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6023_ _2486_ vssd1 vssd1 vccd1 vccd1 _2487_ sky130_fd_sc_hd__buf_2
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6856_ net100 _0315_ vssd1 vssd1 vccd1 vccd1 net28 sky130_fd_sc_hd__dfxtp_2
X_3999_ _0488_ _3097_ vssd1 vssd1 vccd1 vccd1 _0513_ sky130_fd_sc_hd__nor2_2
XFILLER_10_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6787_ net191 _0246_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[33\]
+ sky130_fd_sc_hd__dfxtp_1
X_5807_ _3026_ _2307_ vssd1 vssd1 vccd1 vccd1 _2308_ sky130_fd_sc_hd__nor2_1
X_5738_ _0503_ _0365_ vssd1 vssd1 vccd1 vccd1 _2239_ sky130_fd_sc_hd__nand2_1
XFILLER_13_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5669_ _3061_ _3082_ vssd1 vssd1 vccd1 vccd1 _2171_ sky130_fd_sc_hd__nand2_1
XFILLER_89_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4971_ _0416_ _0396_ _0399_ _0443_ _1477_ vssd1 vssd1 vccd1 vccd1 _1478_ sky130_fd_sc_hd__a221oi_2
X_6710_ net114 _0169_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[87\]
+ sky130_fd_sc_hd__dfxtp_1
X_3922_ egd_top.BitStream_buffer.BS_buffer\[55\] vssd1 vssd1 vccd1 vccd1 _0436_ sky130_fd_sc_hd__clkbuf_4
X_3853_ _3045_ _0339_ vssd1 vssd1 vccd1 vccd1 _0367_ sky130_fd_sc_hd__nand2_2
X_3784_ _3104_ _3297_ vssd1 vssd1 vccd1 vccd1 _3318_ sky130_fd_sc_hd__nand2_2
X_5523_ _0647_ _0422_ _2025_ vssd1 vssd1 vccd1 vccd1 _2026_ sky130_fd_sc_hd__o21ai_1
X_5454_ _1016_ _3318_ vssd1 vssd1 vccd1 vccd1 _1957_ sky130_fd_sc_hd__or2_1
X_4405_ _0582_ egd_top.BitStream_buffer.BS_buffer\[12\] vssd1 vssd1 vccd1 vccd1 _0917_
+ sky130_fd_sc_hd__nand2_1
X_5385_ _3301_ _3327_ vssd1 vssd1 vccd1 vccd1 _1889_ sky130_fd_sc_hd__nand2_1
X_4336_ _3306_ _3319_ vssd1 vssd1 vccd1 vccd1 _0848_ sky130_fd_sc_hd__or2_1
XFILLER_59_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4267_ egd_top.BitStream_buffer.BS_buffer\[89\] vssd1 vssd1 vccd1 vccd1 _0780_ sky130_fd_sc_hd__clkbuf_4
XFILLER_74_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4198_ _0709_ _3056_ _0710_ vssd1 vssd1 vccd1 vccd1 _0711_ sky130_fd_sc_hd__o21ai_1
X_6006_ _3001_ _2465_ _2474_ _2477_ vssd1 vssd1 vccd1 vccd1 _0255_ sky130_fd_sc_hd__o211a_1
XFILLER_39_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6839_ net83 _0298_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[127\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_24_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__2898_ _2898_ vssd1 vssd1 vccd1 vccd1 clknet_0__2898_ sky130_fd_sc_hd__clkbuf_16
XFILLER_50_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5170_ _0519_ _0487_ _0527_ _0490_ _1675_ vssd1 vssd1 vccd1 vccd1 _1676_ sky130_fd_sc_hd__a221oi_1
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4121_ _0370_ _0365_ vssd1 vssd1 vccd1 vccd1 _0634_ sky130_fd_sc_hd__nand2_1
X_4052_ egd_top.BitStream_buffer.BS_buffer\[4\] vssd1 vssd1 vccd1 vccd1 _0566_ sky130_fd_sc_hd__clkbuf_4
XFILLER_68_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput4 la_data_in_58_43[12] vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__clkbuf_1
XFILLER_64_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4954_ _1409_ _1425_ _1443_ _1461_ vssd1 vssd1 vccd1 vccd1 _1462_ sky130_fd_sc_hd__and4_1
XFILLER_51_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3905_ _0418_ vssd1 vssd1 vccd1 vccd1 _0419_ sky130_fd_sc_hd__buf_2
X_4885_ _1383_ _1387_ _1390_ _1392_ vssd1 vssd1 vccd1 vccd1 _1393_ sky130_fd_sc_hd__and4_1
XFILLER_20_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3836_ _0349_ vssd1 vssd1 vccd1 vccd1 _0350_ sky130_fd_sc_hd__buf_2
XFILLER_20_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6624_ clknet_1_1__leaf__2882_ vssd1 vssd1 vccd1 vccd1 _2893_ sky130_fd_sc_hd__buf_1
X_3767_ _3300_ vssd1 vssd1 vccd1 vccd1 _3301_ sky130_fd_sc_hd__buf_6
X_5506_ _3186_ _0583_ _0579_ _3180_ _2008_ vssd1 vssd1 vccd1 vccd1 _2009_ sky130_fd_sc_hd__a221oi_1
X_3698_ _3231_ vssd1 vssd1 vccd1 vccd1 _3232_ sky130_fd_sc_hd__clkbuf_2
X_6486_ _2844_ _2845_ _2926_ vssd1 vssd1 vccd1 vccd1 _2849_ sky130_fd_sc_hd__a21oi_2
X_5437_ _1927_ _1940_ vssd1 vssd1 vccd1 vccd1 _1941_ sky130_fd_sc_hd__nand2_1
XFILLER_10_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5368_ _0922_ _0558_ _1869_ _1870_ _1871_ vssd1 vssd1 vccd1 vccd1 _1872_ sky130_fd_sc_hd__o2111a_1
XFILLER_86_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5299_ _0633_ _0530_ _0865_ _0534_ vssd1 vssd1 vccd1 vccd1 _1804_ sky130_fd_sc_hd__o22a_1
X_4319_ _0829_ _3240_ _0830_ vssd1 vssd1 vccd1 vccd1 _0831_ sky130_fd_sc_hd__o21ai_1
XFILLER_19_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_271 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_32 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4670_ _0804_ _3089_ _1177_ _1178_ _1179_ vssd1 vssd1 vccd1 vccd1 _1180_ sky130_fd_sc_hd__o2111a_1
XFILLER_14_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3621_ _3154_ vssd1 vssd1 vccd1 vccd1 _3155_ sky130_fd_sc_hd__buf_2
X_3552_ _3057_ egd_top.BitStream_buffer.pc\[2\] _3032_ vssd1 vssd1 vccd1 vccd1 _3086_
+ sky130_fd_sc_hd__and3_1
X_6340_ _2710_ _2660_ vssd1 vssd1 vccd1 vccd1 _2711_ sky130_fd_sc_hd__or2_1
X_6271_ _2641_ vssd1 vssd1 vccd1 vccd1 _2642_ sky130_fd_sc_hd__inv_2
X_3483_ _3017_ _2976_ _3002_ _3019_ vssd1 vssd1 vccd1 vccd1 _0300_ sky130_fd_sc_hd__o211a_1
X_5222_ _3313_ _0785_ vssd1 vssd1 vccd1 vccd1 _1727_ sky130_fd_sc_hd__nand2_1
X_5153_ _0965_ _0425_ vssd1 vssd1 vccd1 vccd1 _1659_ sky130_fd_sc_hd__or2_1
X_4104_ _0483_ _0617_ vssd1 vssd1 vccd1 vccd1 _0618_ sky130_fd_sc_hd__nor2_1
X_5084_ _3128_ _3039_ _0722_ _3048_ _1589_ vssd1 vssd1 vccd1 vccd1 _1590_ sky130_fd_sc_hd__a221oi_2
XFILLER_56_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6626__3 clknet_1_1__leaf__2893_ vssd1 vssd1 vccd1 vccd1 net37 sky130_fd_sc_hd__inv_2
X_4035_ _0548_ egd_top.BitStream_buffer.BS_buffer\[28\] vssd1 vssd1 vccd1 vccd1 _0549_
+ sky130_fd_sc_hd__nand2_1
XFILLER_71_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5986_ _2464_ vssd1 vssd1 vccd1 vccd1 _2466_ sky130_fd_sc_hd__buf_2
X_4937_ _3202_ egd_top.BitStream_buffer.BS_buffer\[122\] vssd1 vssd1 vccd1 vccd1 _1445_
+ sky130_fd_sc_hd__nand2_1
X_4868_ _0605_ _0491_ vssd1 vssd1 vccd1 vccd1 _1376_ sky130_fd_sc_hd__nand2_1
X_3819_ _3338_ _3340_ _3341_ _0323_ _0332_ vssd1 vssd1 vccd1 vccd1 _0333_ sky130_fd_sc_hd__a221oi_1
X_4799_ _0527_ _0504_ _0531_ _0508_ _1307_ vssd1 vssd1 vccd1 vccd1 _1308_ sky130_fd_sc_hd__a221oi_1
XFILLER_21_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6469_ _2832_ vssd1 vssd1 vccd1 vccd1 _2833_ sky130_fd_sc_hd__inv_2
XFILLER_75_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_26 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6545__90 clknet_1_0__leaf__2885_ vssd1 vssd1 vccd1 vccd1 net124 sky130_fd_sc_hd__inv_2
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_83 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5840_ _3085_ _3329_ _2339_ vssd1 vssd1 vccd1 vccd1 _2340_ sky130_fd_sc_hd__o21ai_1
XFILLER_34_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5771_ _1076_ _3194_ _3197_ _0566_ _2271_ vssd1 vssd1 vccd1 vccd1 _2272_ sky130_fd_sc_hd__a221oi_1
X_4722_ _3126_ _3070_ vssd1 vssd1 vccd1 vccd1 _1231_ sky130_fd_sc_hd__nand2_1
XFILLER_14_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4653_ _3310_ _3322_ vssd1 vssd1 vccd1 vccd1 _1163_ sky130_fd_sc_hd__nand2_1
X_3604_ egd_top.BitStream_buffer.BS_buffer\[123\] vssd1 vssd1 vccd1 vccd1 _3138_ sky130_fd_sc_hd__buf_2
X_4584_ _0879_ _0402_ _1093_ vssd1 vssd1 vccd1 vccd1 _1094_ sky130_fd_sc_hd__o21ai_1
X_3535_ _3035_ _3068_ vssd1 vssd1 vccd1 vccd1 _3069_ sky130_fd_sc_hd__nor2_1
X_6323_ _2693_ vssd1 vssd1 vccd1 vccd1 _2694_ sky130_fd_sc_hd__inv_2
X_6254_ _2622_ _2623_ _2624_ vssd1 vssd1 vccd1 vccd1 _2625_ sky130_fd_sc_hd__and3_1
X_3466_ _2989_ _3006_ vssd1 vssd1 vccd1 vccd1 _3007_ sky130_fd_sc_hd__nand2_1
XFILLER_88_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5205_ _3127_ _3164_ vssd1 vssd1 vccd1 vccd1 _1710_ sky130_fd_sc_hd__nand2_1
XFILLER_69_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3397_ _2950_ vssd1 vssd1 vccd1 vccd1 _2951_ sky130_fd_sc_hd__inv_2
X_6185_ _2582_ _2583_ _2584_ vssd1 vssd1 vccd1 vccd1 _2585_ sky130_fd_sc_hd__a21bo_1
XFILLER_69_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5136_ _3100_ _3340_ _0714_ _0323_ _1641_ vssd1 vssd1 vccd1 vccd1 _1642_ sky130_fd_sc_hd__a221oi_1
X_6562__105 clknet_1_0__leaf__2887_ vssd1 vssd1 vccd1 vccd1 net139 sky130_fd_sc_hd__inv_2
XFILLER_29_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5067_ egd_top.BitStream_buffer.BS_buffer\[78\] vssd1 vssd1 vccd1 vccd1 _1574_ sky130_fd_sc_hd__inv_2
X_4018_ _0531_ vssd1 vssd1 vccd1 vccd1 _0532_ sky130_fd_sc_hd__inv_2
XFILLER_72_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5969_ _3005_ _2442_ _2446_ _2455_ vssd1 vssd1 vccd1 vccd1 _0270_ sky130_fd_sc_hd__o211a_1
XFILLER_52_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5823_ _3038_ _3075_ vssd1 vssd1 vccd1 vccd1 _2323_ sky130_fd_sc_hd__nand2_1
XFILLER_22_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_274 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5754_ _2983_ _3106_ _2252_ _2253_ _2254_ vssd1 vssd1 vccd1 vccd1 _2255_ sky130_fd_sc_hd__o2111a_1
XFILLER_22_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5685_ _0621_ egd_top.BitStream_buffer.BS_buffer\[12\] vssd1 vssd1 vccd1 vccd1 _2187_
+ sky130_fd_sc_hd__nand2_1
X_4705_ _3317_ _3299_ _1211_ _1212_ _1213_ vssd1 vssd1 vccd1 vccd1 _1214_ sky130_fd_sc_hd__o2111a_1
X_4636_ _3224_ egd_top.BitStream_buffer.BS_buffer\[74\] vssd1 vssd1 vccd1 vccd1 _1146_
+ sky130_fd_sc_hd__nand2_1
XFILLER_89_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4567_ _1002_ _1075_ _1077_ vssd1 vssd1 vccd1 vccd1 _1078_ sky130_fd_sc_hd__nand3_1
X_6306_ _2641_ _2667_ vssd1 vssd1 vccd1 vccd1 _2677_ sky130_fd_sc_hd__nor2_2
XFILLER_89_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3518_ _3051_ _3031_ _3032_ vssd1 vssd1 vccd1 vccd1 _3052_ sky130_fd_sc_hd__and3_2
X_4498_ _3294_ _3311_ vssd1 vssd1 vccd1 vccd1 _1009_ sky130_fd_sc_hd__nand2_1
X_3449_ _2989_ _2993_ vssd1 vssd1 vccd1 vccd1 _2994_ sky130_fd_sc_hd__nand2_1
X_6237_ _2608_ _3328_ vssd1 vssd1 vccd1 vccd1 _2615_ sky130_fd_sc_hd__nand2_1
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6168_ _3014_ _2555_ _2570_ _2571_ vssd1 vssd1 vccd1 vccd1 _0187_ sky130_fd_sc_hd__o211a_1
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5119_ _3268_ _3216_ _3272_ _3220_ _1624_ vssd1 vssd1 vccd1 vccd1 _1625_ sky130_fd_sc_hd__a221oi_1
XFILLER_84_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6099_ _2970_ _2940_ vssd1 vssd1 vccd1 vccd1 _2531_ sky130_fd_sc_hd__nand2_2
XFILLER_45_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f__2895_ clknet_0__2895_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__2895_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_48_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5470_ _2983_ _3089_ _1970_ _1971_ _1972_ vssd1 vssd1 vccd1 vccd1 _1973_ sky130_fd_sc_hd__o2111a_1
XFILLER_8_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4421_ egd_top.BitStream_buffer.BitStream_buffer_output\[13\] vssd1 vssd1 vccd1 vccd1
+ _0933_ sky130_fd_sc_hd__inv_2
X_4352_ _0354_ _0342_ _0345_ _0347_ _0863_ vssd1 vssd1 vccd1 vccd1 _0864_ sky130_fd_sc_hd__a221oi_1
XTAP_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4283_ _0628_ _0795_ vssd1 vssd1 vccd1 vccd1 _0296_ sky130_fd_sc_hd__nor2_1
XFILLER_86_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6022_ _2485_ vssd1 vssd1 vccd1 vccd1 _2486_ sky130_fd_sc_hd__clkbuf_2
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6855_ net99 _0314_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BitStream_buffer_valid_n
+ sky130_fd_sc_hd__dfxtp_1
X_3998_ _0511_ vssd1 vssd1 vccd1 vccd1 _0512_ sky130_fd_sc_hd__clkbuf_4
X_5806_ _2248_ _2305_ _2306_ vssd1 vssd1 vccd1 vccd1 _2307_ sky130_fd_sc_hd__nand3_1
XFILLER_13_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6786_ net190 _0245_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[34\]
+ sky130_fd_sc_hd__dfxtp_4
X_5737_ _0513_ _0364_ vssd1 vssd1 vccd1 vccd1 _2238_ sky130_fd_sc_hd__nand2_1
XFILLER_13_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5668_ _2159_ _2163_ _2166_ _2169_ vssd1 vssd1 vccd1 vccd1 _2170_ sky130_fd_sc_hd__and4_1
X_4619_ _0496_ _0509_ vssd1 vssd1 vccd1 vccd1 _1129_ sky130_fd_sc_hd__nand2_1
X_5599_ _0560_ _0491_ vssd1 vssd1 vccd1 vccd1 _2101_ sky130_fd_sc_hd__nand2_1
XFILLER_89_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6568__111 clknet_1_0__leaf__2887_ vssd1 vssd1 vccd1 vccd1 net145 sky130_fd_sc_hd__inv_2
XFILLER_1_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_54 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4970_ _0653_ _0403_ _1476_ vssd1 vssd1 vccd1 vccd1 _1477_ sky130_fd_sc_hd__o21ai_1
X_3921_ _0434_ vssd1 vssd1 vccd1 vccd1 _0435_ sky130_fd_sc_hd__buf_6
XFILLER_32_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3852_ _0365_ vssd1 vssd1 vccd1 vccd1 _0366_ sky130_fd_sc_hd__inv_2
X_5522_ _0448_ _0425_ vssd1 vssd1 vccd1 vccd1 _2025_ sky130_fd_sc_hd__or2_1
X_3783_ egd_top.BitStream_buffer.BS_buffer\[85\] vssd1 vssd1 vccd1 vccd1 _3317_ sky130_fd_sc_hd__clkinv_2
X_5453_ _3309_ _3040_ vssd1 vssd1 vccd1 vccd1 _1956_ sky130_fd_sc_hd__nand2_1
X_4404_ _0578_ _0583_ vssd1 vssd1 vccd1 vccd1 _0916_ sky130_fd_sc_hd__nand2_1
X_5384_ _0708_ _3333_ _1886_ _1887_ vssd1 vssd1 vccd1 vccd1 _1888_ sky130_fd_sc_hd__a211oi_1
XFILLER_5_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4335_ _3314_ _3311_ vssd1 vssd1 vccd1 vccd1 _0847_ sky130_fd_sc_hd__nand2_1
XFILLER_59_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4266_ egd_top.BitStream_buffer.BS_buffer\[90\] vssd1 vssd1 vccd1 vccd1 _0779_ sky130_fd_sc_hd__clkinv_2
X_4197_ _3061_ _3094_ vssd1 vssd1 vccd1 vccd1 _0710_ sky130_fd_sc_hd__nand2_1
XFILLER_39_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6005_ _2471_ _0520_ vssd1 vssd1 vccd1 vccd1 _2477_ sky130_fd_sc_hd__nand2_1
XFILLER_42_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6838_ net82 _0297_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BitStream_buffer_output\[15\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__2897_ _2897_ vssd1 vssd1 vccd1 vccd1 clknet_0__2897_ sky130_fd_sc_hd__clkbuf_16
XFILLER_10_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6769_ net173 _0228_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[51\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_2_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6622__160 clknet_1_1__leaf__2892_ vssd1 vssd1 vccd1 vccd1 net194 sky130_fd_sc_hd__inv_2
XFILLER_5_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4120_ egd_top.BitStream_buffer.BS_buffer\[34\] vssd1 vssd1 vccd1 vccd1 _0633_ sky130_fd_sc_hd__inv_2
X_4051_ _0564_ vssd1 vssd1 vccd1 vccd1 _0565_ sky130_fd_sc_hd__buf_2
XFILLER_1_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput5 la_data_in_58_43[13] vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4953_ _1447_ _1452_ _1457_ _1460_ vssd1 vssd1 vccd1 vccd1 _1461_ sky130_fd_sc_hd__and4_1
XFILLER_51_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3904_ _0417_ vssd1 vssd1 vccd1 vccd1 _0418_ sky130_fd_sc_hd__clkbuf_2
XFILLER_51_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4884_ _0702_ _0522_ _0366_ _0525_ _1391_ vssd1 vssd1 vccd1 vccd1 _1392_ sky130_fd_sc_hd__o221a_1
XFILLER_20_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3835_ _3087_ _0339_ vssd1 vssd1 vccd1 vccd1 _0349_ sky130_fd_sc_hd__nand2_1
X_3766_ _3290_ _3046_ vssd1 vssd1 vccd1 vccd1 _3300_ sky130_fd_sc_hd__nor2_2
X_5505_ _0586_ _3183_ _2007_ vssd1 vssd1 vccd1 vccd1 _2008_ sky130_fd_sc_hd__o21ai_1
X_6485_ _2837_ _2847_ vssd1 vssd1 vccd1 vccd1 _2848_ sky130_fd_sc_hd__nand2_1
X_5436_ _1930_ _1934_ _1936_ _1939_ vssd1 vssd1 vccd1 vccd1 _1940_ sky130_fd_sc_hd__and4_1
X_3697_ _3052_ _3213_ vssd1 vssd1 vccd1 vccd1 _3231_ sky130_fd_sc_hd__and2_1
XFILLER_10_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5367_ _0602_ _0571_ vssd1 vssd1 vccd1 vccd1 _1871_ sky130_fd_sc_hd__or2_1
X_5298_ egd_top.BitStream_buffer.BS_buffer\[29\] _0504_ _0537_ _0508_ _1802_ vssd1
+ vssd1 vccd1 vccd1 _1803_ sky130_fd_sc_hd__a221oi_1
XFILLER_87_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4318_ _3243_ _3230_ vssd1 vssd1 vccd1 vccd1 _0830_ sky130_fd_sc_hd__nand2_1
XFILLER_59_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4249_ _3252_ _3251_ _3268_ _3255_ _0761_ vssd1 vssd1 vccd1 vccd1 _0762_ sky130_fd_sc_hd__a221oi_1
XFILLER_19_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3620_ _3052_ _3142_ vssd1 vssd1 vccd1 vccd1 _3154_ sky130_fd_sc_hd__and2_1
X_3551_ egd_top.BitStream_buffer.BS_buffer\[103\] vssd1 vssd1 vccd1 vccd1 _3085_ sky130_fd_sc_hd__clkinv_2
X_6270_ _2638_ _2640_ vssd1 vssd1 vccd1 vccd1 _2641_ sky130_fd_sc_hd__nand2_1
X_3482_ _2989_ _3018_ vssd1 vssd1 vccd1 vccd1 _3019_ sky130_fd_sc_hd__nand2_1
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5221_ _3309_ _3341_ vssd1 vssd1 vccd1 vccd1 _1726_ sky130_fd_sc_hd__nand2_1
X_5152_ _1648_ _1651_ _1654_ _1657_ vssd1 vssd1 vccd1 vccd1 _1658_ sky130_fd_sc_hd__and4_1
X_4103_ _0552_ _0616_ vssd1 vssd1 vccd1 vccd1 _0617_ sky130_fd_sc_hd__nand2_1
X_5083_ _0721_ _3056_ _1588_ vssd1 vssd1 vccd1 vccd1 _1589_ sky130_fd_sc_hd__o21ai_1
XFILLER_56_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4034_ _0547_ vssd1 vssd1 vccd1 vccd1 _0548_ sky130_fd_sc_hd__buf_4
XFILLER_64_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5985_ _2464_ vssd1 vssd1 vccd1 vccd1 _2465_ sky130_fd_sc_hd__buf_2
X_4936_ _3193_ egd_top.BitStream_buffer.BS_buffer\[124\] vssd1 vssd1 vccd1 vccd1 _1444_
+ sky130_fd_sc_hd__nand2_1
X_4867_ _0608_ _0502_ vssd1 vssd1 vccd1 vccd1 _1375_ sky130_fd_sc_hd__nand2_1
XANTENNA_10 _2303_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3818_ _0324_ _0327_ _0331_ vssd1 vssd1 vccd1 vccd1 _0332_ sky130_fd_sc_hd__o21ai_1
X_4798_ _0699_ _0512_ _1306_ vssd1 vssd1 vccd1 vccd1 _1307_ sky130_fd_sc_hd__o21ai_1
XFILLER_21_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3749_ egd_top.BitStream_buffer.BS_buffer\[78\] vssd1 vssd1 vccd1 vccd1 _3283_ sky130_fd_sc_hd__clkbuf_4
X_6468_ _2923_ _2699_ _2693_ vssd1 vssd1 vccd1 vccd1 _2832_ sky130_fd_sc_hd__or3_2
X_5419_ _2980_ _3089_ _1920_ _1921_ _1922_ vssd1 vssd1 vccd1 vccd1 _1923_ sky130_fd_sc_hd__o2111a_1
X_6399_ net17 _2700_ _2739_ _2768_ vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__a31o_2
XFILLER_87_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5770_ _0591_ _3200_ _2270_ vssd1 vssd1 vccd1 vccd1 _2271_ sky130_fd_sc_hd__o21ai_1
XFILLER_34_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4721_ _0721_ _3106_ _1227_ _1228_ _1229_ vssd1 vssd1 vccd1 vccd1 _1230_ sky130_fd_sc_hd__o2111a_1
X_4652_ _3314_ _3334_ vssd1 vssd1 vccd1 vccd1 _1162_ sky130_fd_sc_hd__nand2_1
X_3603_ _3136_ vssd1 vssd1 vccd1 vccd1 _3137_ sky130_fd_sc_hd__buf_4
X_4583_ _0405_ _0412_ vssd1 vssd1 vccd1 vccd1 _1093_ sky130_fd_sc_hd__nand2_1
X_3534_ _3067_ vssd1 vssd1 vccd1 vccd1 _3068_ sky130_fd_sc_hd__clkinv_2
X_6322_ _2691_ _2692_ vssd1 vssd1 vccd1 vccd1 _2693_ sky130_fd_sc_hd__nand2_1
X_6253_ egd_top.BitStream_buffer.BitStream_buffer_output\[14\] vssd1 vssd1 vccd1 vccd1
+ _2624_ sky130_fd_sc_hd__clkinv_2
X_3465_ egd_top.BitStream_buffer.BS_buffer\[121\] vssd1 vssd1 vccd1 vccd1 _3006_ sky130_fd_sc_hd__clkinv_2
X_5204_ _0746_ _3069_ _3191_ _3074_ _1708_ vssd1 vssd1 vccd1 vccd1 _1709_ sky130_fd_sc_hd__a221oi_1
X_3396_ _2948_ _2949_ vssd1 vssd1 vccd1 vccd1 _2950_ sky130_fd_sc_hd__nand2_1
X_6184_ egd_top.BitStream_buffer.pc_previous\[3\] egd_top.BitStream_buffer.exp_golomb_len\[3\]
+ vssd1 vssd1 vccd1 vccd1 _2584_ sky130_fd_sc_hd__nand2_1
X_5135_ _3102_ _0327_ _1640_ vssd1 vssd1 vccd1 vccd1 _1641_ sky130_fd_sc_hd__o21ai_1
X_5066_ _3264_ _3233_ _3236_ _3248_ _1572_ vssd1 vssd1 vccd1 vccd1 _1573_ sky130_fd_sc_hd__a221oi_2
XFILLER_84_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4017_ egd_top.BitStream_buffer.BS_buffer\[26\] vssd1 vssd1 vccd1 vccd1 _0531_ sky130_fd_sc_hd__clkbuf_4
XFILLER_37_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5968_ _2449_ _0586_ vssd1 vssd1 vccd1 vccd1 _2455_ sky130_fd_sc_hd__nand2_1
X_4919_ _3223_ egd_top.BitStream_buffer.BS_buffer\[76\] vssd1 vssd1 vccd1 vccd1 _1427_
+ sky130_fd_sc_hd__nand2_1
X_5899_ _2388_ _2391_ _2395_ _2398_ vssd1 vssd1 vccd1 vccd1 _2399_ sky130_fd_sc_hd__and4_1
XFILLER_32_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_507 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5822_ _2312_ _2315_ _2317_ _2321_ vssd1 vssd1 vccd1 vccd1 _2322_ sky130_fd_sc_hd__and4_1
XFILLER_34_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5753_ _2990_ _3088_ vssd1 vssd1 vccd1 vccd1 _2254_ sky130_fd_sc_hd__or2_1
XFILLER_34_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4704_ _3301_ _3311_ vssd1 vssd1 vccd1 vccd1 _1213_ sky130_fd_sc_hd__nand2_1
X_5684_ _2157_ _2185_ vssd1 vssd1 vccd1 vccd1 _2186_ sky130_fd_sc_hd__nor2_1
XFILLER_30_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4635_ _3225_ vssd1 vssd1 vccd1 vccd1 _1145_ sky130_fd_sc_hd__clkbuf_4
X_4566_ _0622_ _1076_ vssd1 vssd1 vccd1 vccd1 _1077_ sky130_fd_sc_hd__nand2_1
X_3517_ _3050_ vssd1 vssd1 vccd1 vccd1 _3051_ sky130_fd_sc_hd__inv_2
X_6305_ _2672_ _2675_ vssd1 vssd1 vccd1 vccd1 _2676_ sky130_fd_sc_hd__nor2b_1
X_4497_ _3291_ _0774_ vssd1 vssd1 vccd1 vccd1 _1008_ sky130_fd_sc_hd__nand2_1
X_6685__57 clknet_1_0__leaf__2898_ vssd1 vssd1 vccd1 vccd1 net91 sky130_fd_sc_hd__inv_2
X_3448_ egd_top.BitStream_buffer.BS_buffer\[117\] vssd1 vssd1 vccd1 vccd1 _2993_ sky130_fd_sc_hd__clkinv_2
X_6236_ _3001_ _2602_ _2611_ _2614_ vssd1 vssd1 vccd1 vccd1 _0168_ sky130_fd_sc_hd__o211a_1
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6167_ _2561_ _1025_ vssd1 vssd1 vccd1 vccd1 _2571_ sky130_fd_sc_hd__nand2_1
X_3379_ _2932_ egd_top.BitStream_buffer.pc\[4\] egd_top.BitStream_buffer.pc\[5\] vssd1
+ vssd1 vccd1 vccd1 _2933_ sky130_fd_sc_hd__and3_2
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5118_ _3277_ _1145_ _1623_ vssd1 vssd1 vccd1 vccd1 _1624_ sky130_fd_sc_hd__o21ai_1
XFILLER_84_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6098_ _3023_ _2511_ _2528_ _2530_ vssd1 vssd1 vccd1 vccd1 _0216_ sky130_fd_sc_hd__o211a_1
XFILLER_84_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5049_ _3310_ _0785_ vssd1 vssd1 vccd1 vccd1 _1556_ sky130_fd_sc_hd__nand2_1
XFILLER_43_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1__f__2894_ clknet_0__2894_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__2894_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_68_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4420_ _0860_ _0929_ _0931_ vssd1 vssd1 vccd1 vccd1 _0932_ sky130_fd_sc_hd__nand3_1
X_4351_ _0861_ _0350_ _0862_ vssd1 vssd1 vccd1 vccd1 _0863_ sky130_fd_sc_hd__o21ai_1
XTAP_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4282_ _3027_ _0794_ vssd1 vssd1 vccd1 vccd1 _0795_ sky130_fd_sc_hd__nor2_1
XFILLER_58_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6021_ egd_top.BitStream_buffer.buffer_index\[6\] _2938_ egd_top.BitStream_buffer.buffer_index\[4\]
+ _2437_ vssd1 vssd1 vccd1 vccd1 _2485_ sky130_fd_sc_hd__or4_1
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6854_ net98 _0313_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[112\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_50_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3997_ _3087_ _0484_ vssd1 vssd1 vccd1 vccd1 _0511_ sky130_fd_sc_hd__nand2_1
X_5805_ _0621_ egd_top.BitStream_buffer.BS_buffer\[13\] vssd1 vssd1 vccd1 vccd1 _2306_
+ sky130_fd_sc_hd__nand2_1
XFILLER_10_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6785_ net189 _0244_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[35\]
+ sky130_fd_sc_hd__dfxtp_1
X_5736_ _0907_ _0494_ _2234_ _2235_ _2236_ vssd1 vssd1 vccd1 vccd1 _2237_ sky130_fd_sc_hd__o2111a_1
X_5667_ _0579_ _3176_ _0585_ _3180_ _2168_ vssd1 vssd1 vccd1 vccd1 _2169_ sky130_fd_sc_hd__a221oi_1
X_4618_ egd_top.BitStream_buffer.BS_buffer\[22\] vssd1 vssd1 vccd1 vccd1 _1128_ sky130_fd_sc_hd__clkinv_2
X_5598_ _2088_ _2092_ _2096_ _2099_ vssd1 vssd1 vccd1 vccd1 _2100_ sky130_fd_sc_hd__and4_1
X_4549_ _3003_ _3199_ _1057_ _1058_ _1059_ vssd1 vssd1 vccd1 vccd1 _1060_ sky130_fd_sc_hd__o2111a_1
XFILLER_1_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6219_ _2603_ _0767_ vssd1 vssd1 vccd1 vccd1 _2605_ sky130_fd_sc_hd__nand2_1
XFILLER_85_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_186 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6649__24 clknet_1_0__leaf__2895_ vssd1 vssd1 vccd1 vccd1 net58 sky130_fd_sc_hd__inv_2
XFILLER_79_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6664__38 clknet_1_0__leaf__2896_ vssd1 vssd1 vccd1 vccd1 net72 sky130_fd_sc_hd__inv_2
XFILLER_91_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_476 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3920_ _0433_ vssd1 vssd1 vccd1 vccd1 _0434_ sky130_fd_sc_hd__buf_6
XFILLER_63_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3851_ egd_top.BitStream_buffer.BS_buffer\[33\] vssd1 vssd1 vccd1 vccd1 _0365_ sky130_fd_sc_hd__clkbuf_4
XFILLER_81_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3782_ _3314_ _3315_ vssd1 vssd1 vccd1 vccd1 _3316_ sky130_fd_sc_hd__nand2_1
X_5521_ _2014_ _2017_ _2020_ _2023_ vssd1 vssd1 vccd1 vccd1 _2024_ sky130_fd_sc_hd__and4_1
XFILLER_8_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5452_ _3313_ _3341_ vssd1 vssd1 vccd1 vccd1 _1955_ sky130_fd_sc_hd__nand2_1
X_4403_ _0586_ _0558_ _0912_ _0913_ _0914_ vssd1 vssd1 vccd1 vccd1 _0915_ sky130_fd_sc_hd__o2111a_1
X_5383_ _3094_ _3323_ _3325_ _0716_ vssd1 vssd1 vccd1 vccd1 _1887_ sky130_fd_sc_hd__a22o_1
XFILLER_5_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4334_ _3310_ _3334_ vssd1 vssd1 vccd1 vccd1 _0846_ sky130_fd_sc_hd__nand2_1
X_6004_ _2998_ _2465_ _2474_ _2476_ vssd1 vssd1 vccd1 vccd1 _0256_ sky130_fd_sc_hd__o211a_1
X_4265_ _0771_ _3319_ _0773_ _0775_ _0777_ vssd1 vssd1 vccd1 vccd1 _0778_ sky130_fd_sc_hd__o2111a_1
X_4196_ egd_top.BitStream_buffer.BS_buffer\[99\] vssd1 vssd1 vccd1 vccd1 _0709_ sky130_fd_sc_hd__clkinv_2
XFILLER_67_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_359 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6598__138 clknet_1_0__leaf__2890_ vssd1 vssd1 vccd1 vccd1 net172 sky130_fd_sc_hd__inv_2
XFILLER_23_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_0__2896_ _2896_ vssd1 vssd1 vccd1 vccd1 clknet_0__2896_ sky130_fd_sc_hd__clkbuf_16
X_6837_ net81 _0296_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BitStream_buffer_output\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_24_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6768_ net172 _0227_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[52\]
+ sky130_fd_sc_hd__dfxtp_1
X_5719_ _0564_ egd_top.BitStream_buffer.BS_buffer\[17\] vssd1 vssd1 vccd1 vccd1 _2220_
+ sky130_fd_sc_hd__nand2_1
XFILLER_2_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4050_ _0559_ _3091_ vssd1 vssd1 vccd1 vccd1 _0564_ sky130_fd_sc_hd__nor2_2
XFILLER_68_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput6 la_data_in_58_43[14] vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__clkbuf_1
XFILLER_64_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4952_ _0930_ _3175_ _1076_ _3179_ _1459_ vssd1 vssd1 vccd1 vccd1 _1460_ sky130_fd_sc_hd__a221oi_1
X_4883_ _0907_ _0529_ _0995_ _0533_ vssd1 vssd1 vccd1 vccd1 _1391_ sky130_fd_sc_hd__o22a_1
X_3903_ _3058_ _2933_ vssd1 vssd1 vccd1 vccd1 _0417_ sky130_fd_sc_hd__and2_1
X_3834_ _0347_ vssd1 vssd1 vccd1 vccd1 _0348_ sky130_fd_sc_hd__inv_2
XFILLER_32_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3765_ _3298_ vssd1 vssd1 vccd1 vccd1 _3299_ sky130_fd_sc_hd__clkbuf_4
X_5504_ _3175_ _0553_ vssd1 vssd1 vccd1 vccd1 _2007_ sky130_fd_sc_hd__nand2_1
X_6484_ _2846_ _2684_ vssd1 vssd1 vccd1 vccd1 _2847_ sky130_fd_sc_hd__nand2_1
X_3696_ egd_top.BitStream_buffer.BS_buffer\[66\] vssd1 vssd1 vccd1 vccd1 _3230_ sky130_fd_sc_hd__clkbuf_4
X_5435_ _0623_ _3194_ _3197_ _0792_ _1938_ vssd1 vssd1 vccd1 vccd1 _1939_ sky130_fd_sc_hd__a221oi_1
X_5366_ _0561_ egd_top.BitStream_buffer.BS_buffer\[16\] vssd1 vssd1 vccd1 vccd1 _1870_
+ sky130_fd_sc_hd__nand2_1
XFILLER_59_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5297_ _0995_ _0512_ _1801_ vssd1 vssd1 vccd1 vccd1 _1802_ sky130_fd_sc_hd__o21ai_1
X_4317_ egd_top.BitStream_buffer.BS_buffer\[67\] vssd1 vssd1 vccd1 vccd1 _0829_ sky130_fd_sc_hd__clkinv_2
XFILLER_19_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4248_ _0759_ _3260_ _0760_ vssd1 vssd1 vccd1 vccd1 _0761_ sky130_fd_sc_hd__o21ai_1
XFILLER_74_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6643__19 clknet_1_0__leaf__2894_ vssd1 vssd1 vccd1 vccd1 net53 sky130_fd_sc_hd__inv_2
X_4179_ _0498_ vssd1 vssd1 vccd1 vccd1 _0692_ sky130_fd_sc_hd__inv_2
XFILLER_67_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6606__145 clknet_1_1__leaf__2891_ vssd1 vssd1 vccd1 vccd1 net179 sky130_fd_sc_hd__inv_2
XFILLER_55_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3550_ _3066_ _3069_ _3070_ _3074_ _3083_ vssd1 vssd1 vccd1 vccd1 _3084_ sky130_fd_sc_hd__a221oi_1
X_3481_ egd_top.BitStream_buffer.BS_buffer\[125\] vssd1 vssd1 vccd1 vccd1 _3018_ sky130_fd_sc_hd__clkinv_2
X_5220_ _3328_ _3298_ _1722_ _1723_ _1724_ vssd1 vssd1 vccd1 vccd1 _1725_ sky130_fd_sc_hd__o2111a_1
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5151_ _0443_ _0396_ _0399_ _0655_ _1656_ vssd1 vssd1 vccd1 vccd1 _1657_ sky130_fd_sc_hd__a221oi_1
X_4102_ _0573_ _0590_ _0601_ _0615_ vssd1 vssd1 vccd1 vccd1 _0616_ sky130_fd_sc_hd__and4_1
X_5082_ _3061_ _3118_ vssd1 vssd1 vccd1 vccd1 _1588_ sky130_fd_sc_hd__nand2_1
XFILLER_84_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4033_ _0488_ _3068_ vssd1 vssd1 vccd1 vccd1 _0547_ sky130_fd_sc_hd__nor2_2
XFILLER_49_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5984_ _2463_ vssd1 vssd1 vccd1 vccd1 _2464_ sky130_fd_sc_hd__clkbuf_2
X_4935_ _1429_ _1434_ _1439_ _1442_ vssd1 vssd1 vccd1 vccd1 _1443_ sky130_fd_sc_hd__and4_1
X_4866_ _0670_ _0592_ _0554_ _0596_ _1373_ vssd1 vssd1 vccd1 vccd1 _1374_ sky130_fd_sc_hd__o221a_1
XANTENNA_11 _2992_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4797_ _0514_ egd_top.BitStream_buffer.BS_buffer\[27\] vssd1 vssd1 vccd1 vccd1 _1306_
+ sky130_fd_sc_hd__nand2_1
XFILLER_20_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3817_ _0329_ _0330_ vssd1 vssd1 vccd1 vccd1 _0331_ sky130_fd_sc_hd__nand2_1
X_3748_ _3281_ vssd1 vssd1 vccd1 vccd1 _3282_ sky130_fd_sc_hd__clkbuf_4
X_6536_ clknet_1_0__leaf__2883_ vssd1 vssd1 vccd1 vccd1 _2885_ sky130_fd_sc_hd__buf_1
X_3679_ _3212_ vssd1 vssd1 vccd1 vccd1 _3213_ sky130_fd_sc_hd__buf_2
X_6467_ _2822_ _2830_ vssd1 vssd1 vccd1 vccd1 _2831_ sky130_fd_sc_hd__nand2_1
X_5418_ _1035_ _3106_ vssd1 vssd1 vccd1 vccd1 _1922_ sky130_fd_sc_hd__or2_1
X_6398_ _2765_ _2767_ _2736_ vssd1 vssd1 vccd1 vccd1 _2768_ sky130_fd_sc_hd__and3_1
X_5349_ _0477_ _3256_ vssd1 vssd1 vccd1 vccd1 _1853_ sky130_fd_sc_hd__nand2_1
XFILLER_87_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4720_ _1025_ _3088_ vssd1 vssd1 vccd1 vccd1 _1229_ sky130_fd_sc_hd__or2_1
X_4651_ _3311_ _3292_ _0772_ _3295_ _1160_ vssd1 vssd1 vccd1 vccd1 _1161_ sky130_fd_sc_hd__a221oi_1
X_3602_ _3135_ vssd1 vssd1 vccd1 vccd1 _3136_ sky130_fd_sc_hd__clkbuf_2
X_4582_ _0401_ _0384_ _1089_ _1090_ _1091_ vssd1 vssd1 vccd1 vccd1 _1092_ sky130_fd_sc_hd__o2111a_1
X_3533_ _2920_ _3029_ vssd1 vssd1 vccd1 vccd1 _3067_ sky130_fd_sc_hd__nor2_4
X_6321_ _2636_ _2640_ vssd1 vssd1 vccd1 vccd1 _2692_ sky130_fd_sc_hd__nand2_1
X_3464_ net13 vssd1 vssd1 vccd1 vccd1 _3005_ sky130_fd_sc_hd__clkbuf_4
X_6551__95 clknet_1_1__leaf__2886_ vssd1 vssd1 vccd1 vccd1 net129 sky130_fd_sc_hd__inv_2
X_6252_ egd_top.BitStream_buffer.BitStream_buffer_valid_n egd_top.BitStream_buffer.BitStream_buffer_output\[15\]
+ vssd1 vssd1 vccd1 vccd1 _2623_ sky130_fd_sc_hd__nor2_4
XFILLER_88_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_310 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5203_ egd_top.BitStream_buffer.BS_buffer\[119\] _3078_ _3080_ egd_top.BitStream_buffer.BS_buffer\[120\]
+ vssd1 vssd1 vccd1 vccd1 _1708_ sky130_fd_sc_hd__a22o_1
X_6183_ egd_top.BitStream_buffer.pc_previous\[3\] egd_top.BitStream_buffer.exp_golomb_len\[3\]
+ vssd1 vssd1 vccd1 vccd1 _2583_ sky130_fd_sc_hd__or2_1
X_5134_ _0329_ _3094_ vssd1 vssd1 vccd1 vccd1 _1640_ sky130_fd_sc_hd__nand2_1
X_3395_ _2908_ _2906_ net34 net32 vssd1 vssd1 vccd1 vccd1 _2949_ sky130_fd_sc_hd__and4_1
XFILLER_57_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5065_ _3257_ _3240_ _1571_ vssd1 vssd1 vccd1 vccd1 _1572_ sky130_fd_sc_hd__o21ai_1
X_4016_ _0529_ vssd1 vssd1 vccd1 vccd1 _0530_ sky130_fd_sc_hd__buf_2
XFILLER_80_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5967_ _3001_ _2442_ _2446_ _2454_ vssd1 vssd1 vccd1 vccd1 _0271_ sky130_fd_sc_hd__o211a_1
X_4918_ egd_top.BitStream_buffer.BS_buffer\[77\] vssd1 vssd1 vccd1 vccd1 _1426_ sky130_fd_sc_hd__clkinv_2
XFILLER_40_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5898_ _3248_ _0470_ _3252_ _0473_ _2397_ vssd1 vssd1 vccd1 vccd1 _2398_ sky130_fd_sc_hd__a221oi_1
XFILLER_32_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4849_ _0432_ _0467_ vssd1 vssd1 vccd1 vccd1 _1357_ sky130_fd_sc_hd__nand2_1
X_6519_ _2865_ _2879_ vssd1 vssd1 vccd1 vccd1 _2880_ sky130_fd_sc_hd__nand2_1
XFILLER_0_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5821_ _0771_ _3260_ _2318_ _2319_ _2320_ vssd1 vssd1 vccd1 vccd1 _2321_ sky130_fd_sc_hd__o2111a_1
X_5752_ _3093_ _3164_ vssd1 vssd1 vccd1 vccd1 _2253_ sky130_fd_sc_hd__nand2_1
X_4703_ _3294_ _3334_ vssd1 vssd1 vccd1 vccd1 _1212_ sky130_fd_sc_hd__nand2_1
X_5683_ _2170_ _2184_ vssd1 vssd1 vccd1 vccd1 _2185_ sky130_fd_sc_hd__nand2_1
XFILLER_30_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4634_ egd_top.BitStream_buffer.BS_buffer\[75\] vssd1 vssd1 vccd1 vccd1 _1144_ sky130_fd_sc_hd__clkinv_2
X_4565_ egd_top.BitStream_buffer.BS_buffer\[3\] vssd1 vssd1 vccd1 vccd1 _1076_ sky130_fd_sc_hd__clkbuf_4
X_3516_ _2929_ egd_top.BitStream_buffer.pc\[1\] vssd1 vssd1 vccd1 vccd1 _3050_ sky130_fd_sc_hd__nand2_1
X_6304_ egd_top.BitStream_buffer.BitStream_buffer_output\[5\] _2673_ _2674_ vssd1
+ vssd1 vccd1 vccd1 _2675_ sky130_fd_sc_hd__o21a_1
X_4496_ egd_top.BitStream_buffer.BS_buffer\[83\] vssd1 vssd1 vccd1 vccd1 _1007_ sky130_fd_sc_hd__clkinv_2
XFILLER_89_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3447_ net2 vssd1 vssd1 vccd1 vccd1 _2992_ sky130_fd_sc_hd__buf_4
X_6235_ _2608_ _0776_ vssd1 vssd1 vccd1 vccd1 _2614_ sky130_fd_sc_hd__nand2_1
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3378_ egd_top.BitStream_buffer.pc\[6\] vssd1 vssd1 vccd1 vccd1 _2932_ sky130_fd_sc_hd__clkinv_2
X_6166_ _2904_ vssd1 vssd1 vccd1 vccd1 _2570_ sky130_fd_sc_hd__buf_2
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_195 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6097_ _2509_ _0474_ vssd1 vssd1 vccd1 vccd1 _2530_ sky130_fd_sc_hd__nand2_1
X_5117_ _3224_ _3283_ vssd1 vssd1 vccd1 vccd1 _1623_ sky130_fd_sc_hd__nand2_1
X_5048_ _3314_ _3327_ vssd1 vssd1 vccd1 vccd1 _1555_ sky130_fd_sc_hd__nand2_1
XFILLER_72_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6530__76 clknet_1_0__leaf__2884_ vssd1 vssd1 vccd1 vccd1 net110 sky130_fd_sc_hd__inv_2
XFILLER_0_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1__f__2893_ clknet_0__2893_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__2893_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_88_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4350_ _0353_ _0375_ vssd1 vssd1 vccd1 vccd1 _0862_ sky130_fd_sc_hd__nand2_1
X_4281_ _0707_ _0791_ _0793_ vssd1 vssd1 vccd1 vccd1 _0794_ sky130_fd_sc_hd__nand3_1
XTAP_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6020_ _3023_ _2466_ _2474_ _2484_ vssd1 vssd1 vccd1 vccd1 _0248_ sky130_fd_sc_hd__o211a_1
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6853_ net97 _0312_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[113\]
+ sky130_fd_sc_hd__dfxtp_2
X_5804_ _2277_ _2304_ vssd1 vssd1 vccd1 vccd1 _2305_ sky130_fd_sc_hd__nor2_1
XFILLER_62_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3996_ _0509_ vssd1 vssd1 vccd1 vccd1 _0510_ sky130_fd_sc_hd__inv_2
X_6784_ net188 _0243_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[36\]
+ sky130_fd_sc_hd__dfxtp_1
X_5735_ _0496_ egd_top.BitStream_buffer.BS_buffer\[32\] vssd1 vssd1 vccd1 vccd1 _2236_
+ sky130_fd_sc_hd__nand2_1
X_5666_ _0679_ _3183_ _2167_ vssd1 vssd1 vccd1 vccd1 _2168_ sky130_fd_sc_hd__o21ai_1
XFILLER_30_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4617_ _1116_ _1120_ _1122_ _1126_ vssd1 vssd1 vccd1 vccd1 _1127_ sky130_fd_sc_hd__and4_1
X_5597_ _3256_ _0470_ _3264_ _0473_ _2098_ vssd1 vssd1 vccd1 vccd1 _2099_ sky130_fd_sc_hd__a221oi_1
X_4548_ _3196_ egd_top.BitStream_buffer.BS_buffer\[122\] vssd1 vssd1 vccd1 vccd1 _1059_
+ sky130_fd_sc_hd__nand2_1
X_4479_ _0986_ _0494_ _0987_ _0988_ _0989_ vssd1 vssd1 vccd1 vccd1 _0990_ sky130_fd_sc_hd__o2111a_1
XFILLER_77_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6218_ _2966_ _2602_ _2570_ _2604_ vssd1 vssd1 vccd1 vccd1 _0176_ sky130_fd_sc_hd__o211a_1
XFILLER_57_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6149_ _2553_ vssd1 vssd1 vccd1 vccd1 _2561_ sky130_fd_sc_hd__buf_2
XFILLER_57_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_198 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6575__117 clknet_1_1__leaf__2888_ vssd1 vssd1 vccd1 vccd1 net151 sky130_fd_sc_hd__inv_2
XFILLER_5_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3850_ egd_top.BitStream_buffer.BS_buffer\[35\] vssd1 vssd1 vccd1 vccd1 _0364_ sky130_fd_sc_hd__clkbuf_4
X_3781_ egd_top.BitStream_buffer.BS_buffer\[84\] vssd1 vssd1 vccd1 vccd1 _3315_ sky130_fd_sc_hd__clkbuf_4
XFILLER_74_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5520_ _0436_ _0396_ _0399_ _0454_ _2022_ vssd1 vssd1 vccd1 vccd1 _2023_ sky130_fd_sc_hd__a221oi_1
X_5451_ _0850_ _3298_ _1951_ _1952_ _1953_ vssd1 vssd1 vccd1 vccd1 _1954_ sky130_fd_sc_hd__o2111a_1
X_4402_ _0554_ _0571_ vssd1 vssd1 vccd1 vccd1 _0914_ sky130_fd_sc_hd__or2_1
X_5382_ _0709_ _3330_ vssd1 vssd1 vccd1 vccd1 _1886_ sky130_fd_sc_hd__nor2_1
X_4333_ _3315_ _3292_ _0774_ _3295_ _0844_ vssd1 vssd1 vccd1 vccd1 _0845_ sky130_fd_sc_hd__a221oi_1
X_4264_ _0776_ _3307_ vssd1 vssd1 vccd1 vccd1 _0777_ sky130_fd_sc_hd__or2_1
XFILLER_86_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6003_ _2471_ _0510_ vssd1 vssd1 vccd1 vccd1 _2476_ sky130_fd_sc_hd__nand2_1
XFILLER_86_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4195_ egd_top.BitStream_buffer.BS_buffer\[98\] vssd1 vssd1 vccd1 vccd1 _0708_ sky130_fd_sc_hd__clkbuf_4
XFILLER_82_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6836_ net80 _0295_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BitStream_buffer_output\[13\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__2895_ _2895_ vssd1 vssd1 vccd1 vccd1 clknet_0__2895_ sky130_fd_sc_hd__clkbuf_16
XFILLER_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_330 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6767_ net171 _0226_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[53\]
+ sky130_fd_sc_hd__dfxtp_1
X_5718_ _0560_ _0498_ vssd1 vssd1 vccd1 vccd1 _2219_ sky130_fd_sc_hd__nand2_1
X_3979_ _0488_ _3053_ vssd1 vssd1 vccd1 vccd1 _0493_ sky130_fd_sc_hd__nor2_1
XFILLER_50_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5649_ _3224_ _3288_ vssd1 vssd1 vccd1 vccd1 _2151_ sky130_fd_sc_hd__nand2_1
XFILLER_40_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_34 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_67 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_66 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_88 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_87 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput7 la_data_in_58_43[15] vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__clkbuf_1
XFILLER_64_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4951_ _0682_ _3183_ _1458_ vssd1 vssd1 vccd1 vccd1 _1459_ sky130_fd_sc_hd__o21ai_1
XFILLER_17_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4882_ _0337_ _0538_ _0346_ _0541_ _1389_ vssd1 vssd1 vccd1 vccd1 _1390_ sky130_fd_sc_hd__a221oi_1
X_3902_ egd_top.BitStream_buffer.BS_buffer\[51\] vssd1 vssd1 vccd1 vccd1 _0416_ sky130_fd_sc_hd__clkbuf_4
XFILLER_17_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3833_ egd_top.BitStream_buffer.BS_buffer\[39\] vssd1 vssd1 vccd1 vccd1 _0347_ sky130_fd_sc_hd__clkbuf_4
X_3764_ _3033_ _3297_ vssd1 vssd1 vccd1 vccd1 _3298_ sky130_fd_sc_hd__nand2_2
X_5503_ _2002_ _2003_ _2004_ _2005_ vssd1 vssd1 vccd1 vccd1 _2006_ sky130_fd_sc_hd__and4_1
X_6483_ _2844_ _2845_ vssd1 vssd1 vccd1 vccd1 _2846_ sky130_fd_sc_hd__nand2_1
X_3695_ _3210_ _3216_ _3217_ _3220_ _3228_ vssd1 vssd1 vccd1 vccd1 _3229_ sky130_fd_sc_hd__a221oi_1
X_5434_ _3024_ _3200_ _1937_ vssd1 vssd1 vccd1 vccd1 _1938_ sky130_fd_sc_hd__o21ai_1
X_5365_ _0565_ egd_top.BitStream_buffer.BS_buffer\[14\] vssd1 vssd1 vccd1 vccd1 _1869_
+ sky130_fd_sc_hd__nand2_1
X_5296_ _0514_ _0540_ vssd1 vssd1 vccd1 vccd1 _1801_ sky130_fd_sc_hd__nand2_1
X_4316_ _3221_ _3216_ _3227_ _3220_ _0827_ vssd1 vssd1 vccd1 vccd1 _0828_ sky130_fd_sc_hd__a221oi_1
XFILLER_59_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4247_ _3263_ _3248_ vssd1 vssd1 vccd1 vccd1 _0760_ sky130_fd_sc_hd__nand2_1
X_4178_ _0675_ _0681_ _0684_ _0690_ vssd1 vssd1 vccd1 vccd1 _0691_ sky130_fd_sc_hd__and4_1
XFILLER_55_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6819_ net63 _0278_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[1\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_50_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_98 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3480_ net9 vssd1 vssd1 vccd1 vccd1 _3017_ sky130_fd_sc_hd__clkbuf_4
X_5150_ _0883_ _0403_ _1655_ vssd1 vssd1 vccd1 vccd1 _1656_ sky130_fd_sc_hd__o21ai_1
XFILLER_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4101_ _0602_ _0604_ _0607_ _0610_ _0614_ vssd1 vssd1 vccd1 vccd1 _0615_ sky130_fd_sc_hd__o2111a_1
X_5081_ _3027_ _1585_ _1587_ vssd1 vssd1 vccd1 vccd1 _0290_ sky130_fd_sc_hd__o21a_1
X_4032_ _0545_ vssd1 vssd1 vccd1 vccd1 _0546_ sky130_fd_sc_hd__buf_2
XFILLER_2_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5983_ egd_top.BitStream_buffer.buffer_index\[6\] egd_top.BitStream_buffer.buffer_index\[5\]
+ _2971_ vssd1 vssd1 vccd1 vccd1 _2463_ sky130_fd_sc_hd__or3_1
XFILLER_37_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4934_ _3315_ _3282_ _0774_ _1153_ _1441_ vssd1 vssd1 vccd1 vccd1 _1442_ sky130_fd_sc_hd__a221oi_1
XFILLER_24_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4865_ _0586_ _0598_ vssd1 vssd1 vccd1 vccd1 _1373_ sky130_fd_sc_hd__or2_1
XANTENNA_12 _0167_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4796_ _0505_ _0487_ _0515_ _0490_ _1304_ vssd1 vssd1 vccd1 vccd1 _1305_ sky130_fd_sc_hd__a221oi_1
X_3816_ egd_top.BitStream_buffer.BS_buffer\[92\] vssd1 vssd1 vccd1 vccd1 _0330_ sky130_fd_sc_hd__clkbuf_4
X_3747_ _3280_ vssd1 vssd1 vccd1 vccd1 _3281_ sky130_fd_sc_hd__clkbuf_2
XFILLER_21_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3678_ _3211_ _3034_ egd_top.BitStream_buffer.pc\[6\] vssd1 vssd1 vccd1 vccd1 _3212_
+ sky130_fd_sc_hd__and3_1
X_6466_ _2827_ _2829_ _2685_ vssd1 vssd1 vccd1 vccd1 _2830_ sky130_fd_sc_hd__o21ai_1
X_5417_ _3093_ _3075_ vssd1 vssd1 vccd1 vccd1 _1921_ sky130_fd_sc_hd__nand2_1
X_6397_ _2766_ _2738_ vssd1 vssd1 vccd1 vccd1 _2767_ sky130_fd_sc_hd__nand2_1
X_5348_ _1360_ _0450_ _1849_ _1850_ _1851_ vssd1 vssd1 vccd1 vccd1 _1852_ sky130_fd_sc_hd__o2111a_1
XFILLER_75_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5279_ _0371_ _0379_ vssd1 vssd1 vccd1 vccd1 _1784_ sky130_fd_sc_hd__nand2_1
XFILLER_47_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4650_ _1158_ _3299_ _1159_ vssd1 vssd1 vccd1 vccd1 _1160_ sky130_fd_sc_hd__o21ai_1
X_3601_ _3110_ _3134_ vssd1 vssd1 vccd1 vccd1 _3135_ sky130_fd_sc_hd__and2_1
Xinput10 la_data_in_58_43[3] vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__clkbuf_1
X_6320_ _2663_ _2690_ _2643_ vssd1 vssd1 vccd1 vccd1 _2691_ sky130_fd_sc_hd__or3b_1
X_4581_ _0381_ egd_top.BitStream_buffer.BS_buffer\[45\] vssd1 vssd1 vccd1 vccd1 _1091_
+ sky130_fd_sc_hd__nand2_1
X_3532_ egd_top.BitStream_buffer.BS_buffer\[108\] vssd1 vssd1 vccd1 vccd1 _3066_ sky130_fd_sc_hd__clkbuf_4
XFILLER_6_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6251_ egd_top.BitStream_buffer.BitStream_buffer_output\[13\] egd_top.BitStream_buffer.BitStream_buffer_output\[12\]
+ vssd1 vssd1 vccd1 vccd1 _2622_ sky130_fd_sc_hd__nor2_1
X_3463_ _3001_ _2975_ _3002_ _3004_ vssd1 vssd1 vccd1 vccd1 _0305_ sky130_fd_sc_hd__o211a_1
X_6182_ _2579_ _2580_ _2581_ vssd1 vssd1 vccd1 vccd1 _2582_ sky130_fd_sc_hd__a21bo_1
X_5202_ egd_top.BitStream_buffer.BitStream_buffer_output\[6\] _2965_ _0627_ vssd1
+ vssd1 vccd1 vccd1 _1707_ sky130_fd_sc_hd__o21ai_1
XFILLER_69_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3394_ _2918_ _2919_ _2947_ vssd1 vssd1 vccd1 vccd1 _2948_ sky130_fd_sc_hd__a21o_1
X_5133_ _0708_ _3324_ _3326_ _3062_ _1638_ vssd1 vssd1 vccd1 vccd1 _1639_ sky130_fd_sc_hd__a221oi_1
XFILLER_57_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5064_ _3243_ _3227_ vssd1 vssd1 vccd1 vccd1 _1571_ sky130_fd_sc_hd__nand2_1
XFILLER_72_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4015_ _0521_ _3043_ vssd1 vssd1 vccd1 vccd1 _0529_ sky130_fd_sc_hd__nand2_2
XFILLER_92_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5966_ _2449_ _0670_ vssd1 vssd1 vccd1 vccd1 _2454_ sky130_fd_sc_hd__nand2_1
X_4917_ _1413_ _1417_ _1421_ _1424_ vssd1 vssd1 vccd1 vccd1 _1425_ sky130_fd_sc_hd__and4_1
X_5897_ _1426_ _2935_ _2396_ vssd1 vssd1 vccd1 vccd1 _2397_ sky130_fd_sc_hd__o21ai_1
X_4848_ _0441_ _0459_ vssd1 vssd1 vccd1 vccd1 _1356_ sky130_fd_sc_hd__nand2_1
XFILLER_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4779_ _0653_ _0422_ _1287_ vssd1 vssd1 vccd1 vccd1 _1288_ sky130_fd_sc_hd__o21ai_1
X_6518_ _2701_ _2876_ vssd1 vssd1 vccd1 vccd1 _2879_ sky130_fd_sc_hd__nor2_1
XFILLER_4_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6449_ egd_top.BitStream_buffer.BitStream_buffer_output\[9\] _2781_ vssd1 vssd1 vccd1
+ vccd1 _2813_ sky130_fd_sc_hd__nor2_1
XFILLER_79_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5820_ _3255_ _0780_ vssd1 vssd1 vccd1 vccd1 _2320_ sky130_fd_sc_hd__nand2_1
X_5751_ _3099_ _3157_ vssd1 vssd1 vccd1 vccd1 _2252_ sky130_fd_sc_hd__nand2_1
X_4702_ _3292_ _0772_ vssd1 vssd1 vccd1 vccd1 _1211_ sky130_fd_sc_hd__nand2_1
X_5682_ _2173_ _2177_ _2180_ _2183_ vssd1 vssd1 vccd1 vccd1 _2184_ sky130_fd_sc_hd__and4_1
XFILLER_8_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4633_ _3221_ _3233_ _3227_ _3236_ _1142_ vssd1 vssd1 vccd1 vccd1 _1143_ sky130_fd_sc_hd__a221oi_1
X_4564_ _1020_ _1039_ _1056_ _1074_ vssd1 vssd1 vccd1 vccd1 _1075_ sky130_fd_sc_hd__and4_1
X_6303_ _2624_ egd_top.BitStream_buffer.BitStream_buffer_output\[13\] _2662_ vssd1
+ vssd1 vccd1 vccd1 _2674_ sky130_fd_sc_hd__or3_1
X_3515_ egd_top.BitStream_buffer.BS_buffer\[98\] vssd1 vssd1 vccd1 vccd1 _3049_ sky130_fd_sc_hd__clkinv_2
XFILLER_89_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6234_ _2998_ _2602_ _2611_ _2613_ vssd1 vssd1 vccd1 vccd1 _0169_ sky130_fd_sc_hd__o211a_1
X_4495_ _0785_ _3324_ _3326_ _3338_ _1005_ vssd1 vssd1 vccd1 vccd1 _1006_ sky130_fd_sc_hd__a221oi_1
X_3446_ _2988_ _2975_ _2913_ _2991_ vssd1 vssd1 vccd1 vccd1 _0309_ sky130_fd_sc_hd__o211a_1
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3377_ _2920_ _2930_ vssd1 vssd1 vccd1 vccd1 _2931_ sky130_fd_sc_hd__nor2_4
X_6165_ _3011_ _2555_ _2558_ _2569_ vssd1 vssd1 vccd1 vccd1 _0188_ sky130_fd_sc_hd__o211a_1
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6096_ _3020_ _2511_ _2528_ _2529_ vssd1 vssd1 vccd1 vccd1 _0217_ sky130_fd_sc_hd__o211a_1
X_5116_ _3248_ _3233_ _3236_ _3252_ _1621_ vssd1 vssd1 vccd1 vccd1 _1622_ sky130_fd_sc_hd__a221oi_1
XFILLER_84_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5047_ _0780_ _3292_ _3322_ _3295_ _1553_ vssd1 vssd1 vccd1 vccd1 _1554_ sky130_fd_sc_hd__a221oi_1
XFILLER_84_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5949_ _2966_ _2442_ _3002_ _2444_ vssd1 vssd1 vccd1 vccd1 _0279_ sky130_fd_sc_hd__o211a_1
XFILLER_4_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__2892_ clknet_0__2892_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__2892_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_88_494 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4280_ _0622_ _0792_ vssd1 vssd1 vccd1 vccd1 _0793_ sky130_fd_sc_hd__nand2_1
XTAP_203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_166 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6852_ net96 _0311_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[114\]
+ sky130_fd_sc_hd__dfxtp_2
X_5803_ _2289_ _2303_ vssd1 vssd1 vccd1 vccd1 _2304_ sky130_fd_sc_hd__nand2_1
X_3995_ egd_top.BitStream_buffer.BS_buffer\[23\] vssd1 vssd1 vccd1 vccd1 _0509_ sky130_fd_sc_hd__clkbuf_4
X_6783_ net187 _0242_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[37\]
+ sky130_fd_sc_hd__dfxtp_1
X_5734_ _0489_ _0537_ vssd1 vssd1 vccd1 vccd1 _2235_ sky130_fd_sc_hd__nand2_1
X_5665_ _3186_ egd_top.BitStream_buffer.BS_buffer\[11\] vssd1 vssd1 vccd1 vccd1 _2167_
+ sky130_fd_sc_hd__nand2_1
X_4616_ _0692_ _0604_ _1123_ _1124_ _1125_ vssd1 vssd1 vccd1 vccd1 _1126_ sky130_fd_sc_hd__o2111a_1
X_5596_ _1144_ _2935_ _2097_ vssd1 vssd1 vccd1 vccd1 _2098_ sky130_fd_sc_hd__o21ai_1
X_4547_ _3193_ egd_top.BitStream_buffer.BS_buffer\[121\] vssd1 vssd1 vccd1 vccd1 _1058_
+ sky130_fd_sc_hd__nand2_1
XFILLER_89_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4478_ _0489_ _0502_ vssd1 vssd1 vccd1 vccd1 _0989_ sky130_fd_sc_hd__nand2_1
XFILLER_89_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3429_ _2966_ _2975_ _2913_ _2978_ vssd1 vssd1 vccd1 vccd1 _0313_ sky130_fd_sc_hd__o211a_1
X_6217_ _2603_ _3296_ vssd1 vssd1 vccd1 vccd1 _2604_ sky130_fd_sc_hd__nand2_1
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6148_ _2985_ _2554_ _2558_ _2560_ vssd1 vssd1 vccd1 vccd1 _0196_ sky130_fd_sc_hd__o211a_1
XFILLER_85_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_47 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6079_ _2995_ _2510_ _2516_ _2520_ vssd1 vssd1 vccd1 vccd1 _0225_ sky130_fd_sc_hd__o211a_1
XFILLER_72_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_13 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3780_ _3313_ vssd1 vssd1 vccd1 vccd1 _3314_ sky130_fd_sc_hd__clkbuf_4
X_5450_ _3300_ _0330_ vssd1 vssd1 vccd1 vccd1 _1953_ sky130_fd_sc_hd__nand2_1
X_4401_ _0561_ _0579_ vssd1 vssd1 vccd1 vccd1 _0913_ sky130_fd_sc_hd__nand2_1
XFILLER_67_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5381_ _1857_ _1884_ vssd1 vssd1 vccd1 vccd1 _1885_ sky130_fd_sc_hd__nor2_1
XFILLER_5_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6629__6 clknet_1_0__leaf__2893_ vssd1 vssd1 vccd1 vccd1 net40 sky130_fd_sc_hd__inv_2
X_4332_ _0842_ _3299_ _0843_ vssd1 vssd1 vccd1 vccd1 _0844_ sky130_fd_sc_hd__o21ai_1
XFILLER_5_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4263_ egd_top.BitStream_buffer.BS_buffer\[88\] vssd1 vssd1 vccd1 vccd1 _0776_ sky130_fd_sc_hd__inv_2
X_6002_ _2995_ _2465_ _2474_ _2475_ vssd1 vssd1 vccd1 vccd1 _0257_ sky130_fd_sc_hd__o211a_1
X_4194_ _0669_ _0691_ _0706_ vssd1 vssd1 vccd1 vccd1 _0707_ sky130_fd_sc_hd__and3_1
XFILLER_67_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6835_ net79 _0294_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BitStream_buffer_output\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_23_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__2894_ _2894_ vssd1 vssd1 vccd1 vccd1 clknet_0__2894_ sky130_fd_sc_hd__clkbuf_16
XFILLER_50_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3978_ _0491_ vssd1 vssd1 vccd1 vccd1 _0492_ sky130_fd_sc_hd__inv_2
X_6766_ net170 _0225_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[54\]
+ sky130_fd_sc_hd__dfxtp_1
X_5717_ _2206_ _2210_ _2214_ _2217_ vssd1 vssd1 vccd1 vccd1 _2218_ sky130_fd_sc_hd__and4_1
XFILLER_40_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5648_ _3283_ _3233_ _3236_ _3276_ _2149_ vssd1 vssd1 vccd1 vccd1 _2150_ sky130_fd_sc_hd__a221oi_2
X_5579_ _2079_ _2080_ vssd1 vssd1 vccd1 vccd1 _2081_ sky130_fd_sc_hd__nor2_1
XFILLER_2_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6581__122 clknet_1_0__leaf__2889_ vssd1 vssd1 vccd1 vccd1 net156 sky130_fd_sc_hd__inv_2
XFILLER_18_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput8 la_data_in_58_43[1] vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__clkbuf_1
XFILLER_91_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4950_ _3185_ _0568_ vssd1 vssd1 vccd1 vccd1 _1458_ sky130_fd_sc_hd__nand2_1
X_4881_ _0865_ _0545_ _1388_ vssd1 vssd1 vccd1 vccd1 _1389_ sky130_fd_sc_hd__o21ai_1
X_3901_ _0414_ vssd1 vssd1 vccd1 vccd1 _0415_ sky130_fd_sc_hd__buf_2
X_3832_ egd_top.BitStream_buffer.BS_buffer\[37\] vssd1 vssd1 vccd1 vccd1 _0346_ sky130_fd_sc_hd__clkbuf_4
X_5502_ _3136_ _0568_ vssd1 vssd1 vccd1 vccd1 _2005_ sky130_fd_sc_hd__nand2_1
X_3763_ _3289_ vssd1 vssd1 vccd1 vccd1 _3297_ sky130_fd_sc_hd__clkinv_2
X_3694_ _3221_ _3224_ _3226_ _3227_ vssd1 vssd1 vccd1 vccd1 _3228_ sky130_fd_sc_hd__a22o_1
X_6482_ _2715_ _2811_ _2717_ vssd1 vssd1 vccd1 vccd1 _2845_ sky130_fd_sc_hd__o21ai_2
X_5433_ _3203_ _0741_ vssd1 vssd1 vccd1 vccd1 _1937_ sky130_fd_sc_hd__nand2_1
X_5364_ _1859_ _1861_ _1864_ _1867_ vssd1 vssd1 vccd1 vccd1 _1868_ sky130_fd_sc_hd__and4_1
XFILLER_10_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4315_ _3256_ _3224_ _3226_ _3264_ vssd1 vssd1 vccd1 vccd1 _0827_ sky130_fd_sc_hd__a22o_1
X_5295_ _0527_ _0487_ _0531_ _0490_ _1799_ vssd1 vssd1 vccd1 vccd1 _1800_ sky130_fd_sc_hd__a221oi_1
XFILLER_87_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4246_ egd_top.BitStream_buffer.BS_buffer\[73\] vssd1 vssd1 vccd1 vccd1 _0759_ sky130_fd_sc_hd__clkinv_2
X_4177_ _0685_ _0604_ _0686_ _0687_ _0689_ vssd1 vssd1 vccd1 vccd1 _0690_ sky130_fd_sc_hd__o2111a_1
XFILLER_74_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6818_ net62 _0277_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_50_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6749_ net153 _0208_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[71\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_51_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4100_ _0611_ _0613_ vssd1 vssd1 vccd1 vccd1 _0614_ sky130_fd_sc_hd__or2_1
XFILLER_69_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5080_ _1586_ _3027_ _2905_ vssd1 vssd1 vccd1 vccd1 _1587_ sky130_fd_sc_hd__a21oi_1
X_4031_ _0544_ vssd1 vssd1 vccd1 vccd1 _0545_ sky130_fd_sc_hd__clkinv_2
XFILLER_2_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6633__10 clknet_1_1__leaf__2893_ vssd1 vssd1 vccd1 vccd1 net44 sky130_fd_sc_hd__inv_2
XFILLER_37_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5982_ _3023_ _2443_ _2458_ _2462_ vssd1 vssd1 vccd1 vccd1 _0264_ sky130_fd_sc_hd__o211a_1
X_4933_ _1007_ _3273_ _1440_ vssd1 vssd1 vccd1 vccd1 _1441_ sky130_fd_sc_hd__o21ai_1
XFILLER_32_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4864_ _0922_ _0575_ _1369_ _1370_ _1371_ vssd1 vssd1 vccd1 vccd1 _1372_ sky130_fd_sc_hd__o2111a_1
XFILLER_60_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_13 _0257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4795_ _0510_ _0495_ _1303_ vssd1 vssd1 vccd1 vccd1 _1304_ sky130_fd_sc_hd__o21ai_1
X_3815_ _0328_ vssd1 vssd1 vccd1 vccd1 _0329_ sky130_fd_sc_hd__buf_4
X_3746_ _3076_ _3212_ vssd1 vssd1 vccd1 vccd1 _3280_ sky130_fd_sc_hd__and2_1
XFILLER_9_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6465_ _2823_ _2828_ vssd1 vssd1 vccd1 vccd1 _2829_ sky130_fd_sc_hd__nor2_1
XFILLER_21_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5416_ _3099_ _3169_ vssd1 vssd1 vccd1 vccd1 _1920_ sky130_fd_sc_hd__nand2_1
X_3677_ egd_top.BitStream_buffer.pc\[4\] vssd1 vssd1 vccd1 vccd1 _3211_ sky130_fd_sc_hd__inv_2
X_6396_ _2764_ _2684_ vssd1 vssd1 vccd1 vccd1 _2766_ sky130_fd_sc_hd__nand2_1
X_6612__151 clknet_1_0__leaf__2891_ vssd1 vssd1 vccd1 vccd1 net185 sky130_fd_sc_hd__inv_2
X_5347_ _0829_ _0464_ vssd1 vssd1 vccd1 vccd1 _1851_ sky130_fd_sc_hd__or2_1
XFILLER_87_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5278_ _1772_ _1775_ _1779_ _1782_ vssd1 vssd1 vccd1 vccd1 _1783_ sky130_fd_sc_hd__and4_1
XFILLER_87_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4229_ _3181_ egd_top.BitStream_buffer.BS_buffer\[127\] egd_top.BitStream_buffer.BS_buffer\[125\]
+ _3175_ vssd1 vssd1 vccd1 vccd1 _0742_ sky130_fd_sc_hd__a22o_1
XFILLER_46_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_58 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3600_ egd_top.BitStream_buffer.pc\[6\] egd_top.BitStream_buffer.pc\[4\] egd_top.BitStream_buffer.pc\[5\]
+ vssd1 vssd1 vccd1 vccd1 _3134_ sky130_fd_sc_hd__and3_2
Xinput11 la_data_in_58_43[4] vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__clkbuf_1
X_4580_ _0377_ egd_top.BitStream_buffer.BS_buffer\[44\] vssd1 vssd1 vccd1 vccd1 _1090_
+ sky130_fd_sc_hd__nand2_1
X_3531_ _3028_ _3039_ _3040_ _3048_ _3064_ vssd1 vssd1 vccd1 vccd1 _3065_ sky130_fd_sc_hd__a221oi_1
XFILLER_6_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6697__68 clknet_1_0__leaf__2899_ vssd1 vssd1 vccd1 vccd1 net102 sky130_fd_sc_hd__inv_2
X_6250_ _3023_ _2603_ _2611_ _2621_ vssd1 vssd1 vccd1 vccd1 _0161_ sky130_fd_sc_hd__o211a_1
X_3462_ _2989_ _3003_ vssd1 vssd1 vccd1 vccd1 _3004_ sky130_fd_sc_hd__nand2_1
XFILLER_69_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3393_ _2917_ _2937_ _2940_ _2946_ vssd1 vssd1 vccd1 vccd1 _2947_ sky130_fd_sc_hd__a31o_1
X_6181_ egd_top.BitStream_buffer.pc_previous\[2\] egd_top.BitStream_buffer.exp_golomb_len\[2\]
+ vssd1 vssd1 vccd1 vccd1 _2581_ sky130_fd_sc_hd__nand2_1
X_5201_ _3027_ _1704_ _1706_ vssd1 vssd1 vccd1 vccd1 _0289_ sky130_fd_sc_hd__o21a_1
XFILLER_69_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5132_ _1169_ _3330_ _1637_ vssd1 vssd1 vccd1 vccd1 _1638_ sky130_fd_sc_hd__o21ai_1
XFILLER_84_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_326 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5063_ _3302_ _3251_ _3288_ _3255_ _1569_ vssd1 vssd1 vccd1 vccd1 _1570_ sky130_fd_sc_hd__a221oi_1
X_4014_ _0527_ vssd1 vssd1 vccd1 vccd1 _0528_ sky130_fd_sc_hd__inv_2
XFILLER_37_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5965_ _2998_ _2442_ _2446_ _2453_ vssd1 vssd1 vccd1 vccd1 _0272_ sky130_fd_sc_hd__o211a_1
X_4916_ _3204_ _3078_ _0746_ _3080_ _1423_ vssd1 vssd1 vccd1 vccd1 _1424_ sky130_fd_sc_hd__a221oi_2
X_5896_ _0477_ _3268_ vssd1 vssd1 vccd1 vccd1 _2396_ sky130_fd_sc_hd__nand2_1
X_4847_ _3238_ _0450_ _1352_ _1353_ _1354_ vssd1 vssd1 vccd1 vccd1 _1355_ sky130_fd_sc_hd__o2111a_1
XFILLER_20_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4778_ _0437_ _0425_ vssd1 vssd1 vccd1 vccd1 _1287_ sky130_fd_sc_hd__or2_1
X_3729_ _3262_ vssd1 vssd1 vccd1 vccd1 _3263_ sky130_fd_sc_hd__buf_6
X_6517_ _2737_ _2695_ vssd1 vssd1 vccd1 vccd1 _2878_ sky130_fd_sc_hd__nor2_1
X_6448_ _2635_ _2811_ vssd1 vssd1 vccd1 vccd1 _2812_ sky130_fd_sc_hd__nor2_1
X_6379_ _2680_ _2748_ _2732_ vssd1 vssd1 vccd1 vccd1 _2749_ sky130_fd_sc_hd__nand3_1
XFILLER_57_24 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6619__157 clknet_1_0__leaf__2892_ vssd1 vssd1 vccd1 vccd1 net191 sky130_fd_sc_hd__inv_2
XFILLER_7_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5750_ _3070_ _3039_ _3075_ _3048_ _2250_ vssd1 vssd1 vccd1 vccd1 _2251_ sky130_fd_sc_hd__a221oi_1
XFILLER_22_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5681_ _3133_ _0726_ _3138_ _3081_ _2182_ vssd1 vssd1 vccd1 vccd1 _2183_ sky130_fd_sc_hd__a221oi_1
XFILLER_30_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4701_ _3341_ _3324_ _3326_ _3028_ _1209_ vssd1 vssd1 vccd1 vccd1 _1210_ sky130_fd_sc_hd__a221oi_1
XFILLER_30_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4632_ _3210_ _3242_ _0752_ _3217_ vssd1 vssd1 vccd1 vccd1 _1142_ sky130_fd_sc_hd__a22o_1
X_4563_ _1060_ _1065_ _1070_ _1073_ vssd1 vssd1 vccd1 vccd1 _1074_ sky130_fd_sc_hd__and4_1
X_3514_ _3047_ vssd1 vssd1 vccd1 vccd1 _3048_ sky130_fd_sc_hd__buf_6
X_6302_ _2663_ _2668_ vssd1 vssd1 vccd1 vccd1 _2673_ sky130_fd_sc_hd__nand2_1
X_4494_ _1003_ _3329_ _1004_ vssd1 vssd1 vccd1 vccd1 _1005_ sky130_fd_sc_hd__o21ai_1
XFILLER_89_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3445_ _2989_ _2990_ vssd1 vssd1 vccd1 vccd1 _2991_ sky130_fd_sc_hd__nand2_1
X_6233_ _2608_ _3306_ vssd1 vssd1 vccd1 vccd1 _2613_ sky130_fd_sc_hd__nand2_1
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3376_ _2921_ _2929_ vssd1 vssd1 vccd1 vccd1 _2930_ sky130_fd_sc_hd__or2_1
X_6164_ _2561_ _0804_ vssd1 vssd1 vccd1 vccd1 _2569_ sky130_fd_sc_hd__nand2_1
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6095_ _2509_ _0955_ vssd1 vssd1 vccd1 vccd1 _2529_ sky130_fd_sc_hd__nand2_1
X_5115_ _0759_ _3240_ _1620_ vssd1 vssd1 vccd1 vccd1 _1621_ sky130_fd_sc_hd__o21ai_1
XFILLER_84_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5046_ _3306_ _3299_ _1552_ vssd1 vssd1 vccd1 vccd1 _1553_ sky130_fd_sc_hd__o21ai_1
XFILLER_27_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5948_ _2443_ _1602_ vssd1 vssd1 vccd1 vccd1 _2444_ sky130_fd_sc_hd__nand2_1
XFILLER_40_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5879_ _0371_ _0407_ vssd1 vssd1 vccd1 vccd1 _2379_ sky130_fd_sc_hd__nand2_1
XFILLER_4_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6676__49 clknet_1_1__leaf__2897_ vssd1 vssd1 vccd1 vccd1 net83 sky130_fd_sc_hd__inv_2
Xclkbuf_1_1__f__2891_ clknet_0__2891_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__2891_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_29_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_66 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6851_ net95 _0310_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[115\]
+ sky130_fd_sc_hd__dfxtp_1
X_5802_ _2292_ _2296_ _2299_ _2302_ vssd1 vssd1 vccd1 vccd1 _2303_ sky130_fd_sc_hd__and4_1
X_3994_ _0507_ vssd1 vssd1 vccd1 vccd1 _0508_ sky130_fd_sc_hd__buf_6
XFILLER_22_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6782_ net186 _0241_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[38\]
+ sky130_fd_sc_hd__dfxtp_1
X_5733_ _0486_ egd_top.BitStream_buffer.BS_buffer\[29\] vssd1 vssd1 vccd1 vccd1 _2234_
+ sky130_fd_sc_hd__nand2_1
XFILLER_13_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5664_ _0930_ _3194_ _3197_ _1076_ _2165_ vssd1 vssd1 vccd1 vccd1 _2166_ sky130_fd_sc_hd__a221oi_1
X_4615_ _0922_ _0612_ vssd1 vssd1 vccd1 vccd1 _1125_ sky130_fd_sc_hd__or2_1
X_5595_ _0476_ egd_top.BitStream_buffer.BS_buffer\[74\] vssd1 vssd1 vccd1 vccd1 _2097_
+ sky130_fd_sc_hd__nand2_1
X_4546_ _3202_ _3198_ vssd1 vssd1 vccd1 vccd1 _1057_ sky130_fd_sc_hd__nand2_1
X_4477_ _0496_ _0515_ vssd1 vssd1 vccd1 vccd1 _0988_ sky130_fd_sc_hd__nand2_1
X_3428_ _2976_ _2977_ vssd1 vssd1 vccd1 vccd1 _2978_ sky130_fd_sc_hd__nand2_1
X_6216_ _2601_ vssd1 vssd1 vccd1 vccd1 _2603_ sky130_fd_sc_hd__buf_2
XFILLER_85_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3359_ _2911_ _2906_ _2905_ vssd1 vssd1 vccd1 vccd1 _2914_ sky130_fd_sc_hd__a21o_1
X_6147_ _2555_ _0709_ vssd1 vssd1 vccd1 vccd1 _2560_ sky130_fd_sc_hd__nand2_1
XFILLER_85_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6078_ _2517_ _0653_ vssd1 vssd1 vccd1 vccd1 _2520_ sky130_fd_sc_hd__nand2_1
X_5029_ _1525_ _1529_ _1532_ _1535_ vssd1 vssd1 vccd1 vccd1 _1536_ sky130_fd_sc_hd__and4_1
XFILLER_54_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_46 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4400_ _0565_ _0562_ vssd1 vssd1 vccd1 vccd1 _0912_ sky130_fd_sc_hd__nand2_1
X_5380_ _1868_ _1883_ vssd1 vssd1 vccd1 vccd1 _1884_ sky130_fd_sc_hd__nand2_1
XFILLER_5_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4331_ _3301_ _3293_ vssd1 vssd1 vccd1 vccd1 _0843_ sky130_fd_sc_hd__nand2_1
X_4262_ _3314_ _0774_ vssd1 vssd1 vccd1 vccd1 _0775_ sky130_fd_sc_hd__nand2_1
XFILLER_39_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6001_ _2471_ _1128_ vssd1 vssd1 vccd1 vccd1 _2475_ sky130_fd_sc_hd__nand2_1
X_4193_ _0695_ _0698_ _0701_ _0705_ vssd1 vssd1 vccd1 vccd1 _0706_ sky130_fd_sc_hd__and4_1
XFILLER_79_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6834_ net78 _0293_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BitStream_buffer_output\[11\]
+ sky130_fd_sc_hd__dfxtp_2
Xclkbuf_0__2893_ _2893_ vssd1 vssd1 vccd1 vccd1 clknet_0__2893_ sky130_fd_sc_hd__clkbuf_16
XFILLER_35_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3977_ egd_top.BitStream_buffer.BS_buffer\[18\] vssd1 vssd1 vccd1 vccd1 _0491_ sky130_fd_sc_hd__clkbuf_4
X_6765_ net169 _0224_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[55\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_50_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5716_ _3252_ _0477_ _3268_ _2936_ _2216_ vssd1 vssd1 vccd1 vccd1 _2217_ sky130_fd_sc_hd__a221oi_1
X_5647_ _1426_ _3240_ _2148_ vssd1 vssd1 vccd1 vccd1 _2149_ sky130_fd_sc_hd__o21ai_1
X_5578_ _3087_ _0416_ _0339_ _0412_ _0352_ vssd1 vssd1 vccd1 vccd1 _2080_ sky130_fd_sc_hd__a32o_1
X_4529_ _3215_ _3227_ vssd1 vssd1 vccd1 vccd1 _1040_ sky130_fd_sc_hd__nand2_1
XFILLER_2_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput9 la_data_in_58_43[2] vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__clkbuf_1
XFILLER_49_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4880_ _0547_ egd_top.BitStream_buffer.BS_buffer\[34\] vssd1 vssd1 vccd1 vccd1 _1388_
+ sky130_fd_sc_hd__nand2_1
XFILLER_32_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3900_ _0413_ vssd1 vssd1 vccd1 vccd1 _0414_ sky130_fd_sc_hd__clkbuf_2
XFILLER_44_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3831_ _0344_ vssd1 vssd1 vccd1 vccd1 _0345_ sky130_fd_sc_hd__buf_6
X_6631__8 clknet_1_0__leaf__2893_ vssd1 vssd1 vccd1 vccd1 net42 sky130_fd_sc_hd__inv_2
X_3762_ egd_top.BitStream_buffer.BS_buffer\[80\] vssd1 vssd1 vccd1 vccd1 _3296_ sky130_fd_sc_hd__clkinv_2
X_5501_ _3144_ _1076_ vssd1 vssd1 vccd1 vccd1 _2004_ sky130_fd_sc_hd__nand2_1
X_6481_ _2842_ _2843_ _2681_ vssd1 vssd1 vccd1 vccd1 _2844_ sky130_fd_sc_hd__nand3_1
X_3693_ egd_top.BitStream_buffer.BS_buffer\[71\] vssd1 vssd1 vccd1 vccd1 _3227_ sky130_fd_sc_hd__clkbuf_4
X_5432_ _0553_ _3180_ _0585_ _3186_ _1935_ vssd1 vssd1 vccd1 vccd1 _1936_ sky130_fd_sc_hd__a221oi_1
X_5363_ _0375_ _0539_ _0379_ _0542_ _1866_ vssd1 vssd1 vccd1 vccd1 _1867_ sky130_fd_sc_hd__a221oi_2
X_4314_ _0812_ _0825_ vssd1 vssd1 vccd1 vccd1 _0826_ sky130_fd_sc_hd__nand2_1
XFILLER_87_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5294_ _0524_ _0495_ _1798_ vssd1 vssd1 vccd1 vccd1 _1799_ sky130_fd_sc_hd__o21ai_1
X_4245_ _3227_ _3224_ _3256_ _3226_ _0757_ vssd1 vssd1 vccd1 vccd1 _0758_ sky130_fd_sc_hd__a221oi_1
X_4176_ _0688_ _0613_ vssd1 vssd1 vccd1 vccd1 _0689_ sky130_fd_sc_hd__or2_1
XFILLER_55_413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6817_ net61 _0276_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_23_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6748_ net152 _0207_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[72\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_50_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6679_ clknet_1_0__leaf__2882_ vssd1 vssd1 vccd1 vccd1 _2898_ sky130_fd_sc_hd__buf_1
XFILLER_2_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6548__92 clknet_1_0__leaf__2886_ vssd1 vssd1 vccd1 vccd1 net126 sky130_fd_sc_hd__inv_2
XFILLER_41_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6588__129 clknet_1_0__leaf__2889_ vssd1 vssd1 vccd1 vccd1 net163 sky130_fd_sc_hd__inv_2
XFILLER_69_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4030_ _0488_ _3072_ vssd1 vssd1 vccd1 vccd1 _0544_ sky130_fd_sc_hd__nor2_1
X_5981_ _2441_ _0602_ vssd1 vssd1 vccd1 vccd1 _2462_ sky130_fd_sc_hd__nand2_1
X_4932_ _3270_ egd_top.BitStream_buffer.BS_buffer\[82\] vssd1 vssd1 vccd1 vccd1 _1440_
+ sky130_fd_sc_hd__nand2_1
XFILLER_17_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4863_ _0602_ _0587_ vssd1 vssd1 vccd1 vccd1 _1371_ sky130_fd_sc_hd__or2_1
X_6602_ clknet_1_1__leaf__2883_ vssd1 vssd1 vccd1 vccd1 _2891_ sky130_fd_sc_hd__buf_1
XANTENNA_14 _2992_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4794_ _0497_ _0519_ vssd1 vssd1 vccd1 vccd1 _1303_ sky130_fd_sc_hd__nand2_1
X_3814_ _3290_ _3068_ vssd1 vssd1 vccd1 vccd1 _0328_ sky130_fd_sc_hd__nor2_2
XFILLER_20_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3745_ _3278_ vssd1 vssd1 vccd1 vccd1 _3279_ sky130_fd_sc_hd__clkbuf_4
X_6464_ _2767_ _2786_ vssd1 vssd1 vccd1 vccd1 _2828_ sky130_fd_sc_hd__nor2_1
X_5415_ _3109_ _3039_ _3118_ _3048_ _1918_ vssd1 vssd1 vccd1 vccd1 _1919_ sky130_fd_sc_hd__a221oi_2
X_3676_ egd_top.BitStream_buffer.BS_buffer\[68\] vssd1 vssd1 vccd1 vccd1 _3210_ sky130_fd_sc_hd__clkbuf_4
X_6395_ _2739_ _2764_ vssd1 vssd1 vccd1 vccd1 _2765_ sky130_fd_sc_hd__nand2_1
X_5346_ _0458_ _3210_ vssd1 vssd1 vccd1 vccd1 _1850_ sky130_fd_sc_hd__nand2_1
X_5277_ _3217_ _0470_ _3221_ _0473_ _1781_ vssd1 vssd1 vccd1 vccd1 _1782_ sky130_fd_sc_hd__a221oi_1
X_4228_ egd_top.BitStream_buffer.BS_buffer\[126\] vssd1 vssd1 vccd1 vccd1 _0741_ sky130_fd_sc_hd__buf_2
XFILLER_46_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4159_ _0561_ _0553_ vssd1 vssd1 vccd1 vccd1 _0672_ sky130_fd_sc_hd__nand2_1
XFILLER_55_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput12 la_data_in_58_43[5] vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__clkbuf_1
X_3530_ _3049_ _3056_ _3063_ vssd1 vssd1 vccd1 vccd1 _3064_ sky130_fd_sc_hd__o21ai_1
X_3461_ egd_top.BitStream_buffer.BS_buffer\[120\] vssd1 vssd1 vccd1 vccd1 _3003_ sky130_fd_sc_hd__clkinv_2
X_5200_ _1705_ _3027_ _2905_ vssd1 vssd1 vccd1 vccd1 _1706_ sky130_fd_sc_hd__a21oi_1
X_3392_ _2943_ _2945_ _2918_ vssd1 vssd1 vccd1 vccd1 _2946_ sky130_fd_sc_hd__a21oi_1
X_6180_ egd_top.BitStream_buffer.pc_previous\[2\] egd_top.BitStream_buffer.exp_golomb_len\[2\]
+ vssd1 vssd1 vccd1 vccd1 _2580_ sky130_fd_sc_hd__or2_1
XFILLER_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5131_ _3333_ _3028_ vssd1 vssd1 vccd1 vccd1 _1637_ sky130_fd_sc_hd__nand2_1
X_5062_ _3277_ _3260_ _1568_ vssd1 vssd1 vccd1 vccd1 _1569_ sky130_fd_sc_hd__o21ai_1
XFILLER_69_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4013_ egd_top.BitStream_buffer.BS_buffer\[25\] vssd1 vssd1 vccd1 vccd1 _0527_ sky130_fd_sc_hd__clkbuf_4
XFILLER_84_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f__2899_ clknet_0__2899_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__2899_
+ sky130_fd_sc_hd__clkbuf_16
X_5964_ _2449_ _0554_ vssd1 vssd1 vccd1 vccd1 _2453_ sky130_fd_sc_hd__nand2_1
X_4915_ _2983_ _0728_ _1422_ vssd1 vssd1 vccd1 vccd1 _1423_ sky130_fd_sc_hd__o21ai_1
XFILLER_52_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5895_ _0759_ _0450_ _2392_ _2393_ _2394_ vssd1 vssd1 vccd1 vccd1 _2395_ sky130_fd_sc_hd__o2111a_1
XFILLER_40_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4846_ _0474_ _0463_ vssd1 vssd1 vccd1 vccd1 _1354_ sky130_fd_sc_hd__or2_1
XFILLER_32_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6516_ _2870_ _2701_ _2876_ vssd1 vssd1 vccd1 vccd1 _2877_ sky130_fd_sc_hd__nand3_1
X_6527__73 clknet_1_0__leaf__2884_ vssd1 vssd1 vccd1 vccd1 net107 sky130_fd_sc_hd__inv_2
X_4777_ _1275_ _1279_ _1282_ _1285_ vssd1 vssd1 vccd1 vccd1 _1286_ sky130_fd_sc_hd__and4_1
X_3728_ _3261_ vssd1 vssd1 vccd1 vccd1 _3262_ sky130_fd_sc_hd__clkbuf_2
XFILLER_4_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3659_ _3192_ vssd1 vssd1 vccd1 vccd1 _3193_ sky130_fd_sc_hd__clkbuf_2
X_6447_ _2781_ vssd1 vssd1 vccd1 vccd1 _2811_ sky130_fd_sc_hd__inv_2
X_6378_ _2626_ _2723_ _2747_ vssd1 vssd1 vccd1 vccd1 _2748_ sky130_fd_sc_hd__o21ai_1
X_6542__87 clknet_1_1__leaf__2885_ vssd1 vssd1 vccd1 vccd1 net121 sky130_fd_sc_hd__inv_2
XFILLER_0_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5329_ _0353_ _0874_ vssd1 vssd1 vccd1 vccd1 _1833_ sky130_fd_sc_hd__nand2_1
XFILLER_87_143 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_508 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_36 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5680_ _3003_ _0729_ _2181_ vssd1 vssd1 vccd1 vccd1 _2182_ sky130_fd_sc_hd__o21ai_1
X_4700_ _0784_ _3330_ _1208_ vssd1 vssd1 vccd1 vccd1 _1209_ sky130_fd_sc_hd__o21ai_1
X_4631_ _1112_ _1127_ _1140_ vssd1 vssd1 vccd1 vccd1 _1141_ sky130_fd_sc_hd__and3_1
XFILLER_30_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4562_ _3187_ _3176_ _0623_ _3179_ _1072_ vssd1 vssd1 vccd1 vccd1 _1073_ sky130_fd_sc_hd__a221oi_1
X_3513_ _3041_ _3046_ vssd1 vssd1 vccd1 vccd1 _3047_ sky130_fd_sc_hd__nor2_2
X_6301_ _2661_ _2666_ _2671_ vssd1 vssd1 vccd1 vccd1 _2672_ sky130_fd_sc_hd__nand3_1
X_4493_ _3332_ _3327_ vssd1 vssd1 vccd1 vccd1 _1004_ sky130_fd_sc_hd__nand2_1
X_3444_ egd_top.BitStream_buffer.BS_buffer\[116\] vssd1 vssd1 vccd1 vccd1 _2990_ sky130_fd_sc_hd__inv_2
X_6232_ _2995_ _2602_ _2611_ _2612_ vssd1 vssd1 vccd1 vccd1 _0170_ sky130_fd_sc_hd__o211a_1
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3375_ _2925_ _2928_ vssd1 vssd1 vccd1 vccd1 _2929_ sky130_fd_sc_hd__nand2_2
X_6163_ _3008_ _2555_ _2558_ _2568_ vssd1 vssd1 vccd1 vccd1 _0189_ sky130_fd_sc_hd__o211a_1
XFILLER_84_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6094_ _2904_ vssd1 vssd1 vccd1 vccd1 _2528_ sky130_fd_sc_hd__buf_2
X_5114_ _3243_ _3256_ vssd1 vssd1 vccd1 vccd1 _1620_ sky130_fd_sc_hd__nand2_1
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5045_ _3301_ _3334_ vssd1 vssd1 vccd1 vccd1 _1552_ sky130_fd_sc_hd__nand2_1
XFILLER_27_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5947_ _2441_ vssd1 vssd1 vccd1 vccd1 _2443_ sky130_fd_sc_hd__buf_2
XFILLER_43_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5878_ _0429_ _0378_ _0436_ _0382_ _2377_ vssd1 vssd1 vccd1 vccd1 _2378_ sky130_fd_sc_hd__a221oi_1
X_4829_ _0870_ _0350_ _1336_ vssd1 vssd1 vccd1 vccd1 _1337_ sky130_fd_sc_hd__o21ai_1
XFILLER_21_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__2890_ clknet_0__2890_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__2890_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_75_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1 egd_top.BitStream_buffer.buffer_index\[5\] vssd1 vssd1 vccd1 vccd1 net196 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_81_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6850_ net94 _0309_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[116\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_47_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5801_ _3118_ _3340_ _3066_ _0323_ _2301_ vssd1 vssd1 vccd1 vccd1 _2302_ sky130_fd_sc_hd__a221oi_1
X_6781_ net185 _0240_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[39\]
+ sky130_fd_sc_hd__dfxtp_1
X_3993_ _0506_ vssd1 vssd1 vccd1 vccd1 _0507_ sky130_fd_sc_hd__inv_2
X_5732_ _2222_ _2226_ _2228_ _2232_ vssd1 vssd1 vccd1 vccd1 _2233_ sky130_fd_sc_hd__and4_1
XFILLER_50_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5663_ _0594_ _3200_ _2164_ vssd1 vssd1 vccd1 vccd1 _2165_ sky130_fd_sc_hd__o21ai_1
X_4614_ _0605_ egd_top.BitStream_buffer.BS_buffer\[16\] vssd1 vssd1 vccd1 vccd1 _1124_
+ sky130_fd_sc_hd__nand2_1
X_5594_ _3238_ _0439_ _2093_ _2094_ _2095_ vssd1 vssd1 vccd1 vccd1 _2096_ sky130_fd_sc_hd__o2111a_1
X_4545_ _1042_ _1047_ _1052_ _1055_ vssd1 vssd1 vccd1 vccd1 _1056_ sky130_fd_sc_hd__and4_1
XFILLER_89_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4476_ _0486_ _0498_ vssd1 vssd1 vccd1 vccd1 _0987_ sky130_fd_sc_hd__nand2_1
X_6215_ _2601_ vssd1 vssd1 vccd1 vccd1 _2602_ sky130_fd_sc_hd__buf_2
X_3427_ egd_top.BitStream_buffer.BS_buffer\[112\] vssd1 vssd1 vccd1 vccd1 _2977_ sky130_fd_sc_hd__inv_2
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3358_ net32 _2912_ _2913_ _2907_ vssd1 vssd1 vccd1 vccd1 _0319_ sky130_fd_sc_hd__o211a_1
X_6146_ _2982_ _2554_ _2558_ _2559_ vssd1 vssd1 vccd1 vccd1 _0197_ sky130_fd_sc_hd__o211a_1
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6077_ _2992_ _2510_ _2516_ _2519_ vssd1 vssd1 vccd1 vccd1 _0226_ sky130_fd_sc_hd__o211a_1
X_6681__53 clknet_1_0__leaf__2898_ vssd1 vssd1 vccd1 vccd1 net87 sky130_fd_sc_hd__inv_2
X_5028_ _0746_ _0726_ _3191_ _3081_ _1534_ vssd1 vssd1 vccd1 vccd1 _1535_ sky130_fd_sc_hd__a221oi_1
XFILLER_72_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4330_ egd_top.BitStream_buffer.BS_buffer\[82\] vssd1 vssd1 vccd1 vccd1 _0842_ sky130_fd_sc_hd__clkinv_2
X_4261_ egd_top.BitStream_buffer.BS_buffer\[85\] vssd1 vssd1 vccd1 vccd1 _0774_ sky130_fd_sc_hd__clkbuf_4
X_6000_ _2901_ vssd1 vssd1 vccd1 vccd1 _2474_ sky130_fd_sc_hd__buf_2
X_4192_ _0540_ _0539_ egd_top.BitStream_buffer.BS_buffer\[32\] _0542_ _0704_ vssd1
+ vssd1 vccd1 vccd1 _0705_ sky130_fd_sc_hd__a221oi_1
XFILLER_67_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6833_ net77 _0292_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BitStream_buffer_output\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_24_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__2892_ _2892_ vssd1 vssd1 vccd1 vccd1 clknet_0__2892_ sky130_fd_sc_hd__clkbuf_16
X_3976_ _0489_ vssd1 vssd1 vccd1 vccd1 _0490_ sky130_fd_sc_hd__buf_6
X_6764_ net168 _0223_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[56\]
+ sky130_fd_sc_hd__dfxtp_1
X_5715_ _0833_ _0472_ _2215_ vssd1 vssd1 vccd1 vccd1 _2216_ sky130_fd_sc_hd__o21ai_1
X_5646_ _3243_ _3268_ vssd1 vssd1 vccd1 vccd1 _2148_ sky130_fd_sc_hd__nand2_1
X_5577_ egd_top.BitStream_buffer.BS_buffer\[48\] _0341_ _0344_ _0948_ vssd1 vssd1
+ vccd1 vccd1 _2079_ sky130_fd_sc_hd__a22o_1
X_4528_ _1024_ _1029_ _1034_ _1038_ vssd1 vssd1 vccd1 vccd1 _1039_ sky130_fd_sc_hd__and4_1
XFILLER_2_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4459_ _0954_ _0959_ _0964_ _0969_ vssd1 vssd1 vccd1 vccd1 _0970_ sky130_fd_sc_hd__and4_1
XFILLER_49_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6129_ _3014_ _2533_ _2543_ _2548_ vssd1 vssd1 vccd1 vccd1 _0203_ sky130_fd_sc_hd__o211a_1
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_355 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6660__34 clknet_1_0__leaf__2896_ vssd1 vssd1 vccd1 vccd1 net68 sky130_fd_sc_hd__inv_2
XFILLER_36_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_80 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3830_ _0343_ vssd1 vssd1 vccd1 vccd1 _0344_ sky130_fd_sc_hd__clkbuf_2
X_3761_ _3294_ vssd1 vssd1 vccd1 vccd1 _3295_ sky130_fd_sc_hd__buf_6
X_5500_ _3140_ _0562_ vssd1 vssd1 vccd1 vccd1 _2003_ sky130_fd_sc_hd__nand2_1
XFILLER_72_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3692_ _3225_ vssd1 vssd1 vccd1 vccd1 _3226_ sky130_fd_sc_hd__inv_2
X_6480_ _2802_ _2804_ _2840_ vssd1 vssd1 vccd1 vccd1 _2843_ sky130_fd_sc_hd__nand3_1
X_5431_ _3181_ _0579_ _0562_ _3176_ vssd1 vssd1 vccd1 vccd1 _1935_ sky130_fd_sc_hd__a22o_1
X_5362_ _0348_ _0546_ _1865_ vssd1 vssd1 vccd1 vccd1 _1866_ sky130_fd_sc_hd__o21ai_1
X_4313_ _0815_ _0819_ _0821_ _0824_ vssd1 vssd1 vccd1 vccd1 _0825_ sky130_fd_sc_hd__and4_1
XFILLER_87_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5293_ _0497_ egd_top.BitStream_buffer.BS_buffer\[28\] vssd1 vssd1 vccd1 vccd1 _1798_
+ sky130_fd_sc_hd__nand2_1
X_4244_ _0755_ _3218_ _0756_ vssd1 vssd1 vccd1 vccd1 _0757_ sky130_fd_sc_hd__o21ai_1
XFILLER_19_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6565__108 clknet_1_1__leaf__2887_ vssd1 vssd1 vccd1 vccd1 net142 sky130_fd_sc_hd__inv_2
X_4175_ egd_top.BitStream_buffer.BS_buffer\[14\] vssd1 vssd1 vccd1 vccd1 _0688_ sky130_fd_sc_hd__inv_2
XFILLER_67_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6816_ net60 _0275_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[4\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_23_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6747_ net151 _0206_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[73\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_50_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3959_ _0472_ vssd1 vssd1 vccd1 vccd1 _0473_ sky130_fd_sc_hd__inv_2
X_5629_ _3301_ _0785_ vssd1 vssd1 vccd1 vccd1 _2131_ sky130_fd_sc_hd__nand2_1
XFILLER_2_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5980_ _3020_ _2443_ _2458_ _2461_ vssd1 vssd1 vccd1 vccd1 _0265_ sky130_fd_sc_hd__o211a_1
XFILLER_17_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4931_ _1435_ _1436_ _1437_ _1438_ vssd1 vssd1 vccd1 vccd1 _1439_ sky130_fd_sc_hd__and4_1
XFILLER_45_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4862_ _0577_ egd_top.BitStream_buffer.BS_buffer\[14\] vssd1 vssd1 vccd1 vccd1 _1370_
+ sky130_fd_sc_hd__nand2_1
XFILLER_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3813_ _0326_ vssd1 vssd1 vccd1 vccd1 _0327_ sky130_fd_sc_hd__buf_2
XFILLER_20_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_15 _2992_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4793_ _1286_ _1301_ vssd1 vssd1 vccd1 vccd1 _1302_ sky130_fd_sc_hd__nand2_1
X_3744_ _2931_ _3213_ vssd1 vssd1 vccd1 vccd1 _3278_ sky130_fd_sc_hd__nand2_1
X_3675_ _3132_ _3208_ vssd1 vssd1 vccd1 vccd1 _3209_ sky130_fd_sc_hd__nand2_1
X_6463_ _2824_ _2826_ vssd1 vssd1 vccd1 vccd1 _2827_ sky130_fd_sc_hd__nor2_1
X_5414_ _1025_ _3056_ _1917_ vssd1 vssd1 vccd1 vccd1 _1918_ sky130_fd_sc_hd__o21ai_1
X_6394_ _2750_ _2763_ vssd1 vssd1 vccd1 vccd1 _2764_ sky130_fd_sc_hd__nand2_2
X_5345_ _0453_ _3230_ vssd1 vssd1 vccd1 vccd1 _1849_ sky130_fd_sc_hd__nand2_1
X_5276_ _3257_ _2935_ _1780_ vssd1 vssd1 vccd1 vccd1 _1781_ sky130_fd_sc_hd__o21ai_1
X_4227_ _3157_ _3156_ _3204_ _3160_ _0739_ vssd1 vssd1 vccd1 vccd1 _0740_ sky130_fd_sc_hd__a221oi_2
X_4158_ _0565_ _0568_ vssd1 vssd1 vccd1 vccd1 _0671_ sky130_fd_sc_hd__nand2_1
XFILLER_55_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4089_ _2931_ _0556_ vssd1 vssd1 vccd1 vccd1 _0603_ sky130_fd_sc_hd__nand2_1
XFILLER_55_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6594__134 clknet_1_1__leaf__2890_ vssd1 vssd1 vccd1 vccd1 net168 sky130_fd_sc_hd__inv_2
XFILLER_42_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput13 la_data_in_58_43[6] vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__clkbuf_1
XFILLER_6_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3460_ _2901_ vssd1 vssd1 vccd1 vccd1 _3002_ sky130_fd_sc_hd__buf_2
X_3391_ _2944_ egd_top.BitStream_buffer.pc_previous\[6\] _2932_ vssd1 vssd1 vccd1
+ vccd1 _2945_ sky130_fd_sc_hd__a21o_1
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5130_ _0854_ _3308_ _1633_ _1634_ _1635_ vssd1 vssd1 vccd1 vccd1 _1636_ sky130_fd_sc_hd__o2111a_1
X_5061_ _3263_ _0837_ vssd1 vssd1 vccd1 vccd1 _1568_ sky130_fd_sc_hd__nand2_1
X_4012_ _0525_ vssd1 vssd1 vccd1 vccd1 _0526_ sky130_fd_sc_hd__buf_2
XFILLER_77_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_0__f__2898_ clknet_0__2898_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__2898_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_25_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5963_ _2995_ _2442_ _2446_ _2452_ vssd1 vssd1 vccd1 vccd1 _0273_ sky130_fd_sc_hd__o211a_1
X_4914_ _3073_ _3157_ vssd1 vssd1 vccd1 vccd1 _1422_ sky130_fd_sc_hd__nand2_1
X_5894_ _1430_ _0464_ vssd1 vssd1 vccd1 vccd1 _2394_ sky130_fd_sc_hd__or2_1
XFILLER_33_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4845_ _0457_ _3244_ vssd1 vssd1 vccd1 vccd1 _1353_ sky130_fd_sc_hd__nand2_1
XFILLER_32_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4776_ _0948_ _0396_ _0399_ _0412_ _1284_ vssd1 vssd1 vccd1 vccd1 _1285_ sky130_fd_sc_hd__a221oi_1
X_3727_ _3121_ _3212_ vssd1 vssd1 vccd1 vccd1 _3261_ sky130_fd_sc_hd__and2_1
X_6515_ _2695_ _2875_ vssd1 vssd1 vccd1 vccd1 _2876_ sky130_fd_sc_hd__or2_1
X_3658_ _3096_ _3142_ vssd1 vssd1 vccd1 vccd1 _3192_ sky130_fd_sc_hd__and2_1
X_6446_ _2806_ _2809_ _2681_ vssd1 vssd1 vccd1 vccd1 _2810_ sky130_fd_sc_hd__nand3_1
X_3589_ _3122_ vssd1 vssd1 vccd1 vccd1 _3123_ sky130_fd_sc_hd__clkbuf_4
X_6377_ _2723_ egd_top.BitStream_buffer.BitStream_buffer_output\[5\] vssd1 vssd1 vccd1
+ vccd1 _2747_ sky130_fd_sc_hd__nand2_1
XFILLER_87_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5328_ _0393_ _0360_ _0363_ _0400_ _1831_ vssd1 vssd1 vccd1 vccd1 _1832_ sky130_fd_sc_hd__a221oi_2
XFILLER_0_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5259_ _3138_ _3155_ _3173_ _3159_ _1763_ vssd1 vssd1 vccd1 vccd1 _1764_ sky130_fd_sc_hd__a221oi_1
XFILLER_75_306 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4630_ _1131_ _1134_ _1136_ _1139_ vssd1 vssd1 vccd1 vccd1 _1140_ sky130_fd_sc_hd__and4_1
XFILLER_8_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4561_ _0594_ _3183_ _1071_ vssd1 vssd1 vccd1 vccd1 _1072_ sky130_fd_sc_hd__o21ai_1
XFILLER_8_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6300_ _2670_ _1705_ vssd1 vssd1 vccd1 vccd1 _2671_ sky130_fd_sc_hd__nand2_1
X_3512_ _3045_ vssd1 vssd1 vccd1 vccd1 _3046_ sky130_fd_sc_hd__clkinv_2
XFILLER_6_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4492_ egd_top.BitStream_buffer.BS_buffer\[92\] vssd1 vssd1 vccd1 vccd1 _1003_ sky130_fd_sc_hd__clkinv_2
X_3443_ _2974_ vssd1 vssd1 vccd1 vccd1 _2989_ sky130_fd_sc_hd__buf_2
X_6231_ _2608_ _0771_ vssd1 vssd1 vccd1 vccd1 _2612_ sky130_fd_sc_hd__nand2_1
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6162_ _2561_ _0721_ vssd1 vssd1 vccd1 vccd1 _2568_ sky130_fd_sc_hd__nand2_1
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5113_ _0837_ _3259_ _3302_ _3263_ _1618_ vssd1 vssd1 vccd1 vccd1 _1619_ sky130_fd_sc_hd__a221oi_1
X_3374_ _2926_ _2927_ vssd1 vssd1 vccd1 vccd1 _2928_ sky130_fd_sc_hd__nand2_1
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6093_ _3017_ _2511_ _2516_ _2527_ vssd1 vssd1 vccd1 vccd1 _0218_ sky130_fd_sc_hd__o211a_1
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5044_ _1536_ _1550_ vssd1 vssd1 vccd1 vccd1 _1551_ sky130_fd_sc_hd__nand2_1
XFILLER_69_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5946_ _2441_ vssd1 vssd1 vccd1 vccd1 _2442_ sky130_fd_sc_hd__buf_2
X_5877_ _0462_ _0385_ _2376_ vssd1 vssd1 vccd1 vccd1 _2377_ sky130_fd_sc_hd__o21ai_1
X_4828_ _0353_ _0393_ vssd1 vssd1 vccd1 vccd1 _1336_ sky130_fd_sc_hd__nand2_1
X_4759_ _3281_ egd_top.BitStream_buffer.BS_buffer\[83\] vssd1 vssd1 vccd1 vccd1 _1268_
+ sky130_fd_sc_hd__nand2_1
X_6429_ _2795_ _2698_ _2796_ vssd1 vssd1 vccd1 vccd1 _2797_ sky130_fd_sc_hd__nand3_1
XFILLER_68_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2 _2600_ vssd1 vssd1 vccd1 vccd1 net197 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_54_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3992_ _3104_ _0484_ vssd1 vssd1 vccd1 vccd1 _0506_ sky130_fd_sc_hd__nand2_1
X_5800_ _0721_ _0327_ _2300_ vssd1 vssd1 vccd1 vccd1 _2301_ sky130_fd_sc_hd__o21ai_1
X_6780_ net184 _0239_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[40\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_50_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5731_ _0699_ _0603_ _2229_ _2230_ _2231_ vssd1 vssd1 vccd1 vccd1 _2232_ sky130_fd_sc_hd__o2111a_1
X_5662_ _3203_ _0623_ vssd1 vssd1 vccd1 vccd1 _2164_ sky130_fd_sc_hd__nand2_1
X_4613_ _0608_ _0491_ vssd1 vssd1 vccd1 vccd1 _1123_ sky130_fd_sc_hd__nand2_1
X_5593_ _0434_ _3237_ vssd1 vssd1 vccd1 vccd1 _2095_ sky130_fd_sc_hd__nand2_1
X_4544_ _3276_ _3270_ _0837_ _3274_ _1054_ vssd1 vssd1 vccd1 vccd1 _1055_ sky130_fd_sc_hd__a221oi_1
X_4475_ _0505_ vssd1 vssd1 vccd1 vccd1 _0986_ sky130_fd_sc_hd__inv_2
X_6214_ net197 vssd1 vssd1 vccd1 vccd1 _2601_ sky130_fd_sc_hd__inv_2
X_6666__40 clknet_1_1__leaf__2896_ vssd1 vssd1 vccd1 vccd1 net74 sky130_fd_sc_hd__inv_2
X_3426_ _2974_ vssd1 vssd1 vccd1 vccd1 _2976_ sky130_fd_sc_hd__buf_2
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3357_ _2901_ vssd1 vssd1 vccd1 vccd1 _2913_ sky130_fd_sc_hd__clkbuf_4
X_6145_ _2555_ _3049_ vssd1 vssd1 vccd1 vccd1 _2559_ sky130_fd_sc_hd__nand2_1
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6076_ _2517_ _0437_ vssd1 vssd1 vccd1 vccd1 _2519_ sky130_fd_sc_hd__nand2_1
X_5027_ _2986_ _0729_ _1533_ vssd1 vssd1 vccd1 vccd1 _1534_ sky130_fd_sc_hd__o21ai_1
XFILLER_57_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5929_ _2400_ _2428_ vssd1 vssd1 vccd1 vccd1 _2429_ sky130_fd_sc_hd__nor2_1
XFILLER_5_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4260_ _3310_ _0772_ vssd1 vssd1 vccd1 vccd1 _0773_ sky130_fd_sc_hd__nand2_1
X_4191_ _0702_ _0546_ _0703_ vssd1 vssd1 vccd1 vccd1 _0704_ sky130_fd_sc_hd__o21ai_1
XFILLER_86_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6832_ net76 _0291_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BitStream_buffer_output\[9\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_62_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_0__2891_ _2891_ vssd1 vssd1 vccd1 vccd1 clknet_0__2891_ sky130_fd_sc_hd__clkbuf_16
X_3975_ _0488_ _3046_ vssd1 vssd1 vccd1 vccd1 _0489_ sky130_fd_sc_hd__nor2_2
X_6763_ net167 _0222_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[57\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_10_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5714_ _0469_ egd_top.BitStream_buffer.BS_buffer\[73\] vssd1 vssd1 vccd1 vccd1 _2215_
+ sky130_fd_sc_hd__nand2_1
XFILLER_40_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5645_ _3311_ _3251_ _0772_ _3255_ _2146_ vssd1 vssd1 vccd1 vccd1 _2147_ sky130_fd_sc_hd__a221oi_1
XFILLER_40_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5576_ _0443_ _0378_ _0655_ _0382_ _2077_ vssd1 vssd1 vccd1 vccd1 _2078_ sky130_fd_sc_hd__a221oi_1
X_4527_ _3164_ _3078_ _3153_ _3080_ _1037_ vssd1 vssd1 vccd1 vccd1 _1038_ sky130_fd_sc_hd__a221oi_2
X_4458_ _0965_ _0438_ _0966_ _0967_ _0968_ vssd1 vssd1 vccd1 vccd1 _0969_ sky130_fd_sc_hd__o2111a_1
X_3409_ _2954_ _2919_ vssd1 vssd1 vccd1 vccd1 _2961_ sky130_fd_sc_hd__or2b_1
X_4389_ _0511_ vssd1 vssd1 vccd1 vccd1 _0901_ sky130_fd_sc_hd__inv_2
XFILLER_58_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6128_ _2538_ _1149_ vssd1 vssd1 vccd1 vccd1 _2548_ sky130_fd_sc_hd__nand2_1
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6059_ _3023_ _2489_ _2501_ _2507_ vssd1 vssd1 vccd1 vccd1 _0232_ sky130_fd_sc_hd__o211a_1
XFILLER_14_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_367 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6645__21 clknet_1_0__leaf__2894_ vssd1 vssd1 vccd1 vccd1 net55 sky130_fd_sc_hd__inv_2
XFILLER_49_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3760_ _3290_ _3059_ vssd1 vssd1 vccd1 vccd1 _3294_ sky130_fd_sc_hd__nor2_2
XFILLER_20_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5430_ _3173_ _3156_ _3177_ _3160_ _1933_ vssd1 vssd1 vccd1 vccd1 _1934_ sky130_fd_sc_hd__a221oi_1
X_3691_ _3087_ _3213_ vssd1 vssd1 vccd1 vccd1 _3225_ sky130_fd_sc_hd__nand2_1
XFILLER_65_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5361_ _0548_ _0354_ vssd1 vssd1 vccd1 vccd1 _1865_ sky130_fd_sc_hd__nand2_1
X_4312_ _0744_ _3194_ _3197_ _3149_ _0823_ vssd1 vssd1 vccd1 vccd1 _0824_ sky130_fd_sc_hd__a221oi_1
X_5292_ _1783_ _1796_ vssd1 vssd1 vccd1 vccd1 _1797_ sky130_fd_sc_hd__nand2_1
X_4243_ _3216_ _3217_ vssd1 vssd1 vccd1 vccd1 _0756_ sky130_fd_sc_hd__nand2_1
X_4174_ _0606_ egd_top.BitStream_buffer.BS_buffer\[13\] vssd1 vssd1 vccd1 vccd1 _0687_
+ sky130_fd_sc_hd__nand2_1
XFILLER_67_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6815_ net59 _0274_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_6746_ net150 _0205_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[74\]
+ sky130_fd_sc_hd__dfxtp_2
X_3958_ _3071_ _2934_ vssd1 vssd1 vccd1 vccd1 _0472_ sky130_fd_sc_hd__nand2_2
XFILLER_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3889_ _0402_ vssd1 vssd1 vccd1 vccd1 _0403_ sky130_fd_sc_hd__buf_2
X_5628_ _2085_ _2100_ _2115_ _2129_ vssd1 vssd1 vccd1 vccd1 _2130_ sky130_fd_sc_hd__and4_1
X_5559_ _0606_ _0509_ vssd1 vssd1 vccd1 vccd1 _2062_ sky130_fd_sc_hd__nand2_1
XFILLER_58_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_511 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4930_ _3250_ egd_top.BitStream_buffer.BS_buffer\[80\] vssd1 vssd1 vccd1 vccd1 _1438_
+ sky130_fd_sc_hd__nand2_1
X_4861_ _0581_ egd_top.BitStream_buffer.BS_buffer\[16\] vssd1 vssd1 vccd1 vccd1 _1369_
+ sky130_fd_sc_hd__nand2_1
X_3812_ _0325_ vssd1 vssd1 vccd1 vccd1 _0326_ sky130_fd_sc_hd__inv_2
X_4792_ _1289_ _1293_ _1296_ _1300_ vssd1 vssd1 vccd1 vccd1 _1301_ sky130_fd_sc_hd__and4_1
XFILLER_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3743_ _3276_ vssd1 vssd1 vccd1 vccd1 _3277_ sky130_fd_sc_hd__clkinv_2
X_3674_ _3152_ _3172_ _3190_ _3207_ vssd1 vssd1 vccd1 vccd1 _3208_ sky130_fd_sc_hd__and4_1
XFILLER_9_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6462_ _2825_ _2789_ vssd1 vssd1 vccd1 vccd1 _2826_ sky130_fd_sc_hd__nand2_1
X_6571__113 clknet_1_0__leaf__2888_ vssd1 vssd1 vccd1 vccd1 net147 sky130_fd_sc_hd__inv_2
X_5413_ _3061_ _3070_ vssd1 vssd1 vccd1 vccd1 _1917_ sky130_fd_sc_hd__nand2_1
X_6393_ _2756_ _2762_ vssd1 vssd1 vccd1 vccd1 _2763_ sky130_fd_sc_hd__nor2_1
X_5344_ _3244_ _0432_ _0435_ _0751_ _1847_ vssd1 vssd1 vccd1 vccd1 _1848_ sky130_fd_sc_hd__a221oi_1
XFILLER_87_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5275_ _0477_ _3227_ vssd1 vssd1 vccd1 vccd1 _1780_ sky130_fd_sc_hd__nand2_1
X_4226_ _0737_ _0738_ vssd1 vssd1 vccd1 vccd1 _0739_ sky130_fd_sc_hd__nand2_1
XFILLER_87_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4157_ egd_top.BitStream_buffer.BS_buffer\[8\] vssd1 vssd1 vccd1 vccd1 _0670_ sky130_fd_sc_hd__inv_2
X_4088_ egd_top.BitStream_buffer.BS_buffer\[15\] vssd1 vssd1 vccd1 vccd1 _0602_ sky130_fd_sc_hd__clkinv_4
XFILLER_70_226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6729_ net133 _0188_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[107\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_3_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput14 la_data_in_58_43[7] vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__clkbuf_1
XFILLER_6_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3390_ egd_top.BitStream_buffer.buffer_index\[6\] egd_top.BitStream_buffer.buffer_index\[5\]
+ egd_top.BitStream_buffer.buffer_index\[4\] vssd1 vssd1 vccd1 vccd1 _2944_ sky130_fd_sc_hd__or3_1
XFILLER_69_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5060_ _1559_ _1563_ _1566_ vssd1 vssd1 vccd1 vccd1 _1567_ sky130_fd_sc_hd__nor3_1
XFILLER_77_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4011_ _0521_ _3057_ vssd1 vssd1 vccd1 vccd1 _0525_ sky130_fd_sc_hd__nand2_2
XFILLER_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f__2897_ clknet_0__2897_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__2897_
+ sky130_fd_sc_hd__clkbuf_16
X_5962_ _2449_ _0673_ vssd1 vssd1 vccd1 vccd1 _2452_ sky130_fd_sc_hd__nand2_1
XFILLER_37_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4913_ _1035_ _3122_ _1418_ _1419_ _1420_ vssd1 vssd1 vccd1 vccd1 _1421_ sky130_fd_sc_hd__o2111a_1
X_5893_ _0458_ _3256_ vssd1 vssd1 vccd1 vccd1 _2393_ sky130_fd_sc_hd__nand2_1
XFILLER_60_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4844_ _0452_ _0478_ vssd1 vssd1 vccd1 vccd1 _1352_ sky130_fd_sc_hd__nand2_1
X_4775_ _0960_ _0403_ _1283_ vssd1 vssd1 vccd1 vccd1 _1284_ sky130_fd_sc_hd__o21ai_1
X_6514_ _2858_ _2854_ _2855_ vssd1 vssd1 vccd1 vccd1 _2875_ sky130_fd_sc_hd__o21ai_1
XFILLER_20_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3726_ _3259_ vssd1 vssd1 vccd1 vccd1 _3260_ sky130_fd_sc_hd__inv_2
X_3657_ egd_top.BitStream_buffer.BS_buffer\[118\] vssd1 vssd1 vccd1 vccd1 _3191_ sky130_fd_sc_hd__clkbuf_4
X_6445_ _2808_ _2804_ vssd1 vssd1 vccd1 vccd1 _2809_ sky130_fd_sc_hd__nand2_1
X_3588_ _3121_ _3036_ vssd1 vssd1 vccd1 vccd1 _3122_ sky130_fd_sc_hd__nand2_2
X_6376_ _2742_ _2745_ vssd1 vssd1 vccd1 vccd1 _2746_ sky130_fd_sc_hd__nand2_1
X_5327_ _0383_ _0368_ _1830_ vssd1 vssd1 vccd1 vccd1 _1831_ sky130_fd_sc_hd__o21ai_1
XFILLER_57_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5258_ _1761_ _1762_ vssd1 vssd1 vccd1 vccd1 _1763_ sky130_fd_sc_hd__nand2_1
X_5189_ _0679_ _0593_ _0574_ _0599_ _1694_ vssd1 vssd1 vccd1 vccd1 _1695_ sky130_fd_sc_hd__o221a_1
X_4209_ egd_top.BitStream_buffer.BS_buffer\[105\] vssd1 vssd1 vccd1 vccd1 _0722_ sky130_fd_sc_hd__clkbuf_4
XFILLER_28_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4560_ _3185_ _0930_ vssd1 vssd1 vccd1 vccd1 _1071_ sky130_fd_sc_hd__nand2_1
XFILLER_8_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3511_ _3044_ vssd1 vssd1 vccd1 vccd1 _3045_ sky130_fd_sc_hd__buf_6
X_4491_ _0952_ _0970_ _0985_ _1001_ vssd1 vssd1 vccd1 vccd1 _1002_ sky130_fd_sc_hd__and4_1
X_3442_ net3 vssd1 vssd1 vccd1 vccd1 _2988_ sky130_fd_sc_hd__buf_4
X_6230_ _2904_ vssd1 vssd1 vccd1 vccd1 _2611_ sky130_fd_sc_hd__buf_2
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3373_ egd_top.BitStream_buffer.pc_previous\[0\] vssd1 vssd1 vccd1 vccd1 _2927_ sky130_fd_sc_hd__inv_2
X_6161_ _3005_ _2554_ _2558_ _2567_ vssd1 vssd1 vccd1 vccd1 _0190_ sky130_fd_sc_hd__o211a_1
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5112_ _3288_ _3251_ _3255_ _3293_ vssd1 vssd1 vccd1 vccd1 _1618_ sky130_fd_sc_hd__a22o_1
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6092_ _2517_ _0887_ vssd1 vssd1 vccd1 vccd1 _2527_ sky130_fd_sc_hd__nand2_1
X_5043_ _1539_ _1543_ _1546_ _1549_ vssd1 vssd1 vccd1 vccd1 _1550_ sky130_fd_sc_hd__and4_1
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5945_ _2440_ vssd1 vssd1 vccd1 vccd1 _2441_ sky130_fd_sc_hd__clkbuf_2
XFILLER_80_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5876_ _0388_ _0454_ vssd1 vssd1 vccd1 vccd1 _2376_ sky130_fd_sc_hd__nand2_1
X_4827_ egd_top.BitStream_buffer.BitStream_buffer_output\[9\] _2965_ _0627_ vssd1
+ vssd1 vccd1 vccd1 _1335_ sky130_fd_sc_hd__o21ai_1
X_4758_ _1263_ _1264_ _1265_ _1266_ vssd1 vssd1 vccd1 vccd1 _1267_ sky130_fd_sc_hd__and4_1
X_4689_ _0591_ _3183_ _1198_ vssd1 vssd1 vccd1 vccd1 _1199_ sky130_fd_sc_hd__o21ai_1
XFILLER_4_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3709_ _3242_ vssd1 vssd1 vccd1 vccd1 _3243_ sky130_fd_sc_hd__buf_6
X_6428_ _2791_ _2793_ _2792_ vssd1 vssd1 vccd1 vccd1 _2796_ sky130_fd_sc_hd__nand3_1
XFILLER_88_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6359_ _2663_ _2627_ _2681_ vssd1 vssd1 vccd1 vccd1 _2730_ sky130_fd_sc_hd__nand3_1
XFILLER_75_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3 egd_top.BitStream_buffer.buffer_index\[6\] vssd1 vssd1 vccd1 vccd1 net198 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_47_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3991_ egd_top.BitStream_buffer.BS_buffer\[21\] vssd1 vssd1 vccd1 vccd1 _0505_ sky130_fd_sc_hd__clkbuf_4
X_5730_ _0532_ _0612_ vssd1 vssd1 vccd1 vccd1 _2231_ sky130_fd_sc_hd__or2_1
XFILLER_22_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5661_ _0741_ _3156_ _3187_ _3160_ _2162_ vssd1 vssd1 vccd1 vccd1 _2163_ sky130_fd_sc_hd__a221oi_1
XFILLER_30_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4612_ _0673_ _0592_ _0569_ _0596_ _1121_ vssd1 vssd1 vccd1 vccd1 _1122_ sky130_fd_sc_hd__o221a_1
X_5592_ _0432_ _3230_ vssd1 vssd1 vccd1 vccd1 _2094_ sky130_fd_sc_hd__nand2_1
X_4543_ _0842_ _3279_ _1053_ vssd1 vssd1 vccd1 vccd1 _1054_ sky130_fd_sc_hd__o21ai_1
X_4474_ _0974_ _0978_ _0980_ _0984_ vssd1 vssd1 vccd1 vccd1 _0985_ sky130_fd_sc_hd__and4_1
X_6213_ _2967_ net196 _2971_ vssd1 vssd1 vccd1 vccd1 _2600_ sky130_fd_sc_hd__nor3_1
X_3425_ _2974_ vssd1 vssd1 vccd1 vccd1 _2975_ sky130_fd_sc_hd__buf_2
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3356_ _2906_ _2911_ vssd1 vssd1 vccd1 vccd1 _2912_ sky130_fd_sc_hd__nor2_1
X_6144_ _2904_ vssd1 vssd1 vccd1 vccd1 _2558_ sky130_fd_sc_hd__buf_2
XFILLER_85_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6075_ _2988_ _2510_ _2516_ _2518_ vssd1 vssd1 vccd1 vccd1 _0227_ sky130_fd_sc_hd__o211a_1
XFILLER_38_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5026_ _3074_ _3204_ vssd1 vssd1 vccd1 vccd1 _1533_ sky130_fd_sc_hd__nand2_1
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6609__148 clknet_1_1__leaf__2891_ vssd1 vssd1 vccd1 vccd1 net182 sky130_fd_sc_hd__inv_2
XFILLER_38_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_310 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5928_ _2412_ _2427_ vssd1 vssd1 vccd1 vccd1 _2428_ sky130_fd_sc_hd__nand2_1
XFILLER_13_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5859_ _3159_ _0792_ vssd1 vssd1 vccd1 vccd1 _2359_ sky130_fd_sc_hd__nand2_1
XFILLER_70_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_50 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4190_ _0548_ egd_top.BitStream_buffer.BS_buffer\[29\] vssd1 vssd1 vccd1 vccd1 _0703_
+ sky130_fd_sc_hd__nand2_1
XFILLER_5_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_90 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_438 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6831_ net75 _0290_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BitStream_buffer_output\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_23_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__2890_ _2890_ vssd1 vssd1 vccd1 vccd1 clknet_0__2890_ sky130_fd_sc_hd__clkbuf_16
XFILLER_35_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3974_ _0484_ vssd1 vssd1 vccd1 vccd1 _0488_ sky130_fd_sc_hd__clkinv_4
X_6762_ net166 _0221_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[58\]
+ sky130_fd_sc_hd__dfxtp_1
X_5713_ _1297_ _0438_ _2211_ _2212_ _2213_ vssd1 vssd1 vccd1 vccd1 _2214_ sky130_fd_sc_hd__o2111a_1
X_5644_ _1158_ _3260_ _2145_ vssd1 vssd1 vccd1 vccd1 _2146_ sky130_fd_sc_hd__o21ai_1
X_5575_ _0883_ _0385_ _2076_ vssd1 vssd1 vccd1 vccd1 _2077_ sky130_fd_sc_hd__o21ai_1
X_4526_ _1035_ _0728_ _1036_ vssd1 vssd1 vccd1 vccd1 _1037_ sky130_fd_sc_hd__o21ai_1
X_4457_ _0434_ _0459_ vssd1 vssd1 vccd1 vccd1 _0968_ sky130_fd_sc_hd__nand2_1
X_3408_ _2960_ vssd1 vssd1 vccd1 vccd1 _0316_ sky130_fd_sc_hd__inv_2
X_4388_ _0491_ _0487_ _0498_ _0490_ _0899_ vssd1 vssd1 vccd1 vccd1 _0900_ sky130_fd_sc_hd__a221oi_1
XFILLER_85_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6127_ _3011_ _2533_ _2543_ _2547_ vssd1 vssd1 vccd1 vccd1 _0204_ sky130_fd_sc_hd__o211a_1
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6058_ _2486_ _0401_ vssd1 vssd1 vccd1 vccd1 _2507_ sky130_fd_sc_hd__nand2_1
X_5009_ _0606_ _0498_ vssd1 vssd1 vccd1 vccd1 _1516_ sky130_fd_sc_hd__nand2_1
XFILLER_73_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_302 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3690_ _3223_ vssd1 vssd1 vccd1 vccd1 _3224_ sky130_fd_sc_hd__buf_6
X_5360_ _0531_ _0487_ egd_top.BitStream_buffer.BS_buffer\[27\] _0490_ _1863_ vssd1
+ vssd1 vccd1 vccd1 _1864_ sky130_fd_sc_hd__a221oi_1
XFILLER_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4311_ _2999_ _3200_ _0822_ vssd1 vssd1 vccd1 vccd1 _0823_ sky130_fd_sc_hd__o21ai_1
X_5291_ _1786_ _1789_ _1792_ _1795_ vssd1 vssd1 vccd1 vccd1 _1796_ sky130_fd_sc_hd__and4_1
X_4242_ egd_top.BitStream_buffer.BS_buffer\[70\] vssd1 vssd1 vccd1 vccd1 _0755_ sky130_fd_sc_hd__clkinv_2
X_4173_ _0609_ egd_top.BitStream_buffer.BS_buffer\[15\] vssd1 vssd1 vccd1 vccd1 _0686_
+ sky130_fd_sc_hd__nand2_1
XFILLER_55_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6814_ net58 _0273_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_35_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3957_ egd_top.BitStream_buffer.BS_buffer\[61\] vssd1 vssd1 vccd1 vccd1 _0471_ sky130_fd_sc_hd__clkbuf_4
X_6745_ net149 _0204_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[75\]
+ sky130_fd_sc_hd__dfxtp_1
X_3888_ _2931_ _0339_ vssd1 vssd1 vccd1 vccd1 _0402_ sky130_fd_sc_hd__nand2_2
X_5627_ _2119_ _2123_ _2126_ _2128_ vssd1 vssd1 vccd1 vccd1 _2129_ sky130_fd_sc_hd__and4_1
X_5558_ _0611_ _0593_ _0676_ _0596_ _2060_ vssd1 vssd1 vccd1 vccd1 _2061_ sky130_fd_sc_hd__o221a_1
X_4509_ _1006_ _1011_ _1015_ _1019_ vssd1 vssd1 vccd1 vccd1 _1020_ sky130_fd_sc_hd__and4_1
XFILLER_78_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5489_ _0772_ _3270_ _3334_ _3275_ _1991_ vssd1 vssd1 vccd1 vccd1 _1992_ sky130_fd_sc_hd__a221oi_1
XFILLER_76_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4860_ _0611_ _0557_ _1365_ _1366_ _1367_ vssd1 vssd1 vccd1 vccd1 _1368_ sky130_fd_sc_hd__o2111a_1
XFILLER_82_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3811_ _3290_ _3072_ vssd1 vssd1 vccd1 vccd1 _0325_ sky130_fd_sc_hd__nor2_1
XFILLER_32_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6539__84 clknet_1_1__leaf__2885_ vssd1 vssd1 vccd1 vccd1 net118 sky130_fd_sc_hd__inv_2
X_4791_ _3237_ _0477_ _3210_ _2936_ _1299_ vssd1 vssd1 vccd1 vccd1 _1300_ sky130_fd_sc_hd__a221oi_2
XFILLER_20_327 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3742_ egd_top.BitStream_buffer.BS_buffer\[79\] vssd1 vssd1 vccd1 vccd1 _3276_ sky130_fd_sc_hd__clkbuf_4
X_3673_ _3191_ _3194_ _3197_ _3198_ _3206_ vssd1 vssd1 vccd1 vccd1 _3207_ sky130_fd_sc_hd__a221oi_1
X_6461_ _2735_ _2764_ _2684_ vssd1 vssd1 vccd1 vccd1 _2825_ sky130_fd_sc_hd__o21ai_1
X_5412_ _3153_ _3127_ _1914_ _1915_ vssd1 vssd1 vccd1 vccd1 _1916_ sky130_fd_sc_hd__a211oi_1
X_6392_ _2759_ _2761_ vssd1 vssd1 vccd1 vccd1 _2762_ sky130_fd_sc_hd__nand2_1
X_6554__98 clknet_1_1__leaf__2886_ vssd1 vssd1 vccd1 vccd1 net132 sky130_fd_sc_hd__inv_2
X_5343_ _0474_ _0439_ _1846_ vssd1 vssd1 vccd1 vccd1 _1847_ sky130_fd_sc_hd__o21ai_1
XFILLER_87_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5274_ _1297_ _0464_ _1776_ _1777_ _1778_ vssd1 vssd1 vccd1 vccd1 _1779_ sky130_fd_sc_hd__o2111a_1
X_4225_ _3168_ _3164_ vssd1 vssd1 vccd1 vccd1 _0738_ sky130_fd_sc_hd__nand2_1
X_4156_ _0646_ _0668_ vssd1 vssd1 vccd1 vccd1 _0669_ sky130_fd_sc_hd__and2_1
XFILLER_55_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_427 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4087_ _0591_ _0593_ _0594_ _0596_ _0600_ vssd1 vssd1 vccd1 vccd1 _0601_ sky130_fd_sc_hd__o221a_1
XFILLER_70_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4989_ egd_top.BitStream_buffer.BS_buffer\[29\] _0514_ _0537_ _0901_ _1495_ vssd1
+ vssd1 vccd1 vccd1 _1496_ sky130_fd_sc_hd__a221oi_1
XFILLER_11_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6728_ net132 _0187_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[108\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_11_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_500 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_50 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput15 la_data_in_58_43[8] vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__clkbuf_1
XFILLER_10_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4010_ egd_top.BitStream_buffer.BS_buffer\[27\] vssd1 vssd1 vccd1 vccd1 _0524_ sky130_fd_sc_hd__inv_2
XFILLER_77_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0__f__2896_ clknet_0__2896_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__2896_
+ sky130_fd_sc_hd__clkbuf_16
X_5961_ _2992_ _2442_ _2446_ _2451_ vssd1 vssd1 vccd1 vccd1 _0274_ sky130_fd_sc_hd__o211a_1
XFILLER_37_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4912_ _3116_ _3164_ vssd1 vssd1 vccd1 vccd1 _1420_ sky130_fd_sc_hd__nand2_1
XFILLER_52_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5892_ _0453_ _3221_ vssd1 vssd1 vccd1 vccd1 _2392_ sky130_fd_sc_hd__nand2_1
X_4843_ _0454_ _0415_ _0461_ _0419_ _1350_ vssd1 vssd1 vccd1 vccd1 _1351_ sky130_fd_sc_hd__a221oi_1
XFILLER_20_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4774_ _0406_ _0416_ vssd1 vssd1 vccd1 vccd1 _1283_ sky130_fd_sc_hd__nand2_1
X_3725_ _3258_ vssd1 vssd1 vccd1 vccd1 _3259_ sky130_fd_sc_hd__buf_2
X_6513_ _2873_ _2874_ vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__nand2_1
X_6444_ _2807_ _2771_ vssd1 vssd1 vccd1 vccd1 _2808_ sky130_fd_sc_hd__nand2_1
X_3656_ _3173_ _3176_ _3177_ _3180_ _3189_ vssd1 vssd1 vccd1 vccd1 _3190_ sky130_fd_sc_hd__a221oi_1
X_3587_ _3120_ vssd1 vssd1 vccd1 vccd1 _3121_ sky130_fd_sc_hd__buf_6
X_6375_ _2743_ _2744_ vssd1 vssd1 vccd1 vccd1 _2745_ sky130_fd_sc_hd__nand2_1
X_5326_ _0371_ _0389_ vssd1 vssd1 vccd1 vccd1 _1830_ sky130_fd_sc_hd__nand2_1
XFILLER_87_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5257_ _3167_ _3149_ vssd1 vssd1 vccd1 vccd1 _1762_ sky130_fd_sc_hd__nand2_1
X_4208_ egd_top.BitStream_buffer.BS_buffer\[106\] vssd1 vssd1 vccd1 vccd1 _0721_ sky130_fd_sc_hd__clkinv_2
X_5188_ _0586_ _0595_ vssd1 vssd1 vccd1 vccd1 _1694_ sky130_fd_sc_hd__or2_1
XFILLER_56_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4139_ _0647_ _0449_ _0648_ _0649_ _0651_ vssd1 vssd1 vccd1 vccd1 _0652_ sky130_fd_sc_hd__o2111a_1
XFILLER_83_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6533__79 clknet_1_1__leaf__2884_ vssd1 vssd1 vccd1 vccd1 net113 sky130_fd_sc_hd__inv_2
XFILLER_3_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3510_ _3043_ _3031_ _3032_ vssd1 vssd1 vccd1 vccd1 _3044_ sky130_fd_sc_hd__and3_1
X_4490_ _0990_ _0994_ _0998_ _1000_ vssd1 vssd1 vccd1 vccd1 _1001_ sky130_fd_sc_hd__and4_1
XFILLER_6_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3441_ _2985_ _2975_ _2913_ _2987_ vssd1 vssd1 vccd1 vccd1 _0310_ sky130_fd_sc_hd__o211a_1
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3372_ net18 net17 vssd1 vssd1 vccd1 vccd1 _2926_ sky130_fd_sc_hd__nor2_4
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6160_ _2561_ _3119_ vssd1 vssd1 vccd1 vccd1 _2567_ sky130_fd_sc_hd__nand2_1
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5111_ _1601_ _1616_ vssd1 vssd1 vccd1 vccd1 _1617_ sky130_fd_sc_hd__nand2_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6091_ _3014_ _2511_ _2516_ _2526_ vssd1 vssd1 vccd1 vccd1 _0219_ sky130_fd_sc_hd__o211a_1
X_6693__64 clknet_1_0__leaf__2899_ vssd1 vssd1 vccd1 vccd1 net98 sky130_fd_sc_hd__inv_2
X_5042_ _1076_ _3176_ _0566_ _3180_ _1548_ vssd1 vssd1 vccd1 vccd1 _1549_ sky130_fd_sc_hd__a221oi_2
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5944_ _2944_ _2437_ vssd1 vssd1 vccd1 vccd1 _2440_ sky130_fd_sc_hd__or2_1
X_5875_ _0412_ _0342_ _0345_ _0416_ _2374_ vssd1 vssd1 vccd1 vccd1 _2375_ sky130_fd_sc_hd__a221oi_1
X_4826_ _1207_ _1334_ vssd1 vssd1 vccd1 vccd1 _0292_ sky130_fd_sc_hd__nor2_1
X_4757_ _3259_ egd_top.BitStream_buffer.BS_buffer\[77\] vssd1 vssd1 vccd1 vccd1 _1266_
+ sky130_fd_sc_hd__nand2_1
X_4688_ _3186_ _1076_ vssd1 vssd1 vccd1 vccd1 _1198_ sky130_fd_sc_hd__nand2_1
X_3708_ _3241_ vssd1 vssd1 vccd1 vccd1 _3242_ sky130_fd_sc_hd__clkbuf_2
X_3639_ egd_top.BitStream_buffer.BS_buffer\[124\] vssd1 vssd1 vccd1 vccd1 _3173_ sky130_fd_sc_hd__clkbuf_4
X_6427_ net22 _2794_ vssd1 vssd1 vccd1 vccd1 _2795_ sky130_fd_sc_hd__nand2_1
X_6358_ _2727_ _2728_ vssd1 vssd1 vccd1 vccd1 _2729_ sky130_fd_sc_hd__nand2_1
XFILLER_88_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5309_ _0578_ egd_top.BitStream_buffer.BS_buffer\[17\] vssd1 vssd1 vccd1 vccd1 _1814_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6289_ _2644_ _2659_ vssd1 vssd1 vccd1 vccd1 _2660_ sky130_fd_sc_hd__nand2_1
XFILLER_84_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3990_ _0503_ vssd1 vssd1 vccd1 vccd1 _0504_ sky130_fd_sc_hd__clkbuf_4
XFILLER_50_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5660_ _2160_ _2161_ vssd1 vssd1 vccd1 vccd1 _2162_ sky130_fd_sc_hd__nand2_1
XFILLER_15_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4611_ _0554_ _0598_ vssd1 vssd1 vccd1 vccd1 _1121_ sky130_fd_sc_hd__or2_1
X_5591_ _0441_ _3244_ vssd1 vssd1 vccd1 vccd1 _2093_ sky130_fd_sc_hd__nand2_1
X_4542_ _3281_ _3302_ vssd1 vssd1 vccd1 vccd1 _1053_ sky130_fd_sc_hd__nand2_1
X_4473_ _0492_ _0603_ _0981_ _0982_ _0983_ vssd1 vssd1 vccd1 vccd1 _0984_ sky130_fd_sc_hd__o2111a_1
XFILLER_7_470 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3424_ _2973_ vssd1 vssd1 vccd1 vccd1 _2974_ sky130_fd_sc_hd__clkinv_2
X_6212_ _2599_ vssd1 vssd1 vccd1 vccd1 _0177_ sky130_fd_sc_hd__inv_2
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3355_ _2903_ _2910_ vssd1 vssd1 vccd1 vccd1 _2911_ sky130_fd_sc_hd__nor2_1
X_6143_ _2979_ _2554_ _2543_ _2557_ vssd1 vssd1 vccd1 vccd1 _0198_ sky130_fd_sc_hd__o211a_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6074_ _2517_ _0960_ vssd1 vssd1 vccd1 vccd1 _2518_ sky130_fd_sc_hd__nand2_1
X_5025_ _3164_ _3113_ _3117_ _3153_ _1531_ vssd1 vssd1 vccd1 vccd1 _1532_ sky130_fd_sc_hd__a221oi_1
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5927_ _2416_ _2420_ _2422_ _2426_ vssd1 vssd1 vccd1 vccd1 _2427_ sky130_fd_sc_hd__and4_1
XFILLER_53_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5858_ _3162_ _3187_ vssd1 vssd1 vccd1 vccd1 _2358_ sky130_fd_sc_hd__nand2_1
X_4809_ _0676_ _0558_ _1315_ _1316_ _1317_ vssd1 vssd1 vccd1 vccd1 _1318_ sky130_fd_sc_hd__o2111a_1
X_5789_ _3301_ _3338_ vssd1 vssd1 vccd1 vccd1 _2290_ sky130_fd_sc_hd__nand2_1
XFILLER_79_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6672__45 clknet_1_0__leaf__2897_ vssd1 vssd1 vccd1 vccd1 net79 sky130_fd_sc_hd__inv_2
XFILLER_29_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_62 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6830_ net74 _0289_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BitStream_buffer_output\[7\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_90_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6761_ net165 _0220_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[59\]
+ sky130_fd_sc_hd__dfxtp_1
X_3973_ _0486_ vssd1 vssd1 vccd1 vccd1 _0487_ sky130_fd_sc_hd__buf_2
X_5712_ _0434_ _3210_ vssd1 vssd1 vccd1 vccd1 _2213_ sky130_fd_sc_hd__nand2_1
XFILLER_50_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5643_ _3263_ _0774_ vssd1 vssd1 vccd1 vccd1 _2145_ sky130_fd_sc_hd__nand2_1
X_5574_ _0387_ _0429_ vssd1 vssd1 vccd1 vccd1 _2076_ sky130_fd_sc_hd__nand2_1
X_4525_ _3073_ _3169_ vssd1 vssd1 vccd1 vccd1 _1036_ sky130_fd_sc_hd__nand2_1
X_6615__153 clknet_1_0__leaf__2892_ vssd1 vssd1 vccd1 vccd1 net187 sky130_fd_sc_hd__inv_2
X_4456_ _0441_ _0436_ vssd1 vssd1 vccd1 vccd1 _0967_ sky130_fd_sc_hd__nand2_1
X_4387_ _0897_ _0495_ _0898_ vssd1 vssd1 vccd1 vccd1 _0899_ sky130_fd_sc_hd__o21ai_1
X_3407_ net29 _2951_ _2902_ _2959_ vssd1 vssd1 vccd1 vccd1 _2960_ sky130_fd_sc_hd__o211ai_1
X_6126_ _2538_ _1144_ vssd1 vssd1 vccd1 vccd1 _2547_ sky130_fd_sc_hd__nand2_1
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6057_ _3020_ _2489_ _2501_ _2506_ vssd1 vssd1 vccd1 vccd1 _0233_ sky130_fd_sc_hd__o211a_1
X_5008_ _0586_ _0593_ _0679_ _0599_ _1514_ vssd1 vssd1 vccd1 vccd1 _1515_ sky130_fd_sc_hd__o221a_1
XFILLER_26_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_62 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4310_ _3203_ _3191_ vssd1 vssd1 vccd1 vccd1 _0822_ sky130_fd_sc_hd__nand2_1
X_5290_ _0655_ _0396_ _0399_ _0429_ _1794_ vssd1 vssd1 vccd1 vccd1 _1795_ sky130_fd_sc_hd__a221oi_1
X_4241_ _3237_ _3233_ _3210_ _3236_ _0753_ vssd1 vssd1 vccd1 vccd1 _0754_ sky130_fd_sc_hd__a221oi_1
X_6636__12 clknet_1_0__leaf__2894_ vssd1 vssd1 vccd1 vccd1 net46 sky130_fd_sc_hd__inv_2
X_4172_ egd_top.BitStream_buffer.BS_buffer\[16\] vssd1 vssd1 vccd1 vccd1 _0685_ sky130_fd_sc_hd__inv_2
XFILLER_55_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6651__26 clknet_1_0__leaf__2895_ vssd1 vssd1 vccd1 vccd1 net60 sky130_fd_sc_hd__inv_2
X_6813_ net57 _0272_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_3956_ _0469_ vssd1 vssd1 vccd1 vccd1 _0470_ sky130_fd_sc_hd__buf_2
X_6744_ net148 _0203_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[76\]
+ sky130_fd_sc_hd__dfxtp_1
X_5626_ _0940_ _0522_ _1276_ _0533_ _2127_ vssd1 vssd1 vccd1 vccd1 _2128_ sky130_fd_sc_hd__o221a_1
XFILLER_31_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3887_ egd_top.BitStream_buffer.BS_buffer\[47\] vssd1 vssd1 vccd1 vccd1 _0401_ sky130_fd_sc_hd__clkinv_2
X_5557_ _0688_ _0599_ vssd1 vssd1 vccd1 vccd1 _2060_ sky130_fd_sc_hd__or2_1
X_4508_ _3040_ _3339_ _0708_ _0322_ _1018_ vssd1 vssd1 vccd1 vccd1 _1019_ sky130_fd_sc_hd__a221oi_1
XFILLER_2_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5488_ _0779_ _3279_ _1990_ vssd1 vssd1 vccd1 vccd1 _1991_ sky130_fd_sc_hd__o21ai_1
XFILLER_4_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4439_ _0659_ _0403_ _0949_ vssd1 vssd1 vccd1 vccd1 _0950_ sky130_fd_sc_hd__o21ai_1
XFILLER_86_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6109_ _2985_ _2532_ _2528_ _2537_ vssd1 vssd1 vccd1 vccd1 _0212_ sky130_fd_sc_hd__o211a_1
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_391 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4790_ _1297_ _0472_ _1298_ vssd1 vssd1 vccd1 vccd1 _1299_ sky130_fd_sc_hd__o21ai_1
X_3810_ egd_top.BitStream_buffer.BS_buffer\[93\] vssd1 vssd1 vccd1 vccd1 _0324_ sky130_fd_sc_hd__clkinv_2
XFILLER_60_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_339 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3741_ _3274_ vssd1 vssd1 vccd1 vccd1 _3275_ sky130_fd_sc_hd__clkbuf_4
XFILLER_13_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3672_ _2993_ _3200_ _3205_ vssd1 vssd1 vccd1 vccd1 _3206_ sky130_fd_sc_hd__o21ai_1
XFILLER_70_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6460_ _2823_ vssd1 vssd1 vccd1 vccd1 _2824_ sky130_fd_sc_hd__inv_2
X_5411_ _3204_ _3112_ _3116_ _0746_ vssd1 vssd1 vccd1 vccd1 _1915_ sky130_fd_sc_hd__a22o_1
X_6391_ _2632_ _2760_ _2660_ vssd1 vssd1 vccd1 vccd1 _2761_ sky130_fd_sc_hd__a21o_1
X_5342_ _0442_ _0478_ vssd1 vssd1 vccd1 vccd1 _1846_ sky130_fd_sc_hd__nand2_1
X_5273_ _1043_ _0449_ vssd1 vssd1 vccd1 vccd1 _1778_ sky130_fd_sc_hd__or2_1
X_4224_ _3163_ _3153_ vssd1 vssd1 vccd1 vccd1 _0737_ sky130_fd_sc_hd__nand2_1
XFILLER_68_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4155_ _0652_ _0658_ _0662_ _0667_ vssd1 vssd1 vccd1 vccd1 _0668_ sky130_fd_sc_hd__and4_1
XFILLER_55_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4086_ _0597_ _0599_ vssd1 vssd1 vccd1 vccd1 _0600_ sky130_fd_sc_hd__or2_1
XFILLER_70_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4988_ egd_top.BitStream_buffer.BS_buffer\[27\] _0503_ _0508_ egd_top.BitStream_buffer.BS_buffer\[28\]
+ vssd1 vssd1 vccd1 vccd1 _1495_ sky130_fd_sc_hd__a22o_1
XFILLER_23_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3939_ _0452_ vssd1 vssd1 vccd1 vccd1 _0453_ sky130_fd_sc_hd__clkbuf_4
X_6727_ net131 _0186_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[109\]
+ sky130_fd_sc_hd__dfxtp_1
X_5609_ _0608_ _0531_ vssd1 vssd1 vccd1 vccd1 _2111_ sky130_fd_sc_hd__nand2_1
XFILLER_11_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6699__70 clknet_1_1__leaf__2899_ vssd1 vssd1 vccd1 vccd1 net104 sky130_fd_sc_hd__inv_2
XFILLER_87_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput16 la_data_in_58_43[9] vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__clkbuf_1
XFILLER_10_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_504 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f__2895_ clknet_0__2895_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__2895_
+ sky130_fd_sc_hd__clkbuf_16
X_5960_ _2449_ _0569_ vssd1 vssd1 vccd1 vccd1 _2451_ sky130_fd_sc_hd__nand2_1
X_4911_ _3112_ _3169_ vssd1 vssd1 vccd1 vccd1 _1419_ sky130_fd_sc_hd__nand2_1
X_5891_ _3210_ _0432_ _0435_ _3217_ _2390_ vssd1 vssd1 vccd1 vccd1 _2391_ sky130_fd_sc_hd__a221oi_1
XFILLER_33_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4842_ _0883_ _0422_ _1349_ vssd1 vssd1 vccd1 vccd1 _1350_ sky130_fd_sc_hd__o21ai_1
X_4773_ _0400_ _0378_ _0407_ _0382_ _1281_ vssd1 vssd1 vccd1 vccd1 _1282_ sky130_fd_sc_hd__a221oi_1
X_3724_ _3124_ _3212_ vssd1 vssd1 vccd1 vccd1 _3258_ sky130_fd_sc_hd__and2_1
X_6512_ _2833_ _2846_ vssd1 vssd1 vccd1 vccd1 _2874_ sky130_fd_sc_hd__nand2_1
X_3655_ _3021_ _3183_ _3188_ vssd1 vssd1 vccd1 vccd1 _3189_ sky130_fd_sc_hd__o21ai_1
X_6443_ _2748_ _2773_ vssd1 vssd1 vccd1 vccd1 _2807_ sky130_fd_sc_hd__nor2_1
X_3586_ _3043_ _3031_ egd_top.BitStream_buffer.pc\[3\] vssd1 vssd1 vccd1 vccd1 _3120_
+ sky130_fd_sc_hd__and3_1
X_6374_ _2678_ _1945_ vssd1 vssd1 vccd1 vccd1 _2744_ sky130_fd_sc_hd__nand2_1
X_5325_ _1707_ _1829_ vssd1 vssd1 vccd1 vccd1 _0288_ sky130_fd_sc_hd__nor2_1
XFILLER_87_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5256_ _3162_ _3133_ vssd1 vssd1 vccd1 vccd1 _1761_ sky130_fd_sc_hd__nand2_1
XFILLER_87_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4207_ _0713_ _3106_ _0715_ _0717_ _0719_ vssd1 vssd1 vccd1 vccd1 _0720_ sky130_fd_sc_hd__o2111a_1
X_5187_ _0692_ _0576_ _1690_ _1691_ _1692_ vssd1 vssd1 vccd1 vccd1 _1693_ sky130_fd_sc_hd__o2111a_1
XFILLER_68_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4138_ _0650_ _0463_ vssd1 vssd1 vccd1 vccd1 _0651_ sky130_fd_sc_hd__or2_1
XFILLER_83_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_515 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4069_ egd_top.BitStream_buffer.BS_buffer\[10\] vssd1 vssd1 vccd1 vccd1 _0583_ sky130_fd_sc_hd__clkbuf_4
XFILLER_71_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_114 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3440_ _2976_ _2986_ vssd1 vssd1 vccd1 vccd1 _2987_ sky130_fd_sc_hd__nand2_1
X_3371_ _2924_ egd_top.BitStream_buffer.pc_previous\[0\] vssd1 vssd1 vccd1 vccd1 _2925_
+ sky130_fd_sc_hd__nand2_2
X_6678__51 clknet_1_1__leaf__2897_ vssd1 vssd1 vccd1 vccd1 net85 sky130_fd_sc_hd__inv_2
X_5110_ _1605_ _1609_ _1612_ _1615_ vssd1 vssd1 vccd1 vccd1 _1616_ sky130_fd_sc_hd__and4_1
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6090_ _2517_ _0647_ vssd1 vssd1 vccd1 vccd1 _2526_ sky130_fd_sc_hd__nand2_1
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5041_ _0569_ _3183_ _1547_ vssd1 vssd1 vccd1 vccd1 _1548_ sky130_fd_sc_hd__o21ai_1
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5943_ _2439_ vssd1 vssd1 vccd1 vccd1 _0280_ sky130_fd_sc_hd__clkbuf_1
XFILLER_18_291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5874_ _0437_ _0350_ _2373_ vssd1 vssd1 vccd1 vccd1 _2374_ sky130_fd_sc_hd__o21ai_1
X_4825_ _3026_ _1333_ vssd1 vssd1 vccd1 vccd1 _1334_ sky130_fd_sc_hd__nor2_1
XFILLER_21_467 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4756_ _3250_ egd_top.BitStream_buffer.BS_buffer\[79\] vssd1 vssd1 vccd1 vccd1 _1265_
+ sky130_fd_sc_hd__nand2_1
X_4687_ _3133_ _3194_ _3197_ _3138_ _1196_ vssd1 vssd1 vccd1 vccd1 _1197_ sky130_fd_sc_hd__a221oi_1
X_3707_ _3033_ _3212_ vssd1 vssd1 vccd1 vccd1 _3241_ sky130_fd_sc_hd__and2_1
X_3638_ _3153_ _3156_ _3157_ _3160_ _3171_ vssd1 vssd1 vccd1 vccd1 _3172_ sky130_fd_sc_hd__a221oi_1
X_6426_ _2793_ vssd1 vssd1 vccd1 vccd1 _2794_ sky130_fd_sc_hd__inv_2
X_3569_ _3043_ egd_top.BitStream_buffer.pc\[2\] _3032_ vssd1 vssd1 vccd1 vccd1 _3103_
+ sky130_fd_sc_hd__and3_1
XFILLER_68_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6357_ _2678_ egd_top.BitStream_buffer.BitStream_buffer_output\[3\] vssd1 vssd1 vccd1
+ vccd1 _2728_ sky130_fd_sc_hd__nand2_1
X_5308_ _0685_ _0558_ _1810_ _1811_ _1812_ vssd1 vssd1 vccd1 vccd1 _1813_ sky130_fd_sc_hd__o2111a_1
X_6288_ _2658_ _2623_ vssd1 vssd1 vccd1 vccd1 _2659_ sky130_fd_sc_hd__nand2_2
X_6584__125 clknet_1_1__leaf__2889_ vssd1 vssd1 vccd1 vccd1 net159 sky130_fd_sc_hd__inv_2
X_5239_ _3235_ _3268_ vssd1 vssd1 vccd1 vccd1 _1744_ sky130_fd_sc_hd__nand2_1
XFILLER_48_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4610_ _0602_ _0576_ _1117_ _1118_ _1119_ vssd1 vssd1 vccd1 vccd1 _1120_ sky130_fd_sc_hd__o2111a_1
XFILLER_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5590_ _1430_ _0450_ _2089_ _2090_ _2091_ vssd1 vssd1 vccd1 vccd1 _2092_ sky130_fd_sc_hd__o2111a_1
XFILLER_30_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4541_ _1048_ _1049_ _1050_ _1051_ vssd1 vssd1 vccd1 vccd1 _1052_ sky130_fd_sc_hd__and4_1
X_4472_ _0685_ _0612_ vssd1 vssd1 vccd1 vccd1 _0983_ sky130_fd_sc_hd__or2_1
X_3423_ _2967_ _2972_ vssd1 vssd1 vccd1 vccd1 _2973_ sky130_fd_sc_hd__nor2_1
X_6211_ _2905_ _2929_ vssd1 vssd1 vccd1 vccd1 _2599_ sky130_fd_sc_hd__or2_1
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6142_ _2555_ _1169_ vssd1 vssd1 vccd1 vccd1 _2557_ sky130_fd_sc_hd__nand2_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3354_ net33 net32 vssd1 vssd1 vccd1 vccd1 _2910_ sky130_fd_sc_hd__nor2_1
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6073_ _2509_ vssd1 vssd1 vccd1 vccd1 _2517_ sky130_fd_sc_hd__buf_2
X_5024_ _2977_ _3123_ _1530_ vssd1 vssd1 vccd1 vccd1 _1531_ sky130_fd_sc_hd__o21ai_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_504 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5926_ _0543_ _0604_ _2423_ _2424_ _2425_ vssd1 vssd1 vccd1 vccd1 _2426_ sky130_fd_sc_hd__o2111a_1
XFILLER_53_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5857_ _0566_ _3193_ _3196_ _0568_ _2356_ vssd1 vssd1 vccd1 vccd1 _2357_ sky130_fd_sc_hd__a221oi_1
XFILLER_70_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4808_ _0679_ _0571_ vssd1 vssd1 vccd1 vccd1 _1317_ sky130_fd_sc_hd__or2_1
X_5788_ _2279_ _2282_ _2285_ _2288_ vssd1 vssd1 vccd1 vccd1 _2289_ sky130_fd_sc_hd__and4_1
XFILLER_21_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4739_ _3163_ _3191_ vssd1 vssd1 vccd1 vccd1 _1248_ sky130_fd_sc_hd__nand2_1
XFILLER_79_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6409_ _2775_ _2777_ vssd1 vssd1 vccd1 vccd1 _2778_ sky130_fd_sc_hd__nand2_1
XFILLER_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6760_ net164 _0219_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[60\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_35_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3972_ _0485_ vssd1 vssd1 vccd1 vccd1 _0486_ sky130_fd_sc_hd__clkbuf_2
XFILLER_62_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5711_ _0442_ _0751_ vssd1 vssd1 vccd1 vccd1 _2212_ sky130_fd_sc_hd__nand2_1
XFILLER_50_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5642_ _2133_ _2137_ _2140_ _2143_ vssd1 vssd1 vccd1 vccd1 _2144_ sky130_fd_sc_hd__and4_1
X_5573_ _0407_ _0360_ _0363_ _0642_ _2074_ vssd1 vssd1 vccd1 vccd1 _2075_ sky130_fd_sc_hd__a221oi_2
X_4524_ egd_top.BitStream_buffer.BS_buffer\[111\] vssd1 vssd1 vccd1 vccd1 _1035_ sky130_fd_sc_hd__inv_2
XFILLER_7_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4455_ _0431_ _0461_ vssd1 vssd1 vccd1 vccd1 _0966_ sky130_fd_sc_hd__nand2_1
X_4386_ _0497_ _0505_ vssd1 vssd1 vccd1 vccd1 _0898_ sky130_fd_sc_hd__nand2_1
X_3406_ _2915_ _2958_ _2951_ vssd1 vssd1 vccd1 vccd1 _2959_ sky130_fd_sc_hd__o21ai_1
X_6125_ _3008_ _2533_ _2543_ _2546_ vssd1 vssd1 vccd1 vccd1 _0205_ sky130_fd_sc_hd__o211a_1
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6056_ _2486_ _1466_ vssd1 vssd1 vccd1 vccd1 _2506_ sky130_fd_sc_hd__nand2_1
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5007_ _0670_ _0596_ vssd1 vssd1 vccd1 vccd1 _1514_ sky130_fd_sc_hd__or2_1
XFILLER_53_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5909_ _0548_ _0389_ vssd1 vssd1 vccd1 vccd1 _2409_ sky130_fd_sc_hd__nand2_1
XFILLER_14_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4240_ _0751_ _3243_ _0752_ _3230_ vssd1 vssd1 vccd1 vccd1 _0753_ sky130_fd_sc_hd__a22o_1
X_4171_ _0597_ _0593_ _0682_ _0599_ _0683_ vssd1 vssd1 vccd1 vccd1 _0684_ sky130_fd_sc_hd__o221a_1
XFILLER_67_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6812_ net56 _0271_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_23_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6743_ net147 _0202_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[77\]
+ sky130_fd_sc_hd__dfxtp_1
X_3955_ _0468_ vssd1 vssd1 vccd1 vccd1 _0469_ sky130_fd_sc_hd__clkinv_2
X_5625_ _1084_ _0529_ _0348_ _0525_ vssd1 vssd1 vccd1 vccd1 _2127_ sky130_fd_sc_hd__o22a_1
X_3886_ egd_top.BitStream_buffer.BS_buffer\[45\] vssd1 vssd1 vccd1 vccd1 _0400_ sky130_fd_sc_hd__clkbuf_4
X_5556_ _1128_ _0576_ _2056_ _2057_ _2058_ vssd1 vssd1 vccd1 vccd1 _2059_ sky130_fd_sc_hd__o2111a_1
X_4507_ _1016_ _0326_ _1017_ vssd1 vssd1 vccd1 vccd1 _1018_ sky130_fd_sc_hd__o21ai_1
X_5487_ _3281_ _0780_ vssd1 vssd1 vccd1 vccd1 _1990_ sky130_fd_sc_hd__nand2_1
X_4438_ _0406_ _0948_ vssd1 vssd1 vccd1 vccd1 _0949_ sky130_fd_sc_hd__nand2_1
X_4369_ _0879_ _0422_ _0880_ vssd1 vssd1 vccd1 vccd1 _0881_ sky130_fd_sc_hd__o21ai_1
X_6108_ _2533_ _0829_ vssd1 vssd1 vccd1 vccd1 _2537_ sky130_fd_sc_hd__nand2_1
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6039_ _2494_ _1276_ vssd1 vssd1 vccd1 vccd1 _2497_ sky130_fd_sc_hd__nand2_1
XFILLER_39_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3740_ _3273_ vssd1 vssd1 vccd1 vccd1 _3274_ sky130_fd_sc_hd__inv_2
XFILLER_20_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3671_ _3203_ _3204_ vssd1 vssd1 vccd1 vccd1 _3205_ sky130_fd_sc_hd__nand2_1
X_5410_ _2986_ _3123_ vssd1 vssd1 vccd1 vccd1 _1914_ sky130_fd_sc_hd__nor2_1
XFILLER_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6390_ _2708_ egd_top.BitStream_buffer.BitStream_buffer_output\[13\] vssd1 vssd1
+ vccd1 vccd1 _2760_ sky130_fd_sc_hd__nand2_1
X_5341_ _0467_ _0415_ _0471_ _0419_ _1844_ vssd1 vssd1 vccd1 vccd1 _1845_ sky130_fd_sc_hd__a221oi_1
XFILLER_87_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5272_ _0453_ _0751_ vssd1 vssd1 vccd1 vccd1 _1777_ sky130_fd_sc_hd__nand2_1
X_4223_ _3138_ _3137_ _3173_ _3141_ _0735_ vssd1 vssd1 vccd1 vccd1 _0736_ sky130_fd_sc_hd__a221oi_1
X_4154_ _0471_ _0469_ _0478_ _0473_ _0666_ vssd1 vssd1 vccd1 vccd1 _0667_ sky130_fd_sc_hd__a221oi_2
XFILLER_83_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4085_ _0598_ vssd1 vssd1 vccd1 vccd1 _0599_ sky130_fd_sc_hd__clkbuf_2
XFILLER_63_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4987_ _1479_ _1493_ vssd1 vssd1 vccd1 vccd1 _1494_ sky130_fd_sc_hd__nand2_1
X_6726_ net130 _0185_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[110\]
+ sky130_fd_sc_hd__dfxtp_1
X_3938_ _0451_ vssd1 vssd1 vccd1 vccd1 _0452_ sky130_fd_sc_hd__clkinv_2
X_6657_ clknet_1_1__leaf__2882_ vssd1 vssd1 vccd1 vccd1 _2896_ sky130_fd_sc_hd__buf_1
X_3869_ egd_top.BitStream_buffer.BS_buffer\[43\] vssd1 vssd1 vccd1 vccd1 _0383_ sky130_fd_sc_hd__clkinv_2
X_5608_ _0688_ _0592_ _0611_ _0596_ _2109_ vssd1 vssd1 vccd1 vccd1 _2110_ sky130_fd_sc_hd__o221a_1
X_5539_ egd_top.BitStream_buffer.BS_buffer\[27\] _0487_ egd_top.BitStream_buffer.BS_buffer\[28\]
+ _0490_ _2041_ vssd1 vssd1 vccd1 vccd1 _2042_ sky130_fd_sc_hd__a221oi_1
XFILLER_11_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput17 la_data_in_60_59[0] vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__clkbuf_4
XFILLER_6_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0__f__2894_ clknet_0__2894_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__2894_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_92_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4910_ _3126_ _3075_ vssd1 vssd1 vccd1 vccd1 _1418_ sky130_fd_sc_hd__nand2_1
X_5890_ _0829_ _0439_ _2389_ vssd1 vssd1 vccd1 vccd1 _2390_ sky130_fd_sc_hd__o21ai_1
XFILLER_18_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4841_ _0653_ _0424_ vssd1 vssd1 vccd1 vccd1 _1349_ sky130_fd_sc_hd__or2_1
XFILLER_33_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4772_ _0423_ _0385_ _1280_ vssd1 vssd1 vccd1 vccd1 _1281_ sky130_fd_sc_hd__o21ai_1
X_6511_ _2872_ _2923_ vssd1 vssd1 vccd1 vccd1 _2873_ sky130_fd_sc_hd__nand2_1
X_3723_ _3256_ vssd1 vssd1 vccd1 vccd1 _3257_ sky130_fd_sc_hd__inv_2
X_3654_ _3186_ _3187_ vssd1 vssd1 vccd1 vccd1 _3188_ sky130_fd_sc_hd__nand2_1
X_6442_ _2802_ _2805_ vssd1 vssd1 vccd1 vccd1 _2806_ sky130_fd_sc_hd__nand2_1
X_6373_ _2663_ _2626_ _2681_ vssd1 vssd1 vccd1 vccd1 _2743_ sky130_fd_sc_hd__nand3_1
X_3585_ egd_top.BitStream_buffer.BS_buffer\[105\] vssd1 vssd1 vccd1 vccd1 _3119_ sky130_fd_sc_hd__inv_2
X_5324_ _3026_ _1828_ vssd1 vssd1 vccd1 vccd1 _1829_ sky130_fd_sc_hd__nor2_1
X_5255_ _1754_ _1755_ _1759_ vssd1 vssd1 vccd1 vccd1 _1760_ sky130_fd_sc_hd__nor3_1
XFILLER_87_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4206_ _0718_ _3088_ vssd1 vssd1 vccd1 vccd1 _0719_ sky130_fd_sc_hd__or2_1
X_5186_ _0922_ _0588_ vssd1 vssd1 vccd1 vccd1 _1692_ sky130_fd_sc_hd__or2_1
XFILLER_68_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4137_ egd_top.BitStream_buffer.BS_buffer\[58\] vssd1 vssd1 vccd1 vccd1 _0650_ sky130_fd_sc_hd__clkinv_2
X_4068_ _0581_ vssd1 vssd1 vccd1 vccd1 _0582_ sky130_fd_sc_hd__buf_4
XFILLER_71_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6709_ net113 _0168_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[88\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_22_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6561__104 clknet_1_1__leaf__2887_ vssd1 vssd1 vccd1 vccd1 net138 sky130_fd_sc_hd__inv_2
XFILLER_47_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3370_ _2922_ _2923_ vssd1 vssd1 vccd1 vccd1 _2924_ sky130_fd_sc_hd__nand2_1
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5040_ _3186_ _0562_ vssd1 vssd1 vccd1 vccd1 _1547_ sky130_fd_sc_hd__nand2_1
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5942_ _2438_ _2901_ _2971_ vssd1 vssd1 vccd1 vccd1 _2439_ sky130_fd_sc_hd__and3_1
XFILLER_18_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5873_ _0353_ _0443_ vssd1 vssd1 vccd1 vccd1 _2373_ sky130_fd_sc_hd__nand2_1
X_4824_ _1272_ _1331_ _1332_ vssd1 vssd1 vccd1 vccd1 _1333_ sky130_fd_sc_hd__nand3_1
X_4755_ _3262_ egd_top.BitStream_buffer.BS_buffer\[78\] vssd1 vssd1 vccd1 vccd1 _1264_
+ sky130_fd_sc_hd__nand2_1
X_3706_ _3239_ vssd1 vssd1 vccd1 vccd1 _3240_ sky130_fd_sc_hd__buf_2
X_4686_ _3006_ _3200_ _1195_ vssd1 vssd1 vccd1 vccd1 _1196_ sky130_fd_sc_hd__o21ai_1
X_3637_ _3165_ _3170_ vssd1 vssd1 vccd1 vccd1 _3171_ sky130_fd_sc_hd__nand2_1
X_6425_ net20 net21 vssd1 vssd1 vccd1 vccd1 _2793_ sky130_fd_sc_hd__nand2_1
X_3568_ egd_top.BitStream_buffer.BS_buffer\[101\] vssd1 vssd1 vccd1 vccd1 _3102_ sky130_fd_sc_hd__clkinv_2
X_6356_ _2663_ egd_top.BitStream_buffer.BitStream_buffer_output\[1\] _2681_ vssd1
+ vssd1 vccd1 vccd1 _2727_ sky130_fd_sc_hd__nand3_1
X_5307_ _0688_ _0571_ vssd1 vssd1 vccd1 vccd1 _1812_ sky130_fd_sc_hd__or2_1
XFILLER_68_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3499_ _3030_ _3031_ _3032_ vssd1 vssd1 vccd1 vccd1 _3033_ sky130_fd_sc_hd__and3_4
X_6287_ _2657_ _2624_ vssd1 vssd1 vccd1 vccd1 _2658_ sky130_fd_sc_hd__nand2_1
XFILLER_29_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5238_ _3243_ _3264_ vssd1 vssd1 vccd1 vccd1 _1743_ sky130_fd_sc_hd__nand2_1
X_5169_ _0532_ _0495_ _1674_ vssd1 vssd1 vccd1 vccd1 _1675_ sky130_fd_sc_hd__o21ai_1
XFILLER_56_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4540_ _3259_ egd_top.BitStream_buffer.BS_buffer\[75\] vssd1 vssd1 vccd1 vccd1 _1051_
+ sky130_fd_sc_hd__nand2_1
X_4471_ _0605_ egd_top.BitStream_buffer.BS_buffer\[15\] vssd1 vssd1 vccd1 vccd1 _0982_
+ sky130_fd_sc_hd__nand2_1
X_6210_ _2598_ vssd1 vssd1 vccd1 vccd1 _0178_ sky130_fd_sc_hd__inv_2
X_3422_ _2938_ _2971_ vssd1 vssd1 vccd1 vccd1 _2972_ sky130_fd_sc_hd__or2_1
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6141_ _2966_ _2554_ _2543_ _2556_ vssd1 vssd1 vccd1 vccd1 _0199_ sky130_fd_sc_hd__o211a_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3353_ _2903_ _2900_ _2905_ _2909_ vssd1 vssd1 vccd1 vccd1 _0320_ sky130_fd_sc_hd__a211oi_1
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6072_ _2904_ vssd1 vssd1 vccd1 vccd1 _2516_ sky130_fd_sc_hd__buf_2
XFILLER_85_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5023_ _3127_ _3082_ vssd1 vssd1 vccd1 vccd1 _1530_ sky130_fd_sc_hd__nand2_1
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5925_ _0524_ _0613_ vssd1 vssd1 vccd1 vccd1 _2425_ sky130_fd_sc_hd__or2_1
XFILLER_80_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5856_ _0597_ _3199_ _2355_ vssd1 vssd1 vccd1 vccd1 _2356_ sky130_fd_sc_hd__o21ai_1
X_4807_ _0565_ _0585_ vssd1 vssd1 vccd1 vccd1 _1316_ sky130_fd_sc_hd__nand2_1
X_5787_ _0780_ _3271_ _3322_ _3275_ _2287_ vssd1 vssd1 vccd1 vccd1 _2288_ sky130_fd_sc_hd__a221oi_1
X_4738_ _3018_ _3145_ _1242_ _1246_ vssd1 vssd1 vccd1 vccd1 _1247_ sky130_fd_sc_hd__o211a_1
X_4669_ _3119_ _3105_ vssd1 vssd1 vccd1 vccd1 _1179_ sky130_fd_sc_hd__or2_1
X_6408_ egd_top.BitStream_buffer.BitStream_buffer_output\[4\] _2723_ _2776_ vssd1
+ vssd1 vccd1 vccd1 _2777_ sky130_fd_sc_hd__o21ai_1
X_6339_ _2708_ _2709_ vssd1 vssd1 vccd1 vccd1 _2710_ sky130_fd_sc_hd__and2_1
XFILLER_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6567__110 clknet_1_1__leaf__2887_ vssd1 vssd1 vccd1 vccd1 net144 sky130_fd_sc_hd__inv_2
XFILLER_79_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3971_ _3033_ _0484_ vssd1 vssd1 vccd1 vccd1 _0485_ sky130_fd_sc_hd__and2_1
XFILLER_35_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5710_ _0431_ _3237_ vssd1 vssd1 vccd1 vccd1 _2211_ sky130_fd_sc_hd__nand2_1
X_6690_ clknet_1_0__leaf__2882_ vssd1 vssd1 vccd1 vccd1 _2899_ sky130_fd_sc_hd__buf_1
X_5641_ _3109_ _3340_ _3118_ _0323_ _2142_ vssd1 vssd1 vccd1 vccd1 _2143_ sky130_fd_sc_hd__a221oi_1
X_5572_ _0870_ _0368_ _2073_ vssd1 vssd1 vccd1 vccd1 _2074_ sky130_fd_sc_hd__o21ai_1
X_4523_ _1030_ _1031_ _1032_ _1033_ vssd1 vssd1 vccd1 vccd1 _1034_ sky130_fd_sc_hd__and4_1
X_4454_ egd_top.BitStream_buffer.BS_buffer\[56\] vssd1 vssd1 vccd1 vccd1 _0965_ sky130_fd_sc_hd__inv_2
X_4385_ _0502_ vssd1 vssd1 vccd1 vccd1 _0897_ sky130_fd_sc_hd__clkinv_2
X_3405_ _2957_ _2916_ vssd1 vssd1 vccd1 vccd1 _2958_ sky130_fd_sc_hd__nand2_1
X_6124_ _2538_ _0833_ vssd1 vssd1 vccd1 vccd1 _2546_ sky130_fd_sc_hd__nand2_1
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6055_ _3017_ _2489_ _2501_ _2505_ vssd1 vssd1 vccd1 vccd1 _0234_ sky130_fd_sc_hd__o211a_1
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5006_ _0492_ _0576_ _1510_ _1511_ _1512_ vssd1 vssd1 vccd1 vccd1 _1513_ sky130_fd_sc_hd__o2111a_1
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5908_ _1276_ _0523_ _0861_ _0526_ _2407_ vssd1 vssd1 vccd1 vccd1 _2408_ sky130_fd_sc_hd__o221a_1
XFILLER_14_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5839_ _3332_ _3100_ vssd1 vssd1 vccd1 vccd1 _2339_ sky130_fd_sc_hd__nand2_1
XFILLER_30_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4170_ _0591_ _0595_ vssd1 vssd1 vccd1 vccd1 _0683_ sky130_fd_sc_hd__or2_1
XFILLER_67_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6811_ net55 _0270_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_35_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6742_ net146 _0201_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[78\]
+ sky130_fd_sc_hd__dfxtp_1
X_3954_ _3067_ _2934_ vssd1 vssd1 vccd1 vccd1 _0468_ sky130_fd_sc_hd__nand2_1
X_3885_ _0398_ vssd1 vssd1 vccd1 vccd1 _0399_ sky130_fd_sc_hd__clkbuf_4
XFILLER_50_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5624_ _0389_ _0538_ _0869_ _0541_ _2125_ vssd1 vssd1 vccd1 vccd1 _2126_ sky130_fd_sc_hd__a221oi_1
XFILLER_31_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5555_ _0897_ _0588_ vssd1 vssd1 vccd1 vccd1 _2058_ sky130_fd_sc_hd__or2_1
X_4506_ _0328_ _3341_ vssd1 vssd1 vccd1 vccd1 _1017_ sky130_fd_sc_hd__nand2_1
X_5486_ _1985_ _1986_ _1987_ _1988_ vssd1 vssd1 vccd1 vccd1 _1989_ sky130_fd_sc_hd__and4_1
XFILLER_6_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4437_ egd_top.BitStream_buffer.BS_buffer\[49\] vssd1 vssd1 vccd1 vccd1 _0948_ sky130_fd_sc_hd__clkbuf_4
XFILLER_86_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6107_ _2982_ _2532_ _2528_ _2536_ vssd1 vssd1 vccd1 vccd1 _0213_ sky130_fd_sc_hd__o211a_1
X_4368_ _0659_ _0425_ vssd1 vssd1 vccd1 vccd1 _0880_ sky130_fd_sc_hd__or2_1
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4299_ _3169_ _0726_ _3164_ _3081_ _0810_ vssd1 vssd1 vccd1 vccd1 _0811_ sky130_fd_sc_hd__a221oi_1
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6038_ _2992_ _2487_ _2488_ _2496_ vssd1 vssd1 vccd1 vccd1 _0242_ sky130_fd_sc_hd__o211a_1
XFILLER_46_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3670_ egd_top.BitStream_buffer.BS_buffer\[116\] vssd1 vssd1 vccd1 vccd1 _3204_ sky130_fd_sc_hd__clkbuf_4
XFILLER_40_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5340_ _0448_ _0422_ _1843_ vssd1 vssd1 vccd1 vccd1 _1844_ sky130_fd_sc_hd__o21ai_1
X_5271_ _0458_ _3237_ vssd1 vssd1 vccd1 vccd1 _1776_ sky130_fd_sc_hd__nand2_1
X_4222_ _3006_ _3145_ _0734_ vssd1 vssd1 vccd1 vccd1 _0735_ sky130_fd_sc_hd__o21ai_1
XFILLER_68_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4153_ _0663_ _2935_ _0665_ vssd1 vssd1 vccd1 vccd1 _0666_ sky130_fd_sc_hd__o21ai_1
X_4084_ _3058_ _0556_ vssd1 vssd1 vccd1 vccd1 _0598_ sky130_fd_sc_hd__nand2_1
XFILLER_28_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4986_ _1482_ _1485_ _1489_ _1492_ vssd1 vssd1 vccd1 vccd1 _1493_ sky130_fd_sc_hd__and4_1
X_6725_ net129 _0184_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[111\]
+ sky130_fd_sc_hd__dfxtp_1
X_3937_ _3124_ _2934_ vssd1 vssd1 vccd1 vccd1 _0451_ sky130_fd_sc_hd__nand2_1
X_3868_ _0381_ vssd1 vssd1 vccd1 vccd1 _0382_ sky130_fd_sc_hd__buf_6
X_5607_ _0602_ _0598_ vssd1 vssd1 vccd1 vccd1 _2109_ sky130_fd_sc_hd__or2_1
X_3799_ _3332_ vssd1 vssd1 vccd1 vccd1 _3333_ sky130_fd_sc_hd__buf_2
X_5538_ _0543_ _0495_ _2040_ vssd1 vssd1 vccd1 vccd1 _2041_ sky130_fd_sc_hd__o21ai_1
XFILLER_11_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5469_ _2977_ _3105_ vssd1 vssd1 vccd1 vccd1 _1972_ sky130_fd_sc_hd__or2_1
XTAP_190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput18 la_data_in_60_59[1] vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__buf_2
XFILLER_42_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__2893_ clknet_0__2893_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__2893_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_52_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4840_ _1338_ _1341_ _1344_ _1347_ vssd1 vssd1 vccd1 vccd1 _1348_ sky130_fd_sc_hd__and4_1
XFILLER_33_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6510_ _2866_ _2871_ vssd1 vssd1 vccd1 vccd1 _2872_ sky130_fd_sc_hd__nand2_1
XFILLER_20_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4771_ _0387_ _0642_ vssd1 vssd1 vccd1 vccd1 _1280_ sky130_fd_sc_hd__nand2_1
XFILLER_9_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3722_ egd_top.BitStream_buffer.BS_buffer\[72\] vssd1 vssd1 vccd1 vccd1 _3256_ sky130_fd_sc_hd__clkbuf_4
X_3653_ egd_top.BitStream_buffer.BS_buffer\[127\] vssd1 vssd1 vccd1 vccd1 _3187_ sky130_fd_sc_hd__clkbuf_4
X_6441_ _2804_ vssd1 vssd1 vccd1 vccd1 _2805_ sky130_fd_sc_hd__inv_2
X_6372_ _2680_ _2732_ vssd1 vssd1 vccd1 vccd1 _2742_ sky130_fd_sc_hd__nand2_1
X_5323_ _1769_ _1826_ _1827_ vssd1 vssd1 vccd1 vccd1 _1828_ sky130_fd_sc_hd__nand3_1
X_3584_ egd_top.BitStream_buffer.BS_buffer\[107\] vssd1 vssd1 vccd1 vccd1 _3118_ sky130_fd_sc_hd__clkbuf_4
X_5254_ _0562_ _3179_ _1756_ _1758_ vssd1 vssd1 vccd1 vccd1 _1759_ sky130_fd_sc_hd__a211o_1
X_5185_ _0578_ egd_top.BitStream_buffer.BS_buffer\[16\] vssd1 vssd1 vccd1 vccd1 _1691_
+ sky130_fd_sc_hd__nand2_1
XFILLER_68_330 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4205_ egd_top.BitStream_buffer.BS_buffer\[104\] vssd1 vssd1 vccd1 vccd1 _0718_ sky130_fd_sc_hd__clkinv_2
XFILLER_68_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4136_ _0452_ _0461_ vssd1 vssd1 vccd1 vccd1 _0649_ sky130_fd_sc_hd__nand2_1
XFILLER_83_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4067_ _0559_ _3111_ vssd1 vssd1 vccd1 vccd1 _0581_ sky130_fd_sc_hd__nor2_2
XFILLER_36_271 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4969_ _0406_ _0655_ vssd1 vssd1 vccd1 vccd1 _1476_ sky130_fd_sc_hd__nand2_1
X_6708_ net112 _0167_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[89\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_22_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5941_ _2437_ _2939_ vssd1 vssd1 vccd1 vccd1 _2438_ sky130_fd_sc_hd__nand2_1
X_5872_ _2322_ _2338_ _2354_ _2371_ vssd1 vssd1 vccd1 vccd1 _2372_ sky130_fd_sc_hd__and4_1
XFILLER_21_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4823_ _0622_ _0568_ vssd1 vssd1 vccd1 vccd1 _1332_ sky130_fd_sc_hd__nand2_1
XFILLER_21_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4754_ _3254_ egd_top.BitStream_buffer.BS_buffer\[80\] vssd1 vssd1 vccd1 vccd1 _1263_
+ sky130_fd_sc_hd__nand2_1
X_3705_ _3045_ _3213_ vssd1 vssd1 vccd1 vccd1 _3239_ sky130_fd_sc_hd__nand2_1
X_4685_ _3203_ _0744_ vssd1 vssd1 vccd1 vccd1 _1195_ sky130_fd_sc_hd__nand2_1
X_3636_ _3168_ _3169_ vssd1 vssd1 vccd1 vccd1 _3170_ sky130_fd_sc_hd__nand2_1
X_6424_ _2791_ _2792_ vssd1 vssd1 vccd1 vccd1 net22 sky130_fd_sc_hd__nand2_1
X_3567_ _3099_ _3100_ vssd1 vssd1 vccd1 vccd1 _3101_ sky130_fd_sc_hd__nand2_1
X_6355_ _2680_ _2725_ vssd1 vssd1 vccd1 vccd1 _2726_ sky130_fd_sc_hd__nand2_1
X_6669__42 clknet_1_1__leaf__2897_ vssd1 vssd1 vccd1 vccd1 net76 sky130_fd_sc_hd__inv_2
X_5306_ _0565_ egd_top.BitStream_buffer.BS_buffer\[13\] vssd1 vssd1 vccd1 vccd1 _1811_
+ sky130_fd_sc_hd__nand2_1
X_6286_ _2654_ _2656_ vssd1 vssd1 vccd1 vccd1 _2657_ sky130_fd_sc_hd__nand2_1
XFILLER_88_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3498_ egd_top.BitStream_buffer.pc\[3\] vssd1 vssd1 vccd1 vccd1 _3032_ sky130_fd_sc_hd__clkinv_2
X_6684__56 clknet_1_0__leaf__2898_ vssd1 vssd1 vccd1 vccd1 net90 sky130_fd_sc_hd__inv_2
X_5237_ _3232_ _3252_ vssd1 vssd1 vccd1 vccd1 _1742_ sky130_fd_sc_hd__nand2_1
X_5168_ _0497_ egd_top.BitStream_buffer.BS_buffer\[27\] vssd1 vssd1 vccd1 vccd1 _1674_
+ sky130_fd_sc_hd__nand2_1
XFILLER_84_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5099_ _0930_ _3137_ _1076_ _3141_ _1604_ vssd1 vssd1 vccd1 vccd1 _1605_ sky130_fd_sc_hd__a221oi_1
XFILLER_83_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4119_ _0346_ _0341_ _0344_ _0354_ _0631_ vssd1 vssd1 vccd1 vccd1 _0632_ sky130_fd_sc_hd__a221oi_1
XFILLER_56_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_196 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_355 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4470_ _0608_ egd_top.BitStream_buffer.BS_buffer\[17\] vssd1 vssd1 vccd1 vccd1 _0981_
+ sky130_fd_sc_hd__nand2_1
XFILLER_7_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3421_ _2970_ egd_top.BitStream_buffer.buffer_index\[4\] vssd1 vssd1 vccd1 vccd1
+ _2971_ sky130_fd_sc_hd__nand2_1
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3352_ _2907_ _2908_ vssd1 vssd1 vccd1 vccd1 _2909_ sky130_fd_sc_hd__and2_1
X_6140_ _2555_ _1016_ vssd1 vssd1 vccd1 vccd1 _2556_ sky130_fd_sc_hd__nand2_1
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6071_ _2985_ _2510_ _2501_ _2515_ vssd1 vssd1 vccd1 vccd1 _0228_ sky130_fd_sc_hd__o211a_1
X_5022_ _0808_ _3089_ _1526_ _1527_ _1528_ vssd1 vssd1 vccd1 vccd1 _1529_ sky130_fd_sc_hd__o2111a_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5924_ _0606_ _0531_ vssd1 vssd1 vccd1 vccd1 _2424_ sky130_fd_sc_hd__nand2_1
XFILLER_53_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5855_ _3202_ _0930_ vssd1 vssd1 vccd1 vccd1 _2355_ sky130_fd_sc_hd__nand2_1
XFILLER_21_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4806_ _0561_ egd_top.BitStream_buffer.BS_buffer\[11\] vssd1 vssd1 vccd1 vccd1 _1315_
+ sky130_fd_sc_hd__nand2_1
XFILLER_61_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5786_ _1003_ _3279_ _2286_ vssd1 vssd1 vccd1 vccd1 _2287_ sky130_fd_sc_hd__o21ai_1
X_4737_ _1243_ _1244_ _1245_ vssd1 vssd1 vccd1 vccd1 _1246_ sky130_fd_sc_hd__and3_1
X_6590__131 clknet_1_1__leaf__2889_ vssd1 vssd1 vccd1 vccd1 net165 sky130_fd_sc_hd__inv_2
X_4668_ _3099_ _3109_ vssd1 vssd1 vccd1 vccd1 _1178_ sky130_fd_sc_hd__nand2_1
X_3619_ egd_top.BitStream_buffer.BS_buffer\[114\] vssd1 vssd1 vccd1 vccd1 _3153_ sky130_fd_sc_hd__clkbuf_4
X_6407_ _2723_ _2649_ vssd1 vssd1 vccd1 vccd1 _2776_ sky130_fd_sc_hd__nand2_1
X_4599_ _0829_ _2935_ _1108_ vssd1 vssd1 vccd1 vccd1 _1109_ sky130_fd_sc_hd__o21ai_1
X_6338_ egd_top.BitStream_buffer.BitStream_buffer_output\[12\] egd_top.BitStream_buffer.BitStream_buffer_output\[11\]
+ vssd1 vssd1 vccd1 vccd1 _2709_ sky130_fd_sc_hd__nand2_1
X_6269_ _2639_ vssd1 vssd1 vccd1 vccd1 _2640_ sky130_fd_sc_hd__inv_2
XFILLER_84_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_391 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6648__23 clknet_1_0__leaf__2895_ vssd1 vssd1 vccd1 vccd1 net57 sky130_fd_sc_hd__inv_2
XFILLER_69_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6663__37 clknet_1_1__leaf__2896_ vssd1 vssd1 vccd1 vccd1 net71 sky130_fd_sc_hd__inv_2
XFILLER_39_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3970_ _2932_ _3034_ egd_top.BitStream_buffer.pc\[4\] vssd1 vssd1 vccd1 vccd1 _0484_
+ sky130_fd_sc_hd__and3_2
XFILLER_62_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5640_ _3119_ _0327_ _2141_ vssd1 vssd1 vccd1 vccd1 _2142_ sky130_fd_sc_hd__o21ai_1
X_5571_ _0371_ _0393_ vssd1 vssd1 vccd1 vccd1 _2073_ sky130_fd_sc_hd__nand2_1
X_4522_ _3038_ _3062_ vssd1 vssd1 vccd1 vccd1 _1033_ sky130_fd_sc_hd__nand2_1
XFILLER_7_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4453_ _0960_ _0421_ _0961_ _0962_ _0963_ vssd1 vssd1 vccd1 vccd1 _0964_ sky130_fd_sc_hd__o2111a_1
X_3404_ net29 net28 vssd1 vssd1 vccd1 vccd1 _2957_ sky130_fd_sc_hd__nand2_1
X_4384_ _0878_ _0895_ vssd1 vssd1 vccd1 vccd1 _0896_ sky130_fd_sc_hd__nand2_1
XFILLER_58_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6123_ _3005_ _2532_ _2543_ _2545_ vssd1 vssd1 vccd1 vccd1 _0206_ sky130_fd_sc_hd__o211a_1
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6054_ _2494_ _0870_ vssd1 vssd1 vccd1 vccd1 _2505_ sky130_fd_sc_hd__nand2_1
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5005_ _0685_ _0588_ vssd1 vssd1 vccd1 vccd1 _1512_ sky130_fd_sc_hd__or2_1
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_420 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5907_ _0348_ _0530_ _0629_ _0534_ vssd1 vssd1 vccd1 vccd1 _2407_ sky130_fd_sc_hd__o22a_1
XFILLER_34_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5838_ _2326_ _2330_ _2334_ _2337_ vssd1 vssd1 vccd1 vccd1 _2338_ sky130_fd_sc_hd__and4_1
X_5769_ _3203_ _0792_ vssd1 vssd1 vccd1 vccd1 _2270_ sky130_fd_sc_hd__nand2_1
XFILLER_89_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6597__137 clknet_1_1__leaf__2890_ vssd1 vssd1 vccd1 vccd1 net171 sky130_fd_sc_hd__inv_2
XFILLER_71_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6810_ net54 _0269_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_23_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3953_ egd_top.BitStream_buffer.BS_buffer\[60\] vssd1 vssd1 vccd1 vccd1 _0467_ sky130_fd_sc_hd__clkbuf_4
X_6741_ net145 _0200_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[79\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_50_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3884_ _0397_ vssd1 vssd1 vccd1 vccd1 _0398_ sky130_fd_sc_hd__clkbuf_2
X_5623_ _0861_ _0545_ _2124_ vssd1 vssd1 vccd1 vccd1 _2125_ sky130_fd_sc_hd__o21ai_1
XFILLER_31_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5554_ _0582_ _0505_ vssd1 vssd1 vccd1 vccd1 _2057_ sky130_fd_sc_hd__nand2_1
X_4505_ egd_top.BitStream_buffer.BS_buffer\[96\] vssd1 vssd1 vccd1 vccd1 _1016_ sky130_fd_sc_hd__inv_2
X_5485_ _3250_ egd_top.BitStream_buffer.BS_buffer\[85\] vssd1 vssd1 vccd1 vccd1 _1988_
+ sky130_fd_sc_hd__nand2_1
X_4436_ _0400_ _0388_ _0407_ _0944_ _0946_ vssd1 vssd1 vccd1 vccd1 _0947_ sky130_fd_sc_hd__a221oi_1
X_4367_ egd_top.BitStream_buffer.BS_buffer\[51\] vssd1 vssd1 vccd1 vccd1 _0879_ sky130_fd_sc_hd__inv_2
XFILLER_76_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6106_ _2533_ _1297_ vssd1 vssd1 vccd1 vccd1 _2536_ sky130_fd_sc_hd__nand2_1
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4298_ _0808_ _0729_ _0809_ vssd1 vssd1 vccd1 vccd1 _0810_ sky130_fd_sc_hd__o21ai_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6642__18 clknet_1_0__leaf__2894_ vssd1 vssd1 vccd1 vccd1 net52 sky130_fd_sc_hd__inv_2
X_6037_ _2494_ _1084_ vssd1 vssd1 vccd1 vccd1 _2496_ sky130_fd_sc_hd__nand2_1
XFILLER_92_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6605__144 clknet_1_0__leaf__2891_ vssd1 vssd1 vccd1 vccd1 net178 sky130_fd_sc_hd__inv_2
XFILLER_32_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5270_ _0664_ _0432_ _0435_ _3244_ _1774_ vssd1 vssd1 vccd1 vccd1 _1775_ sky130_fd_sc_hd__a221oi_1
X_4221_ _3148_ _3133_ vssd1 vssd1 vccd1 vccd1 _0734_ sky130_fd_sc_hd__nand2_1
XFILLER_49_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4152_ _0476_ _0664_ vssd1 vssd1 vccd1 vccd1 _0665_ sky130_fd_sc_hd__nand2_1
X_4083_ egd_top.BitStream_buffer.BS_buffer\[3\] vssd1 vssd1 vccd1 vccd1 _0597_ sky130_fd_sc_hd__inv_2
XFILLER_83_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4985_ _3217_ _0477_ _3221_ _2936_ _1491_ vssd1 vssd1 vccd1 vccd1 _1492_ sky130_fd_sc_hd__a221oi_1
X_3936_ _0449_ vssd1 vssd1 vccd1 vccd1 _0450_ sky130_fd_sc_hd__clkbuf_4
XFILLER_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6724_ net128 _0183_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.pc_previous\[6\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_31_191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3867_ _0380_ vssd1 vssd1 vccd1 vccd1 _0381_ sky130_fd_sc_hd__inv_2
X_5606_ _0986_ _0588_ _2105_ _2106_ _2107_ vssd1 vssd1 vccd1 vccd1 _2108_ sky130_fd_sc_hd__o2111a_1
X_3798_ _3331_ vssd1 vssd1 vccd1 vccd1 _3332_ sky130_fd_sc_hd__clkinv_2
X_5537_ _0497_ _0537_ vssd1 vssd1 vccd1 vccd1 _2040_ sky130_fd_sc_hd__nand2_1
XFILLER_3_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5468_ _3098_ egd_top.BitStream_buffer.BS_buffer\[113\] vssd1 vssd1 vccd1 vccd1 _1971_
+ sky130_fd_sc_hd__nand2_1
X_4419_ _0622_ _0930_ vssd1 vssd1 vccd1 vccd1 _0931_ sky130_fd_sc_hd__nand2_1
X_5399_ _3243_ _3248_ vssd1 vssd1 vccd1 vccd1 _1903_ sky130_fd_sc_hd__nand2_1
XTAP_191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput19 la_data_in_65 vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_22_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0__f__2892_ clknet_0__2892_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__2892_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_18_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4770_ _0347_ _0360_ _0363_ _0375_ _1278_ vssd1 vssd1 vccd1 vccd1 _1279_ sky130_fd_sc_hd__a221oi_1
XFILLER_33_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3721_ _3254_ vssd1 vssd1 vccd1 vccd1 _3255_ sky130_fd_sc_hd__buf_4
X_3652_ _3185_ vssd1 vssd1 vccd1 vccd1 _3186_ sky130_fd_sc_hd__buf_2
X_6440_ egd_top.BitStream_buffer.BitStream_buffer_output\[5\] _2678_ _2803_ vssd1
+ vssd1 vccd1 vccd1 _2804_ sky130_fd_sc_hd__o21ai_2
X_3583_ _3116_ vssd1 vssd1 vccd1 vccd1 _3117_ sky130_fd_sc_hd__buf_2
XFILLER_9_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6371_ _2923_ _2685_ _2695_ _2700_ _2741_ vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__o221ai_4
X_5322_ _0621_ _0585_ vssd1 vssd1 vccd1 vccd1 _1827_ sky130_fd_sc_hd__nand2_1
XFILLER_5_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5253_ _0554_ _3182_ _1757_ vssd1 vssd1 vccd1 vccd1 _1758_ sky130_fd_sc_hd__o21ai_1
X_6550__94 clknet_1_0__leaf__2886_ vssd1 vssd1 vccd1 vccd1 net128 sky130_fd_sc_hd__inv_2
X_5184_ _0582_ _0491_ vssd1 vssd1 vccd1 vccd1 _1690_ sky130_fd_sc_hd__nand2_1
X_4204_ _3093_ _0716_ vssd1 vssd1 vccd1 vccd1 _0717_ sky130_fd_sc_hd__nand2_1
XFILLER_68_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4135_ _0457_ _0447_ vssd1 vssd1 vccd1 vccd1 _0648_ sky130_fd_sc_hd__nand2_1
X_4066_ _0578_ _0579_ vssd1 vssd1 vccd1 vccd1 _0580_ sky130_fd_sc_hd__nand2_1
XFILLER_83_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4968_ _0642_ _0378_ _0874_ _0382_ _1474_ vssd1 vssd1 vccd1 vccd1 _1475_ sky130_fd_sc_hd__a221oi_1
X_4899_ _0709_ _0326_ _1406_ vssd1 vssd1 vccd1 vccd1 _1407_ sky130_fd_sc_hd__o21ai_1
XFILLER_11_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6707_ net111 _0166_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[90\]
+ sky130_fd_sc_hd__dfxtp_1
X_3919_ _3087_ _2933_ vssd1 vssd1 vccd1 vccd1 _0433_ sky130_fd_sc_hd__and2_1
X_6569_ clknet_1_0__leaf__2883_ vssd1 vssd1 vccd1 vccd1 _2888_ sky130_fd_sc_hd__buf_1
XFILLER_78_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_507 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5940_ _2970_ vssd1 vssd1 vccd1 vccd1 _2437_ sky130_fd_sc_hd__inv_2
XFILLER_92_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_326 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5871_ _2357_ _2362_ _2367_ _2370_ vssd1 vssd1 vccd1 vccd1 _2371_ sky130_fd_sc_hd__and4_1
X_4822_ _1302_ _1330_ vssd1 vssd1 vccd1 vccd1 _1331_ sky130_fd_sc_hd__nor2_1
X_4753_ _0755_ _3239_ _1259_ _1260_ _1261_ vssd1 vssd1 vccd1 vccd1 _1262_ sky130_fd_sc_hd__o2111a_1
X_3704_ egd_top.BitStream_buffer.BS_buffer\[65\] vssd1 vssd1 vccd1 vccd1 _3238_ sky130_fd_sc_hd__clkinv_2
X_4684_ _3191_ _3156_ _3198_ _3160_ _1193_ vssd1 vssd1 vccd1 vccd1 _1194_ sky130_fd_sc_hd__a221oi_1
X_6423_ _2923_ _2699_ _2766_ vssd1 vssd1 vccd1 vccd1 _2792_ sky130_fd_sc_hd__or3_1
X_3635_ egd_top.BitStream_buffer.BS_buffer\[112\] vssd1 vssd1 vccd1 vccd1 _3169_ sky130_fd_sc_hd__clkbuf_4
X_3566_ egd_top.BitStream_buffer.BS_buffer\[102\] vssd1 vssd1 vccd1 vccd1 _3100_ sky130_fd_sc_hd__clkbuf_4
X_6354_ _2627_ _2723_ _2724_ vssd1 vssd1 vccd1 vccd1 _2725_ sky130_fd_sc_hd__o21ai_1
X_5305_ _0561_ egd_top.BitStream_buffer.BS_buffer\[15\] vssd1 vssd1 vccd1 vccd1 _1810_
+ sky130_fd_sc_hd__nand2_1
X_3497_ egd_top.BitStream_buffer.pc\[2\] vssd1 vssd1 vccd1 vccd1 _3031_ sky130_fd_sc_hd__clkinv_2
X_6285_ _2655_ egd_top.BitStream_buffer.BitStream_buffer_output\[11\] egd_top.BitStream_buffer.BitStream_buffer_output\[13\]
+ vssd1 vssd1 vccd1 vccd1 _2656_ sky130_fd_sc_hd__a21oi_1
XFILLER_88_448 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5236_ _0767_ _3260_ _1738_ _1739_ _1740_ vssd1 vssd1 vccd1 vccd1 _1741_ sky130_fd_sc_hd__o2111a_1
X_5167_ _1658_ _1672_ vssd1 vssd1 vccd1 vccd1 _1673_ sky130_fd_sc_hd__nand2_1
X_5098_ _1602_ _3145_ _1603_ vssd1 vssd1 vccd1 vccd1 _1604_ sky130_fd_sc_hd__o21ai_1
X_4118_ _0629_ _0349_ _0630_ vssd1 vssd1 vccd1 vccd1 _0631_ sky130_fd_sc_hd__o21ai_1
X_4049_ _0561_ _0562_ vssd1 vssd1 vccd1 vccd1 _0563_ sky130_fd_sc_hd__nand2_1
XFILLER_17_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_507 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_367 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3420_ _2969_ _2961_ vssd1 vssd1 vccd1 vccd1 _2970_ sky130_fd_sc_hd__nand2_2
X_3351_ net33 vssd1 vssd1 vccd1 vccd1 _2908_ sky130_fd_sc_hd__inv_2
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6070_ _2511_ _0879_ vssd1 vssd1 vccd1 vccd1 _2515_ sky130_fd_sc_hd__nand2_1
X_5021_ _1025_ _3106_ vssd1 vssd1 vccd1 vccd1 _1528_ sky130_fd_sc_hd__or2_1
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5923_ _0609_ egd_top.BitStream_buffer.BS_buffer\[28\] vssd1 vssd1 vccd1 vccd1 _2423_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5854_ _2341_ _2345_ _2350_ _2353_ vssd1 vssd1 vccd1 vccd1 _2354_ sky130_fd_sc_hd__and4_1
X_4805_ _1305_ _1308_ _1310_ _1313_ vssd1 vssd1 vccd1 vccd1 _1314_ sky130_fd_sc_hd__and4_1
XFILLER_21_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5785_ _3282_ _3327_ vssd1 vssd1 vccd1 vccd1 _2286_ sky130_fd_sc_hd__nand2_1
X_4736_ _3136_ egd_top.BitStream_buffer.BS_buffer\[127\] vssd1 vssd1 vccd1 vccd1 _1245_
+ sky130_fd_sc_hd__nand2_1
X_4667_ _3093_ _3128_ vssd1 vssd1 vccd1 vccd1 _1177_ sky130_fd_sc_hd__nand2_1
X_3618_ _3133_ _3137_ _3138_ _3141_ _3151_ vssd1 vssd1 vccd1 vccd1 _3152_ sky130_fd_sc_hd__a221oi_1
X_6406_ _2680_ _2732_ _2745_ vssd1 vssd1 vccd1 vccd1 _2775_ sky130_fd_sc_hd__nand3_1
X_4598_ _0476_ egd_top.BitStream_buffer.BS_buffer\[66\] vssd1 vssd1 vccd1 vccd1 _1108_
+ sky130_fd_sc_hd__nand2_1
X_6337_ _2655_ _2631_ vssd1 vssd1 vccd1 vccd1 _2708_ sky130_fd_sc_hd__nand2_1
X_3549_ _3075_ _3078_ _3081_ _3082_ vssd1 vssd1 vccd1 vccd1 _3083_ sky130_fd_sc_hd__a22o_1
XFILLER_88_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6268_ _2623_ _2624_ vssd1 vssd1 vccd1 vccd1 _2639_ sky130_fd_sc_hd__nand2_1
XFILLER_88_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6199_ _2593_ vssd1 vssd1 vccd1 vccd1 _0181_ sky130_fd_sc_hd__inv_2
X_5219_ _3295_ _0330_ vssd1 vssd1 vccd1 vccd1 _1724_ sky130_fd_sc_hd__nand2_1
XFILLER_29_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6574__116 clknet_1_1__leaf__2888_ vssd1 vssd1 vccd1 vccd1 net150 sky130_fd_sc_hd__inv_2
XFILLER_79_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5570_ egd_top.BitStream_buffer.BitStream_buffer_output\[3\] _2965_ _0627_ vssd1
+ vssd1 vccd1 vccd1 _2072_ sky130_fd_sc_hd__o21ai_1
X_4521_ _3054_ egd_top.BitStream_buffer.BS_buffer\[101\] vssd1 vssd1 vccd1 vccd1 _1032_
+ sky130_fd_sc_hd__nand2_1
X_4452_ _0418_ _0429_ vssd1 vssd1 vccd1 vccd1 _0963_ sky130_fd_sc_hd__nand2_1
X_3403_ _2956_ vssd1 vssd1 vccd1 vccd1 _0317_ sky130_fd_sc_hd__inv_2
X_4383_ _0882_ _0886_ _0891_ _0894_ vssd1 vssd1 vccd1 vccd1 _0895_ sky130_fd_sc_hd__and4_1
X_6122_ _2538_ _0759_ vssd1 vssd1 vccd1 vccd1 _2545_ sky130_fd_sc_hd__nand2_1
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6053_ _3014_ _2489_ _2501_ _2504_ vssd1 vssd1 vccd1 vccd1 _0235_ sky130_fd_sc_hd__o211a_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5004_ _0578_ egd_top.BitStream_buffer.BS_buffer\[15\] vssd1 vssd1 vccd1 vccd1 _1511_
+ sky130_fd_sc_hd__nand2_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5906_ egd_top.BitStream_buffer.BS_buffer\[34\] _0504_ _0364_ _0508_ _2405_ vssd1
+ vssd1 vccd1 vccd1 _2406_ sky130_fd_sc_hd__a221oi_1
XFILLER_53_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5837_ _3173_ _3078_ _3177_ _3080_ _2336_ vssd1 vssd1 vccd1 vccd1 _2337_ sky130_fd_sc_hd__a221oi_1
X_5768_ _3187_ _3156_ _0623_ _3160_ _2268_ vssd1 vssd1 vccd1 vccd1 _2269_ sky130_fd_sc_hd__a221oi_1
X_4719_ _3092_ _0722_ vssd1 vssd1 vccd1 vccd1 _1228_ sky130_fd_sc_hd__nand2_1
XFILLER_5_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5699_ _0405_ _0447_ vssd1 vssd1 vccd1 vccd1 _2200_ sky130_fd_sc_hd__nand2_1
XFILLER_1_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_384 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6740_ net144 _0199_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[96\]
+ sky130_fd_sc_hd__dfxtp_2
X_3952_ _0448_ _0450_ _0455_ _0460_ _0465_ vssd1 vssd1 vccd1 vccd1 _0466_ sky130_fd_sc_hd__o2111a_1
X_3883_ _3071_ _0338_ vssd1 vssd1 vccd1 vccd1 _0397_ sky130_fd_sc_hd__and2_1
XFILLER_50_159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5622_ _0547_ _0375_ vssd1 vssd1 vccd1 vccd1 _2124_ sky130_fd_sc_hd__nand2_1
X_5553_ _0578_ _0498_ vssd1 vssd1 vccd1 vccd1 _2056_ sky130_fd_sc_hd__nand2_1
X_4504_ _0779_ _3307_ _1012_ _1013_ _1014_ vssd1 vssd1 vccd1 vccd1 _1015_ sky130_fd_sc_hd__o2111a_1
X_5484_ _3259_ egd_top.BitStream_buffer.BS_buffer\[83\] vssd1 vssd1 vccd1 vccd1 _1987_
+ sky130_fd_sc_hd__nand2_1
X_4435_ _0637_ _0380_ _0945_ vssd1 vssd1 vccd1 vccd1 _0946_ sky130_fd_sc_hd__o21ai_1
XFILLER_6_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4366_ _0864_ _0868_ _0873_ _0877_ vssd1 vssd1 vccd1 vccd1 _0878_ sky130_fd_sc_hd__and4_1
XFILLER_86_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6105_ _2979_ _2532_ _2528_ _2535_ vssd1 vssd1 vccd1 vccd1 _0214_ sky130_fd_sc_hd__o211a_1
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4297_ _3074_ _3082_ vssd1 vssd1 vccd1 vccd1 _0809_ sky130_fd_sc_hd__nand2_1
XFILLER_58_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6036_ _2988_ _2487_ _2488_ _2495_ vssd1 vssd1 vccd1 vccd1 _0243_ sky130_fd_sc_hd__o211a_1
XFILLER_54_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4220_ _0712_ _0720_ _0725_ _0732_ vssd1 vssd1 vccd1 vccd1 _0733_ sky130_fd_sc_hd__and4_1
XFILLER_68_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4151_ egd_top.BitStream_buffer.BS_buffer\[63\] vssd1 vssd1 vccd1 vccd1 _0664_ sky130_fd_sc_hd__clkbuf_4
XFILLER_83_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4082_ _0595_ vssd1 vssd1 vccd1 vccd1 _0596_ sky130_fd_sc_hd__buf_2
XFILLER_83_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4984_ _1043_ _0472_ _1490_ vssd1 vssd1 vccd1 vccd1 _1491_ sky130_fd_sc_hd__o21ai_1
XFILLER_36_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6723_ net127 _0182_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.pc_previous\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_3935_ _3114_ _2934_ vssd1 vssd1 vccd1 vccd1 _0449_ sky130_fd_sc_hd__nand2_2
XFILLER_51_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_468 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5605_ _0510_ _0575_ vssd1 vssd1 vccd1 vccd1 _2107_ sky130_fd_sc_hd__or2_1
X_3866_ _3121_ _0338_ vssd1 vssd1 vccd1 vccd1 _0380_ sky130_fd_sc_hd__nand2_2
X_3797_ _3124_ _3297_ vssd1 vssd1 vccd1 vccd1 _3331_ sky130_fd_sc_hd__nand2_1
XFILLER_11_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5536_ _2024_ _2038_ vssd1 vssd1 vccd1 vccd1 _2039_ sky130_fd_sc_hd__nand2_1
X_5467_ _3092_ _3082_ vssd1 vssd1 vccd1 vccd1 _1970_ sky130_fd_sc_hd__nand2_1
X_4418_ egd_top.BitStream_buffer.BS_buffer\[2\] vssd1 vssd1 vccd1 vccd1 _0930_ sky130_fd_sc_hd__clkbuf_4
X_5398_ _3315_ _3251_ _0774_ _3255_ _1901_ vssd1 vssd1 vccd1 vccd1 _1902_ sky130_fd_sc_hd__a221oi_1
XFILLER_86_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4349_ egd_top.BitStream_buffer.BS_buffer\[41\] vssd1 vssd1 vccd1 vccd1 _0861_ sky130_fd_sc_hd__clkinv_2
XFILLER_86_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6019_ _2464_ _0907_ vssd1 vssd1 vccd1 vccd1 _2484_ sky130_fd_sc_hd__nand2_1
XFILLER_36_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__2891_ clknet_0__2891_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__2891_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_37_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3720_ _3253_ vssd1 vssd1 vccd1 vccd1 _3254_ sky130_fd_sc_hd__buf_4
X_3651_ _3184_ vssd1 vssd1 vccd1 vccd1 _3185_ sky130_fd_sc_hd__clkbuf_2
X_3582_ _3041_ _3115_ vssd1 vssd1 vccd1 vccd1 _3116_ sky130_fd_sc_hd__nor2_2
XFILLER_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6370_ _2701_ _2735_ _2737_ _2740_ vssd1 vssd1 vccd1 vccd1 _2741_ sky130_fd_sc_hd__a211o_1
X_5321_ _1797_ _1825_ vssd1 vssd1 vccd1 vccd1 _1826_ sky130_fd_sc_hd__nor2_1
X_6535__81 clknet_1_1__leaf__2884_ vssd1 vssd1 vccd1 vccd1 net115 sky130_fd_sc_hd__inv_2
XFILLER_87_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5252_ _3185_ _0579_ vssd1 vssd1 vccd1 vccd1 _1757_ sky130_fd_sc_hd__nand2_1
X_5183_ _0602_ _0558_ _1686_ _1687_ _1688_ vssd1 vssd1 vccd1 vccd1 _1689_ sky130_fd_sc_hd__o2111a_1
X_4203_ egd_top.BitStream_buffer.BS_buffer\[101\] vssd1 vssd1 vccd1 vccd1 _0716_ sky130_fd_sc_hd__clkbuf_4
XFILLER_68_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4134_ _0467_ vssd1 vssd1 vccd1 vccd1 _0647_ sky130_fd_sc_hd__clkinv_2
X_6627__4 clknet_1_1__leaf__2893_ vssd1 vssd1 vccd1 vccd1 net38 sky130_fd_sc_hd__inv_2
XFILLER_83_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4065_ egd_top.BitStream_buffer.BS_buffer\[8\] vssd1 vssd1 vccd1 vccd1 _0579_ sky130_fd_sc_hd__clkbuf_4
XFILLER_51_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4967_ _0659_ _0385_ _1473_ vssd1 vssd1 vccd1 vccd1 _1474_ sky130_fd_sc_hd__o21ai_1
X_4898_ _0328_ _0708_ vssd1 vssd1 vccd1 vccd1 _1406_ sky130_fd_sc_hd__nand2_1
X_3918_ _0431_ vssd1 vssd1 vccd1 vccd1 _0432_ sky130_fd_sc_hd__buf_2
X_6706_ net110 _0165_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[91\]
+ sky130_fd_sc_hd__dfxtp_1
X_3849_ _0362_ vssd1 vssd1 vccd1 vccd1 _0363_ sky130_fd_sc_hd__clkbuf_4
XFILLER_3_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5519_ _0650_ _0403_ _2021_ vssd1 vssd1 vccd1 vccd1 _2022_ sky130_fd_sc_hd__o21ai_1
X_6499_ _2695_ _2860_ vssd1 vssd1 vccd1 vccd1 _2861_ sky130_fd_sc_hd__nor2_1
XFILLER_47_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_51 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5870_ _0583_ _3176_ egd_top.BitStream_buffer.BS_buffer\[11\] _3179_ _2369_ vssd1
+ vssd1 vccd1 vccd1 _2370_ sky130_fd_sc_hd__a221oi_1
XFILLER_61_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4821_ _1314_ _1329_ vssd1 vssd1 vccd1 vccd1 _1330_ sky130_fd_sc_hd__nand2_1
XFILLER_21_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4752_ _3235_ _3256_ vssd1 vssd1 vccd1 vccd1 _1261_ sky130_fd_sc_hd__nand2_1
X_4683_ _1191_ _1192_ vssd1 vssd1 vccd1 vccd1 _1193_ sky130_fd_sc_hd__nand2_1
X_3703_ egd_top.BitStream_buffer.BS_buffer\[67\] vssd1 vssd1 vccd1 vccd1 _3237_ sky130_fd_sc_hd__clkbuf_4
X_3634_ _3167_ vssd1 vssd1 vccd1 vccd1 _3168_ sky130_fd_sc_hd__buf_2
X_6422_ _2787_ _2736_ _2790_ vssd1 vssd1 vccd1 vccd1 _2791_ sky130_fd_sc_hd__nand3_1
X_3565_ _3098_ vssd1 vssd1 vccd1 vccd1 _3099_ sky130_fd_sc_hd__buf_4
X_6353_ _2723_ egd_top.BitStream_buffer.BitStream_buffer_output\[4\] vssd1 vssd1 vccd1
+ vccd1 _2724_ sky130_fd_sc_hd__nand2_1
X_5304_ _1800_ _1803_ _1805_ _1808_ vssd1 vssd1 vccd1 vccd1 _1809_ sky130_fd_sc_hd__and4_1
X_3496_ _3029_ vssd1 vssd1 vccd1 vccd1 _3030_ sky130_fd_sc_hd__inv_2
XFILLER_0_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6284_ egd_top.BitStream_buffer.BitStream_buffer_output\[12\] vssd1 vssd1 vccd1 vccd1
+ _2655_ sky130_fd_sc_hd__inv_2
X_5235_ _3263_ _3288_ vssd1 vssd1 vccd1 vccd1 _1740_ sky130_fd_sc_hd__nand2_1
X_5166_ _1661_ _1664_ _1668_ _1671_ vssd1 vssd1 vccd1 vccd1 _1672_ sky130_fd_sc_hd__and4_1
XFILLER_29_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5097_ _3148_ _0792_ vssd1 vssd1 vccd1 vccd1 _1603_ sky130_fd_sc_hd__nand2_1
XFILLER_68_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4117_ _0352_ _0347_ vssd1 vssd1 vccd1 vccd1 _0630_ sky130_fd_sc_hd__nand2_1
XFILLER_17_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4048_ egd_top.BitStream_buffer.BS_buffer\[6\] vssd1 vssd1 vccd1 vccd1 _0562_ sky130_fd_sc_hd__clkbuf_4
XFILLER_71_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5999_ _2992_ _2465_ _2458_ _2473_ vssd1 vssd1 vccd1 vccd1 _0258_ sky130_fd_sc_hd__o211a_1
XFILLER_33_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_416 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3350_ net34 _2906_ net32 vssd1 vssd1 vccd1 vccd1 _2907_ sky130_fd_sc_hd__or3b_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5020_ _3099_ _3070_ vssd1 vssd1 vccd1 vccd1 _1527_ sky130_fd_sc_hd__nand2_1
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5922_ _0685_ _0593_ _0922_ _0599_ _2421_ vssd1 vssd1 vccd1 vccd1 _2422_ sky130_fd_sc_hd__o221a_1
X_5853_ _3066_ _3339_ _3070_ _0322_ _2352_ vssd1 vssd1 vccd1 vccd1 _2353_ sky130_fd_sc_hd__a221oi_1
X_4804_ _0364_ _0539_ _0337_ _0542_ _1312_ vssd1 vssd1 vccd1 vccd1 _1313_ sky130_fd_sc_hd__a221oi_1
XFILLER_61_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5784_ _0772_ _3251_ _3334_ _3255_ _2284_ vssd1 vssd1 vccd1 vccd1 _2285_ sky130_fd_sc_hd__a221oi_1
X_4735_ _3147_ egd_top.BitStream_buffer.BS_buffer\[126\] vssd1 vssd1 vccd1 vccd1 _1244_
+ sky130_fd_sc_hd__nand2_1
XFILLER_21_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4666_ _3094_ _3039_ _0716_ _3048_ _1175_ vssd1 vssd1 vccd1 vccd1 _1176_ sky130_fd_sc_hd__a221oi_2
X_3617_ _3003_ _3145_ _3150_ vssd1 vssd1 vccd1 vccd1 _3151_ sky130_fd_sc_hd__o21ai_1
X_6405_ _2771_ _2745_ _2773_ vssd1 vssd1 vccd1 vccd1 _2774_ sky130_fd_sc_hd__nand3_1
X_4597_ _1105_ _1106_ vssd1 vssd1 vccd1 vccd1 _1107_ sky130_fd_sc_hd__nor2_1
X_3548_ egd_top.BitStream_buffer.BS_buffer\[111\] vssd1 vssd1 vccd1 vccd1 _3082_ sky130_fd_sc_hd__clkbuf_4
X_6336_ _2705_ _2706_ vssd1 vssd1 vccd1 vccd1 _2707_ sky130_fd_sc_hd__nand2_1
XFILLER_0_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6267_ _2633_ _2622_ vssd1 vssd1 vccd1 vccd1 _2638_ sky130_fd_sc_hd__nand2_1
X_3479_ _3014_ _2976_ _3002_ _3016_ vssd1 vssd1 vccd1 vccd1 _0301_ sky130_fd_sc_hd__o211a_1
XFILLER_88_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6198_ _2902_ egd_top.BitStream_buffer.pc\[4\] vssd1 vssd1 vccd1 vccd1 _2593_ sky130_fd_sc_hd__nand2_1
X_5218_ _3300_ _3322_ vssd1 vssd1 vccd1 vccd1 _1723_ sky130_fd_sc_hd__nand2_1
XFILLER_69_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5149_ _0406_ _0429_ vssd1 vssd1 vccd1 vccd1 _1655_ sky130_fd_sc_hd__nand2_1
XFILLER_44_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_55 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4520_ _3047_ egd_top.BitStream_buffer.BS_buffer\[100\] vssd1 vssd1 vccd1 vccd1 _1031_
+ sky130_fd_sc_hd__nand2_1
X_4451_ _0414_ _0655_ vssd1 vssd1 vccd1 vccd1 _0962_ sky130_fd_sc_hd__nand2_1
X_3402_ net30 _2951_ _2902_ _2955_ vssd1 vssd1 vccd1 vccd1 _2956_ sky130_fd_sc_hd__o211ai_1
X_4382_ _0478_ _0470_ _0664_ _0473_ _0893_ vssd1 vssd1 vccd1 vccd1 _0894_ sky130_fd_sc_hd__a221oi_1
X_6121_ _3001_ _2532_ _2543_ _2544_ vssd1 vssd1 vccd1 vccd1 _0207_ sky130_fd_sc_hd__o211a_1
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6052_ _2494_ _0637_ vssd1 vssd1 vccd1 vccd1 _2504_ sky130_fd_sc_hd__nand2_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5003_ _0582_ egd_top.BitStream_buffer.BS_buffer\[17\] vssd1 vssd1 vccd1 vccd1 _1510_
+ sky130_fd_sc_hd__nand2_1
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5905_ _1084_ _0512_ _2404_ vssd1 vssd1 vccd1 vccd1 _2405_ sky130_fd_sc_hd__o21ai_1
XFILLER_14_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5836_ _3009_ _0728_ _2335_ vssd1 vssd1 vccd1 vccd1 _2336_ sky130_fd_sc_hd__o21ai_1
X_5767_ _2266_ _2267_ vssd1 vssd1 vccd1 vccd1 _2268_ sky130_fd_sc_hd__nand2_1
X_4718_ _3098_ _3118_ vssd1 vssd1 vccd1 vccd1 _1227_ sky130_fd_sc_hd__nand2_1
X_5698_ _0655_ _0378_ _0429_ _0382_ _2198_ vssd1 vssd1 vccd1 vccd1 _2199_ sky130_fd_sc_hd__a221oi_1
X_4649_ _3301_ _0774_ vssd1 vssd1 vccd1 vccd1 _1159_ sky130_fd_sc_hd__nand2_1
X_6319_ _2689_ _2625_ vssd1 vssd1 vccd1 vccd1 _2690_ sky130_fd_sc_hd__nor2b_1
XFILLER_1_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_89 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3951_ _0462_ _0464_ vssd1 vssd1 vccd1 vccd1 _0465_ sky130_fd_sc_hd__or2_1
XFILLER_35_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3882_ _0395_ vssd1 vssd1 vccd1 vccd1 _0396_ sky130_fd_sc_hd__clkbuf_4
X_5621_ _0865_ _0511_ _2120_ _2121_ _2122_ vssd1 vssd1 vccd1 vccd1 _2123_ sky130_fd_sc_hd__o2111a_1
X_5552_ _0492_ _0558_ _2052_ _2053_ _2054_ vssd1 vssd1 vccd1 vccd1 _2055_ sky130_fd_sc_hd__o2111a_1
X_4503_ _0776_ _3318_ vssd1 vssd1 vccd1 vccd1 _1014_ sky130_fd_sc_hd__or2_1
X_5483_ _3262_ egd_top.BitStream_buffer.BS_buffer\[84\] vssd1 vssd1 vccd1 vccd1 _1986_
+ sky130_fd_sc_hd__nand2_1
X_4434_ _0377_ _0869_ vssd1 vssd1 vccd1 vccd1 _0945_ sky130_fd_sc_hd__nand2_1
X_4365_ _0407_ _0396_ _0399_ _0642_ _0876_ vssd1 vssd1 vccd1 vccd1 _0877_ sky130_fd_sc_hd__a221oi_1
X_6104_ _2533_ _3238_ vssd1 vssd1 vccd1 vccd1 _2535_ sky130_fd_sc_hd__nand2_1
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6035_ _2494_ _0940_ vssd1 vssd1 vccd1 vccd1 _2495_ sky130_fd_sc_hd__nand2_1
X_4296_ egd_top.BitStream_buffer.BS_buffer\[110\] vssd1 vssd1 vccd1 vccd1 _0808_ sky130_fd_sc_hd__inv_2
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6557__101 clknet_1_0__leaf__2886_ vssd1 vssd1 vccd1 vccd1 net135 sky130_fd_sc_hd__inv_2
X_5819_ _3262_ _0772_ vssd1 vssd1 vccd1 vccd1 _2319_ sky130_fd_sc_hd__nand2_1
X_6799_ net43 _0258_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_41_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4150_ egd_top.BitStream_buffer.BS_buffer\[64\] vssd1 vssd1 vccd1 vccd1 _0663_ sky130_fd_sc_hd__inv_2
X_4081_ _3045_ _0556_ vssd1 vssd1 vccd1 vccd1 _0595_ sky130_fd_sc_hd__nand2_2
XFILLER_36_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4983_ _0470_ _3237_ vssd1 vssd1 vccd1 vccd1 _1490_ sky130_fd_sc_hd__nand2_1
XFILLER_23_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3934_ _0447_ vssd1 vssd1 vccd1 vccd1 _0448_ sky130_fd_sc_hd__clkinv_2
X_6722_ net126 _0181_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.pc_previous\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_23_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3865_ egd_top.BitStream_buffer.BS_buffer\[41\] vssd1 vssd1 vccd1 vccd1 _0379_ sky130_fd_sc_hd__clkbuf_4
X_5604_ _0581_ _0515_ vssd1 vssd1 vccd1 vccd1 _2106_ sky130_fd_sc_hd__nand2_1
X_3796_ _3329_ vssd1 vssd1 vccd1 vccd1 _3330_ sky130_fd_sc_hd__buf_2
XFILLER_11_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5535_ _2027_ _2030_ _2034_ _2037_ vssd1 vssd1 vccd1 vccd1 _2038_ sky130_fd_sc_hd__and4_1
X_5466_ _0727_ _3055_ _1966_ _1967_ _1968_ vssd1 vssd1 vccd1 vccd1 _1969_ sky130_fd_sc_hd__o2111a_1
X_4417_ _0896_ _0928_ vssd1 vssd1 vccd1 vccd1 _0929_ sky130_fd_sc_hd__nor2_1
X_5397_ _0842_ _3260_ _1900_ vssd1 vssd1 vccd1 vccd1 _1901_ sky130_fd_sc_hd__o21ai_1
X_4348_ _0826_ _0859_ vssd1 vssd1 vccd1 vccd1 _0860_ sky130_fd_sc_hd__nor2_1
XFILLER_86_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4279_ egd_top.BitStream_buffer.BS_buffer\[1\] vssd1 vssd1 vccd1 vccd1 _0792_ sky130_fd_sc_hd__clkbuf_4
XTAP_193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6018_ _3020_ _2466_ _2474_ _2483_ vssd1 vssd1 vccd1 vccd1 _0249_ sky130_fd_sc_hd__o211a_1
XFILLER_36_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6611__150 clknet_1_0__leaf__2891_ vssd1 vssd1 vccd1 vccd1 net184 sky130_fd_sc_hd__inv_2
XFILLER_77_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__2890_ clknet_0__2890_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__2890_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_18_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3650_ _2931_ _3134_ vssd1 vssd1 vccd1 vccd1 _3184_ sky130_fd_sc_hd__and2_1
XFILLER_9_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3581_ _3114_ vssd1 vssd1 vccd1 vccd1 _3115_ sky130_fd_sc_hd__inv_2
X_5320_ _1809_ _1824_ vssd1 vssd1 vccd1 vccd1 _1825_ sky130_fd_sc_hd__nand2_1
XFILLER_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5251_ _3067_ _0568_ _3142_ vssd1 vssd1 vccd1 vccd1 _1756_ sky130_fd_sc_hd__and3_1
X_4202_ _3099_ _0714_ vssd1 vssd1 vccd1 vccd1 _0715_ sky130_fd_sc_hd__nand2_1
X_6696__67 clknet_1_1__leaf__2899_ vssd1 vssd1 vccd1 vccd1 net101 sky130_fd_sc_hd__inv_2
X_5182_ _0611_ _0571_ vssd1 vssd1 vccd1 vccd1 _1688_ sky130_fd_sc_hd__or2_1
XFILLER_68_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4133_ _0632_ _0636_ _0641_ _0645_ vssd1 vssd1 vccd1 vccd1 _0646_ sky130_fd_sc_hd__and4_1
X_4064_ _0577_ vssd1 vssd1 vccd1 vccd1 _0578_ sky130_fd_sc_hd__buf_4
XFILLER_91_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4966_ _0388_ _0948_ vssd1 vssd1 vccd1 vccd1 _1473_ sky130_fd_sc_hd__nand2_1
X_6705_ net109 _0164_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[92\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_51_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3917_ _0430_ vssd1 vssd1 vccd1 vccd1 _0431_ sky130_fd_sc_hd__clkbuf_2
X_4897_ _0850_ _3319_ _1402_ _1403_ _1404_ vssd1 vssd1 vccd1 vccd1 _1405_ sky130_fd_sc_hd__o2111a_1
XFILLER_51_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3848_ _0361_ vssd1 vssd1 vccd1 vccd1 _0362_ sky130_fd_sc_hd__clkbuf_2
X_3779_ _3289_ _3091_ vssd1 vssd1 vccd1 vccd1 _3313_ sky130_fd_sc_hd__nor2_2
X_5518_ _0406_ _0461_ vssd1 vssd1 vccd1 vccd1 _2021_ sky130_fd_sc_hd__nand2_1
X_6498_ _2857_ _2681_ _2859_ vssd1 vssd1 vccd1 vccd1 _2860_ sky130_fd_sc_hd__nand3_2
X_5449_ _3294_ _3338_ vssd1 vssd1 vccd1 vccd1 _1952_ sky130_fd_sc_hd__nand2_1
XFILLER_86_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4820_ _1318_ _1322_ _1324_ _1328_ vssd1 vssd1 vccd1 vccd1 _1329_ sky130_fd_sc_hd__and4_1
XFILLER_33_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_299 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4751_ _3232_ egd_top.BitStream_buffer.BS_buffer\[71\] vssd1 vssd1 vccd1 vccd1 _1260_
+ sky130_fd_sc_hd__nand2_1
X_4682_ _3168_ _3204_ vssd1 vssd1 vccd1 vccd1 _1192_ sky130_fd_sc_hd__nand2_1
X_3702_ _3235_ vssd1 vssd1 vccd1 vccd1 _3236_ sky130_fd_sc_hd__clkbuf_4
X_3633_ _3166_ vssd1 vssd1 vccd1 vccd1 _3167_ sky130_fd_sc_hd__buf_2
X_6421_ _2769_ _2765_ _2789_ vssd1 vssd1 vccd1 vccd1 _2790_ sky130_fd_sc_hd__nand3_1
X_6618__156 clknet_1_0__leaf__2892_ vssd1 vssd1 vccd1 vccd1 net190 sky130_fd_sc_hd__inv_2
X_3564_ _3041_ _3097_ vssd1 vssd1 vccd1 vccd1 _3098_ sky130_fd_sc_hd__nor2_2
X_6352_ _2678_ vssd1 vssd1 vccd1 vccd1 _2723_ sky130_fd_sc_hd__buf_6
X_5303_ _0347_ _0539_ _0375_ _0542_ _1807_ vssd1 vssd1 vccd1 vccd1 _1808_ sky130_fd_sc_hd__a221oi_1
X_3495_ _2929_ _2921_ vssd1 vssd1 vccd1 vccd1 _3029_ sky130_fd_sc_hd__nand2_1
X_6283_ _2653_ _2634_ vssd1 vssd1 vccd1 vccd1 _2654_ sky130_fd_sc_hd__nand2_1
X_5234_ _3254_ egd_top.BitStream_buffer.BS_buffer\[84\] vssd1 vssd1 vccd1 vccd1 _1739_
+ sky130_fd_sc_hd__nand2_1
X_5165_ _3221_ _0477_ _3227_ _2936_ _1670_ vssd1 vssd1 vccd1 vccd1 _1671_ sky130_fd_sc_hd__a221oi_1
XFILLER_68_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4116_ egd_top.BitStream_buffer.BS_buffer\[40\] vssd1 vssd1 vccd1 vccd1 _0629_ sky130_fd_sc_hd__inv_2
XFILLER_83_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5096_ egd_top.BitStream_buffer.BS_buffer\[0\] vssd1 vssd1 vccd1 vccd1 _1602_ sky130_fd_sc_hd__clkinv_2
XFILLER_83_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4047_ _0560_ vssd1 vssd1 vccd1 vccd1 _0561_ sky130_fd_sc_hd__buf_2
X_5998_ _2471_ _0986_ vssd1 vssd1 vccd1 vccd1 _2473_ sky130_fd_sc_hd__nand2_1
X_4949_ _1453_ _1454_ _1455_ _1456_ vssd1 vssd1 vccd1 vccd1 _1457_ sky130_fd_sc_hd__and4_1
XFILLER_20_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6675__48 clknet_1_1__leaf__2897_ vssd1 vssd1 vccd1 vccd1 net82 sky130_fd_sc_hd__inv_2
XFILLER_87_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_98 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5921_ _0602_ _0595_ vssd1 vssd1 vccd1 vccd1 _2421_ sky130_fd_sc_hd__or2_1
XFILLER_65_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5852_ _0804_ _0326_ _2351_ vssd1 vssd1 vccd1 vccd1 _2352_ sky130_fd_sc_hd__o21ai_1
X_4803_ _0633_ _0546_ _1311_ vssd1 vssd1 vccd1 vccd1 _1312_ sky130_fd_sc_hd__o21ai_1
X_5783_ _3317_ _3260_ _2283_ vssd1 vssd1 vccd1 vccd1 _2284_ sky130_fd_sc_hd__o21ai_1
XFILLER_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4734_ _3140_ egd_top.BitStream_buffer.BS_buffer\[0\] vssd1 vssd1 vccd1 vccd1 _1243_
+ sky130_fd_sc_hd__nand2_1
XFILLER_9_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4665_ _3100_ _3054_ _3061_ _0714_ vssd1 vssd1 vccd1 vccd1 _1175_ sky130_fd_sc_hd__a22o_1
X_3616_ _3148_ _3149_ vssd1 vssd1 vccd1 vccd1 _3150_ sky130_fd_sc_hd__nand2_1
X_6404_ _2629_ _2723_ _2772_ vssd1 vssd1 vccd1 vccd1 _2773_ sky130_fd_sc_hd__o21ai_1
X_4596_ egd_top.BitStream_buffer.BS_buffer\[54\] _0414_ _0418_ egd_top.BitStream_buffer.BS_buffer\[55\]
+ vssd1 vssd1 vccd1 vccd1 _1106_ sky130_fd_sc_hd__a22o_1
X_3547_ _3080_ vssd1 vssd1 vccd1 vccd1 _3081_ sky130_fd_sc_hd__buf_4
X_6335_ _2624_ _0933_ _2662_ vssd1 vssd1 vccd1 vccd1 _2706_ sky130_fd_sc_hd__or3_1
X_6266_ _2636_ vssd1 vssd1 vccd1 vccd1 _2637_ sky130_fd_sc_hd__clkinv_4
X_3478_ _2989_ _3015_ vssd1 vssd1 vccd1 vccd1 _3016_ sky130_fd_sc_hd__nand2_1
XFILLER_69_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6197_ _2592_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.pc\[4\] sky130_fd_sc_hd__buf_2
X_5217_ _3291_ _3327_ vssd1 vssd1 vccd1 vccd1 _1722_ sky130_fd_sc_hd__nand2_1
X_5148_ _0389_ _0360_ _0363_ _0869_ _1653_ vssd1 vssd1 vccd1 vccd1 _1654_ sky130_fd_sc_hd__a221oi_2
XFILLER_56_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5079_ egd_top.BitStream_buffer.BitStream_buffer_output\[8\] vssd1 vssd1 vccd1 vccd1
+ _1586_ sky130_fd_sc_hd__inv_2
XFILLER_25_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4450_ _0879_ _0424_ vssd1 vssd1 vccd1 vccd1 _0961_ sky130_fd_sc_hd__or2_1
X_4381_ _3238_ _2935_ _0892_ vssd1 vssd1 vccd1 vccd1 _0893_ sky130_fd_sc_hd__o21ai_1
X_3401_ _2952_ _2953_ _2954_ _2951_ vssd1 vssd1 vccd1 vccd1 _2955_ sky130_fd_sc_hd__o31ai_1
X_6120_ _2538_ _3257_ vssd1 vssd1 vccd1 vccd1 _2544_ sky130_fd_sc_hd__nand2_1
X_6639__15 clknet_1_1__leaf__2894_ vssd1 vssd1 vccd1 vccd1 net49 sky130_fd_sc_hd__inv_2
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6654__29 clknet_1_1__leaf__2895_ vssd1 vssd1 vccd1 vccd1 net63 sky130_fd_sc_hd__inv_2
X_6051_ _3011_ _2489_ _2501_ _2503_ vssd1 vssd1 vccd1 vccd1 _0236_ sky130_fd_sc_hd__o211a_1
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5002_ _0688_ _0558_ _1506_ _1507_ _1508_ vssd1 vssd1 vccd1 vccd1 _1509_ sky130_fd_sc_hd__o2111a_1
XFILLER_38_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5904_ _0514_ _0337_ vssd1 vssd1 vccd1 vccd1 _2404_ sky130_fd_sc_hd__nand2_1
XFILLER_53_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5835_ _3073_ egd_top.BitStream_buffer.BS_buffer\[123\] vssd1 vssd1 vccd1 vccd1 _2335_
+ sky130_fd_sc_hd__nand2_1
XFILLER_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5766_ _3168_ _3177_ vssd1 vssd1 vccd1 vccd1 _2267_ sky130_fd_sc_hd__nand2_1
X_4717_ _3085_ _3056_ _1223_ _1224_ _1225_ vssd1 vssd1 vccd1 vccd1 _1226_ sky130_fd_sc_hd__o2111a_1
X_5697_ _0965_ _0385_ _2197_ vssd1 vssd1 vccd1 vccd1 _2198_ sky130_fd_sc_hd__o21ai_1
XFILLER_30_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4648_ egd_top.BitStream_buffer.BS_buffer\[84\] vssd1 vssd1 vccd1 vccd1 _1158_ sky130_fd_sc_hd__inv_2
XFILLER_30_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4579_ _0387_ egd_top.BitStream_buffer.BS_buffer\[46\] vssd1 vssd1 vccd1 vccd1 _1089_
+ sky130_fd_sc_hd__nand2_1
X_6318_ _2629_ _2688_ _2637_ vssd1 vssd1 vccd1 vccd1 _2689_ sky130_fd_sc_hd__a21oi_1
XFILLER_1_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6249_ _2601_ _0854_ vssd1 vssd1 vccd1 vccd1 _2621_ sky130_fd_sc_hd__nand2_1
XFILLER_39_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3950_ _0463_ vssd1 vssd1 vccd1 vccd1 _0464_ sky130_fd_sc_hd__buf_2
XFILLER_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3881_ _0394_ vssd1 vssd1 vccd1 vccd1 _0395_ sky130_fd_sc_hd__clkbuf_2
XFILLER_84_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5620_ _0507_ _0365_ vssd1 vssd1 vccd1 vccd1 _2122_ sky130_fd_sc_hd__nand2_1
X_5551_ _0685_ _0571_ vssd1 vssd1 vccd1 vccd1 _2054_ sky130_fd_sc_hd__or2_1
X_4502_ _3309_ _0780_ vssd1 vssd1 vccd1 vccd1 _1013_ sky130_fd_sc_hd__nand2_1
X_5482_ _3254_ _3311_ vssd1 vssd1 vccd1 vccd1 _1985_ sky130_fd_sc_hd__nand2_1
X_4433_ _0385_ vssd1 vssd1 vccd1 vccd1 _0944_ sky130_fd_sc_hd__inv_2
X_4364_ _0420_ _0403_ _0875_ vssd1 vssd1 vccd1 vccd1 _0876_ sky130_fd_sc_hd__o21ai_1
X_4295_ _3066_ _3113_ _3117_ _3070_ _0806_ vssd1 vssd1 vccd1 vccd1 _0807_ sky130_fd_sc_hd__a221oi_1
X_6103_ _2966_ _2532_ _2528_ _2534_ vssd1 vssd1 vccd1 vccd1 _0215_ sky130_fd_sc_hd__o211a_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6034_ _2486_ vssd1 vssd1 vccd1 vccd1 _2494_ sky130_fd_sc_hd__buf_2
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6798_ net42 _0257_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_5818_ _3250_ egd_top.BitStream_buffer.BS_buffer\[88\] vssd1 vssd1 vccd1 vccd1 _2318_
+ sky130_fd_sc_hd__nand2_1
X_5749_ _1035_ _3056_ _2249_ vssd1 vssd1 vccd1 vccd1 _2250_ sky130_fd_sc_hd__o21ai_1
XFILLER_10_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_25 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4080_ egd_top.BitStream_buffer.BS_buffer\[1\] vssd1 vssd1 vccd1 vccd1 _0594_ sky130_fd_sc_hd__inv_2
XFILLER_83_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4982_ _0663_ _0464_ _1486_ _1487_ _1488_ vssd1 vssd1 vccd1 vccd1 _1489_ sky130_fd_sc_hd__o2111a_1
XFILLER_23_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6721_ net125 _0180_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.pc_previous\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_3933_ egd_top.BitStream_buffer.BS_buffer\[59\] vssd1 vssd1 vccd1 vccd1 _0447_ sky130_fd_sc_hd__clkbuf_4
X_3864_ _0377_ vssd1 vssd1 vccd1 vccd1 _0378_ sky130_fd_sc_hd__buf_2
X_5603_ _0577_ _0502_ vssd1 vssd1 vccd1 vccd1 _2105_ sky130_fd_sc_hd__nand2_1
X_3795_ _3121_ _3297_ vssd1 vssd1 vccd1 vccd1 _3329_ sky130_fd_sc_hd__nand2_2
X_5534_ _3264_ _0477_ _3248_ _2936_ _2036_ vssd1 vssd1 vccd1 vccd1 _2037_ sky130_fd_sc_hd__a221oi_1
X_5465_ _3060_ _3075_ vssd1 vssd1 vccd1 vccd1 _1968_ sky130_fd_sc_hd__nand2_1
X_4416_ _0911_ _0927_ vssd1 vssd1 vccd1 vccd1 _0928_ sky130_fd_sc_hd__nand2_1
X_5396_ _3263_ _3293_ vssd1 vssd1 vccd1 vccd1 _1900_ sky130_fd_sc_hd__nand2_1
X_6587__128 clknet_1_1__leaf__2889_ vssd1 vssd1 vccd1 vccd1 net162 sky130_fd_sc_hd__inv_2
X_4347_ _0841_ _0858_ vssd1 vssd1 vccd1 vccd1 _0859_ sky130_fd_sc_hd__nand2_1
X_4278_ _0750_ _0790_ vssd1 vssd1 vccd1 vccd1 _0791_ sky130_fd_sc_hd__nor2_1
X_6017_ _2464_ _0702_ vssd1 vssd1 vccd1 vccd1 _2483_ sky130_fd_sc_hd__nand2_1
XTAP_194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_98 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_278 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_470 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3580_ _3057_ _3031_ egd_top.BitStream_buffer.pc\[3\] vssd1 vssd1 vccd1 vccd1 _3114_
+ sky130_fd_sc_hd__and3_4
X_5250_ _1076_ _3137_ _3141_ _0566_ vssd1 vssd1 vccd1 vccd1 _1755_ sky130_fd_sc_hd__a22o_1
XFILLER_5_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4201_ egd_top.BitStream_buffer.BS_buffer\[103\] vssd1 vssd1 vccd1 vccd1 _0714_ sky130_fd_sc_hd__clkbuf_4
X_5181_ _0561_ egd_top.BitStream_buffer.BS_buffer\[14\] vssd1 vssd1 vccd1 vccd1 _1687_
+ sky130_fd_sc_hd__nand2_1
X_4132_ egd_top.BitStream_buffer.BS_buffer\[45\] _0395_ _0398_ egd_top.BitStream_buffer.BS_buffer\[46\]
+ _0644_ vssd1 vssd1 vccd1 vccd1 _0645_ sky130_fd_sc_hd__a221oi_2
XFILLER_68_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4063_ _0559_ _3125_ vssd1 vssd1 vccd1 vccd1 _0577_ sky130_fd_sc_hd__nor2_2
XFILLER_3_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4965_ _0379_ _0360_ _0363_ _0389_ _1471_ vssd1 vssd1 vccd1 vccd1 _1472_ sky130_fd_sc_hd__a221oi_1
XFILLER_24_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6704_ net108 _0163_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[93\]
+ sky130_fd_sc_hd__dfxtp_1
X_3916_ _3096_ _2933_ vssd1 vssd1 vccd1 vccd1 _0430_ sky130_fd_sc_hd__and2_1
XFILLER_51_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4896_ _0324_ _3307_ vssd1 vssd1 vccd1 vccd1 _1404_ sky130_fd_sc_hd__or2_1
X_3847_ _3058_ _0338_ vssd1 vssd1 vccd1 vccd1 _0361_ sky130_fd_sc_hd__and2_1
XFILLER_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6635_ clknet_1_1__leaf__2882_ vssd1 vssd1 vccd1 vccd1 _2894_ sky130_fd_sc_hd__buf_1
X_3778_ _3310_ _3311_ vssd1 vssd1 vccd1 vccd1 _3312_ sky130_fd_sc_hd__nand2_1
X_6526__72 clknet_1_0__leaf__2884_ vssd1 vssd1 vccd1 vccd1 net106 sky130_fd_sc_hd__inv_2
X_5517_ _0655_ _0388_ _0429_ _0944_ _2019_ vssd1 vssd1 vccd1 vccd1 _2020_ sky130_fd_sc_hd__a221oi_1
X_6497_ _2802_ _2853_ _2858_ vssd1 vssd1 vccd1 vccd1 _2859_ sky130_fd_sc_hd__nand3_1
X_6541__86 clknet_1_0__leaf__2885_ vssd1 vssd1 vccd1 vccd1 net120 sky130_fd_sc_hd__inv_2
X_5448_ _3291_ _0785_ vssd1 vssd1 vccd1 vccd1 _1951_ sky130_fd_sc_hd__nand2_1
X_5379_ _1872_ _1876_ _1878_ _1882_ vssd1 vssd1 vccd1 vccd1 _1883_ sky130_fd_sc_hd__and4_1
XFILLER_59_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4750_ _3242_ _3217_ vssd1 vssd1 vccd1 vccd1 _1259_ sky130_fd_sc_hd__nand2_1
X_4681_ _3163_ _0746_ vssd1 vssd1 vccd1 vccd1 _1191_ sky130_fd_sc_hd__nand2_1
X_3701_ _3234_ vssd1 vssd1 vccd1 vccd1 _3235_ sky130_fd_sc_hd__clkbuf_2
X_3632_ _3033_ _3134_ vssd1 vssd1 vccd1 vccd1 _3166_ sky130_fd_sc_hd__and2_1
X_6420_ _2788_ _2684_ vssd1 vssd1 vccd1 vccd1 _2789_ sky130_fd_sc_hd__nand2_1
X_6351_ _2707_ _2721_ vssd1 vssd1 vccd1 vccd1 _2722_ sky130_fd_sc_hd__nor2_1
X_5302_ _1276_ _0546_ _1806_ vssd1 vssd1 vccd1 vccd1 _1807_ sky130_fd_sc_hd__o21ai_1
X_3563_ _3096_ vssd1 vssd1 vccd1 vccd1 _3097_ sky130_fd_sc_hd__inv_2
X_6282_ _2652_ _2635_ vssd1 vssd1 vccd1 vccd1 _2653_ sky130_fd_sc_hd__nand2_1
XFILLER_5_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3494_ egd_top.BitStream_buffer.BS_buffer\[96\] vssd1 vssd1 vccd1 vccd1 _3028_ sky130_fd_sc_hd__clkbuf_4
X_5233_ _3251_ _3293_ vssd1 vssd1 vccd1 vccd1 _1738_ sky130_fd_sc_hd__nand2_1
X_5164_ _1360_ _0472_ _1669_ vssd1 vssd1 vccd1 vccd1 _1670_ sky130_fd_sc_hd__o21ai_1
XFILLER_56_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4115_ egd_top.BitStream_buffer.BitStream_buffer_output\[14\] _2965_ _0627_ vssd1
+ vssd1 vccd1 vccd1 _0628_ sky130_fd_sc_hd__o21ai_1
X_5095_ _1590_ _1594_ _1597_ _1600_ vssd1 vssd1 vccd1 vccd1 _1601_ sky130_fd_sc_hd__and4_1
XFILLER_68_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_326 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4046_ _0559_ _3097_ vssd1 vssd1 vccd1 vccd1 _0560_ sky130_fd_sc_hd__nor2_2
XFILLER_83_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5997_ _2988_ _2465_ _2458_ _2472_ vssd1 vssd1 vccd1 vccd1 _0259_ sky130_fd_sc_hd__o211a_1
X_4948_ _3144_ egd_top.BitStream_buffer.BS_buffer\[126\] vssd1 vssd1 vccd1 vccd1 _1456_
+ sky130_fd_sc_hd__nand2_1
X_4879_ _0543_ _0512_ _1384_ _1385_ _1386_ vssd1 vssd1 vccd1 vccd1 _1387_ sky130_fd_sc_hd__o2111a_1
XFILLER_3_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_66 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5920_ _0528_ _0576_ _2417_ _2418_ _2419_ vssd1 vssd1 vccd1 vccd1 _2420_ sky130_fd_sc_hd__o2111a_1
XFILLER_80_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5851_ _0328_ _3109_ vssd1 vssd1 vccd1 vccd1 _2351_ sky130_fd_sc_hd__nand2_1
X_4802_ _0548_ _0365_ vssd1 vssd1 vccd1 vccd1 _1311_ sky130_fd_sc_hd__nand2_1
X_5782_ _3263_ _3311_ vssd1 vssd1 vccd1 vccd1 _2283_ sky130_fd_sc_hd__nand2_1
X_4733_ _0597_ _3182_ _1239_ _1240_ _1241_ vssd1 vssd1 vccd1 vccd1 _1242_ sky130_fd_sc_hd__o2111a_1
X_4664_ _1157_ _1173_ vssd1 vssd1 vccd1 vccd1 _1174_ sky130_fd_sc_hd__nand2_1
X_6403_ _2723_ egd_top.BitStream_buffer.BitStream_buffer_output\[6\] vssd1 vssd1 vccd1
+ vccd1 _2772_ sky130_fd_sc_hd__nand2_1
X_3615_ egd_top.BitStream_buffer.BS_buffer\[121\] vssd1 vssd1 vccd1 vccd1 _3149_ sky130_fd_sc_hd__buf_2
X_4595_ _0960_ _0424_ _0437_ _0421_ vssd1 vssd1 vccd1 vccd1 _1105_ sky130_fd_sc_hd__o22ai_1
X_3546_ _3041_ _3079_ vssd1 vssd1 vccd1 vccd1 _3080_ sky130_fd_sc_hd__nor2_4
X_6334_ _2703_ _2704_ _2669_ vssd1 vssd1 vccd1 vccd1 _2705_ sky130_fd_sc_hd__a21o_1
X_6265_ _2634_ _2635_ _1586_ vssd1 vssd1 vccd1 vccd1 _2636_ sky130_fd_sc_hd__and3_1
X_5216_ _1709_ _1712_ _1716_ _1720_ vssd1 vssd1 vccd1 vccd1 _1721_ sky130_fd_sc_hd__and4_1
X_3477_ egd_top.BitStream_buffer.BS_buffer\[124\] vssd1 vssd1 vccd1 vccd1 _3015_ sky130_fd_sc_hd__clkinv_2
X_6196_ _2591_ _2586_ vssd1 vssd1 vccd1 vccd1 _2592_ sky130_fd_sc_hd__and2_1
XFILLER_84_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5147_ _0861_ _0368_ _1652_ vssd1 vssd1 vccd1 vccd1 _1653_ sky130_fd_sc_hd__o21ai_1
XFILLER_28_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5078_ _1522_ _1583_ _1584_ vssd1 vssd1 vccd1 vccd1 _1585_ sky130_fd_sc_hd__nand3_1
XFILLER_28_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6680__52 clknet_1_1__leaf__2898_ vssd1 vssd1 vccd1 vccd1 net86 sky130_fd_sc_hd__inv_2
X_4029_ egd_top.BitStream_buffer.BS_buffer\[29\] vssd1 vssd1 vccd1 vccd1 _0543_ sky130_fd_sc_hd__inv_2
XFILLER_25_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4380_ _0477_ _3244_ vssd1 vssd1 vccd1 vccd1 _0892_ sky130_fd_sc_hd__nand2_1
X_3400_ net30 net29 vssd1 vssd1 vccd1 vccd1 _2954_ sky130_fd_sc_hd__nor2_1
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6050_ _2494_ _0383_ vssd1 vssd1 vccd1 vccd1 _2503_ sky130_fd_sc_hd__nand2_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5001_ _0676_ _0571_ vssd1 vssd1 vccd1 vccd1 _1508_ sky130_fd_sc_hd__or2_1
XFILLER_78_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5903_ _0537_ _0487_ _0540_ _0490_ _2402_ vssd1 vssd1 vccd1 vccd1 _2403_ sky130_fd_sc_hd__a221oi_1
XFILLER_53_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5834_ _2999_ _3122_ _2331_ _2332_ _2333_ vssd1 vssd1 vccd1 vccd1 _2334_ sky130_fd_sc_hd__o2111a_1
X_5765_ _3163_ _0741_ vssd1 vssd1 vccd1 vccd1 _2266_ sky130_fd_sc_hd__nand2_1
X_4716_ _3048_ _3100_ vssd1 vssd1 vccd1 vccd1 _1225_ sky130_fd_sc_hd__nand2_1
X_5696_ _0387_ _0436_ vssd1 vssd1 vccd1 vccd1 _2197_ sky130_fd_sc_hd__nand2_1
X_4647_ _1143_ _1148_ _1152_ _1156_ vssd1 vssd1 vccd1 vccd1 _1157_ sky130_fd_sc_hd__and4_1
X_4578_ _1084_ _0367_ _1085_ _1086_ _1087_ vssd1 vssd1 vccd1 vccd1 _1088_ sky130_fd_sc_hd__o2111a_1
X_6317_ egd_top.BitStream_buffer.BitStream_buffer_output\[7\] _2687_ vssd1 vssd1 vccd1
+ vccd1 _2688_ sky130_fd_sc_hd__nor2_1
X_3529_ _3061_ _3062_ vssd1 vssd1 vccd1 vccd1 _3063_ sky130_fd_sc_hd__nand2_1
X_6248_ _3020_ _2603_ _2611_ _2620_ vssd1 vssd1 vccd1 vccd1 _0162_ sky130_fd_sc_hd__o211a_1
X_6179_ _2925_ _2578_ _2577_ vssd1 vssd1 vccd1 vccd1 _2579_ sky130_fd_sc_hd__o21ai_2
XFILLER_69_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_424 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3880_ _3067_ _0338_ vssd1 vssd1 vccd1 vccd1 _0394_ sky130_fd_sc_hd__and2_1
X_5550_ _0565_ egd_top.BitStream_buffer.BS_buffer\[15\] vssd1 vssd1 vccd1 vccd1 _2053_
+ sky130_fd_sc_hd__nand2_1
XFILLER_77_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5481_ _1149_ _3240_ _1981_ _1982_ _1983_ vssd1 vssd1 vccd1 vccd1 _1984_ sky130_fd_sc_hd__o2111a_1
X_4501_ _3313_ egd_top.BitStream_buffer.BS_buffer\[87\] vssd1 vssd1 vccd1 vccd1 _1012_
+ sky130_fd_sc_hd__nand2_1
X_4432_ _0346_ _0359_ _0362_ _0354_ _0942_ vssd1 vssd1 vccd1 vccd1 _0943_ sky130_fd_sc_hd__a221oi_1
X_4363_ _0406_ _0874_ vssd1 vssd1 vccd1 vccd1 _0875_ sky130_fd_sc_hd__nand2_1
X_4294_ _0804_ _3123_ _0805_ vssd1 vssd1 vccd1 vccd1 _0806_ sky130_fd_sc_hd__o21ai_1
X_6102_ _2533_ _0663_ vssd1 vssd1 vccd1 vccd1 _2534_ sky130_fd_sc_hd__nand2_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6033_ _2985_ _2487_ _2488_ _2493_ vssd1 vssd1 vccd1 vccd1 _0244_ sky130_fd_sc_hd__o211a_1
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5817_ _3322_ _3271_ _3327_ _3275_ _2316_ vssd1 vssd1 vccd1 vccd1 _2317_ sky130_fd_sc_hd__a221oi_1
XFILLER_10_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6797_ net41 _0256_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_5748_ _3061_ _3169_ vssd1 vssd1 vccd1 vccd1 _2249_ sky130_fd_sc_hd__nand2_1
XFILLER_41_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5679_ _3074_ _3149_ vssd1 vssd1 vccd1 vccd1 _2181_ sky130_fd_sc_hd__nand2_1
XFILLER_1_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6564__107 clknet_1_0__leaf__2887_ vssd1 vssd1 vccd1 vccd1 net141 sky130_fd_sc_hd__inv_2
XFILLER_66_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__2889_ clknet_0__2889_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__2889_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_48_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4981_ _1297_ _0450_ vssd1 vssd1 vccd1 vccd1 _1488_ sky130_fd_sc_hd__or2_1
X_6720_ net124 _0179_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.pc_previous\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_16_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3932_ _0429_ _0432_ _0435_ _0436_ _0445_ vssd1 vssd1 vccd1 vccd1 _0446_ sky130_fd_sc_hd__a221oi_1
XFILLER_51_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3863_ _0376_ vssd1 vssd1 vccd1 vccd1 _0377_ sky130_fd_sc_hd__clkbuf_2
X_5602_ _0692_ _0557_ _2101_ _2102_ _2103_ vssd1 vssd1 vccd1 vccd1 _2104_ sky130_fd_sc_hd__o2111a_1
XFILLER_31_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5533_ _3257_ _0472_ _2035_ vssd1 vssd1 vccd1 vccd1 _2036_ sky130_fd_sc_hd__o21ai_1
X_3794_ egd_top.BitStream_buffer.BS_buffer\[89\] vssd1 vssd1 vccd1 vccd1 _3328_ sky130_fd_sc_hd__clkinv_2
X_5464_ _3047_ _3066_ vssd1 vssd1 vccd1 vccd1 _1967_ sky130_fd_sc_hd__nand2_1
X_4415_ _0915_ _0919_ _0921_ _0926_ vssd1 vssd1 vccd1 vccd1 _0927_ sky130_fd_sc_hd__and4_1
X_5395_ _1888_ _1891_ _1895_ _1898_ vssd1 vssd1 vccd1 vccd1 _1899_ sky130_fd_sc_hd__and4_1
X_4346_ _0845_ _0849_ _0853_ _0857_ vssd1 vssd1 vccd1 vccd1 _0858_ sky130_fd_sc_hd__and4_1
XFILLER_59_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4277_ _0766_ _0789_ vssd1 vssd1 vccd1 vccd1 _0790_ sky130_fd_sc_hd__nand2_1
XTAP_195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6016_ _3017_ _2466_ _2474_ _2482_ vssd1 vssd1 vccd1 vccd1 _0250_ sky130_fd_sc_hd__o211a_1
XFILLER_82_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_427 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6849_ net93 _0308_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[117\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_50_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4200_ egd_top.BitStream_buffer.BS_buffer\[102\] vssd1 vssd1 vccd1 vccd1 _0713_ sky130_fd_sc_hd__clkinv_2
X_5180_ _0565_ egd_top.BitStream_buffer.BS_buffer\[12\] vssd1 vssd1 vccd1 vccd1 _1686_
+ sky130_fd_sc_hd__nand2_1
XFILLER_68_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4131_ _0423_ _0402_ _0643_ vssd1 vssd1 vccd1 vccd1 _0644_ sky130_fd_sc_hd__o21ai_1
X_4062_ _0575_ vssd1 vssd1 vccd1 vccd1 _0576_ sky130_fd_sc_hd__buf_2
XFILLER_56_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4964_ _0629_ _0368_ _1470_ vssd1 vssd1 vccd1 vccd1 _1471_ sky130_fd_sc_hd__o21ai_1
XFILLER_51_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3915_ egd_top.BitStream_buffer.BS_buffer\[54\] vssd1 vssd1 vccd1 vccd1 _0429_ sky130_fd_sc_hd__clkbuf_4
X_6703_ net107 _0162_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[94\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_32_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4895_ _3309_ _0330_ vssd1 vssd1 vccd1 vccd1 _1403_ sky130_fd_sc_hd__nand2_1
X_3846_ _0359_ vssd1 vssd1 vccd1 vccd1 _0360_ sky130_fd_sc_hd__clkbuf_4
X_6593__133 clknet_1_0__leaf__2890_ vssd1 vssd1 vccd1 vccd1 net167 sky130_fd_sc_hd__inv_2
X_3777_ egd_top.BitStream_buffer.BS_buffer\[86\] vssd1 vssd1 vccd1 vccd1 _3311_ sky130_fd_sc_hd__clkbuf_4
X_6496_ _2856_ _2635_ vssd1 vssd1 vccd1 vccd1 _2858_ sky130_fd_sc_hd__nand2_1
X_5516_ _0960_ _0380_ _2018_ vssd1 vssd1 vccd1 vccd1 _2019_ sky130_fd_sc_hd__o21ai_1
X_5447_ _0716_ _3324_ _3326_ _3100_ _1949_ vssd1 vssd1 vccd1 vccd1 _1950_ sky130_fd_sc_hd__a221oi_1
X_5378_ _0528_ _0604_ _1879_ _1880_ _1881_ vssd1 vssd1 vccd1 vccd1 _1882_ sky130_fd_sc_hd__o2111a_1
X_4329_ _0828_ _0832_ _0836_ _0840_ vssd1 vssd1 vccd1 vccd1 _0841_ sky130_fd_sc_hd__and4_1
XFILLER_59_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3700_ _3058_ _3213_ vssd1 vssd1 vccd1 vccd1 _3234_ sky130_fd_sc_hd__and2_1
X_4680_ _0741_ _3137_ _3187_ _3141_ _1189_ vssd1 vssd1 vccd1 vccd1 _1190_ sky130_fd_sc_hd__a221oi_1
X_3631_ _3163_ _3164_ vssd1 vssd1 vccd1 vccd1 _3165_ sky130_fd_sc_hd__nand2_1
X_3562_ _3051_ egd_top.BitStream_buffer.pc\[2\] _3032_ vssd1 vssd1 vccd1 vccd1 _3096_
+ sky130_fd_sc_hd__and3_2
X_6350_ _2711_ _2716_ _2720_ vssd1 vssd1 vccd1 vccd1 _2721_ sky130_fd_sc_hd__nand3_1
X_5301_ _0548_ _0346_ vssd1 vssd1 vccd1 vccd1 _1806_ sky130_fd_sc_hd__nand2_1
X_6281_ _2651_ _1586_ vssd1 vssd1 vccd1 vccd1 _2652_ sky130_fd_sc_hd__nand2_1
X_3493_ _3026_ vssd1 vssd1 vccd1 vccd1 _3027_ sky130_fd_sc_hd__buf_2
XFILLER_88_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5232_ _1725_ _1729_ _1733_ _1736_ vssd1 vssd1 vccd1 vccd1 _1737_ sky130_fd_sc_hd__and4_1
X_5163_ _0470_ _3210_ vssd1 vssd1 vccd1 vccd1 _1669_ sky130_fd_sc_hd__nand2_1
X_4114_ _2904_ vssd1 vssd1 vccd1 vccd1 _0627_ sky130_fd_sc_hd__buf_2
XFILLER_83_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5094_ _3191_ _0726_ _3198_ _3081_ _1599_ vssd1 vssd1 vccd1 vccd1 _1600_ sky130_fd_sc_hd__a221oi_1
XFILLER_56_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4045_ _0556_ vssd1 vssd1 vccd1 vccd1 _0559_ sky130_fd_sc_hd__inv_2
XFILLER_17_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5996_ _2471_ _0897_ vssd1 vssd1 vccd1 vccd1 _2472_ sky130_fd_sc_hd__nand2_1
X_4947_ _3136_ egd_top.BitStream_buffer.BS_buffer\[0\] vssd1 vssd1 vccd1 vccd1 _1455_
+ sky130_fd_sc_hd__nand2_1
XFILLER_33_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4878_ _0507_ egd_top.BitStream_buffer.BS_buffer\[27\] vssd1 vssd1 vccd1 vccd1 _1386_
+ sky130_fd_sc_hd__nand2_1
X_3829_ _3104_ _0339_ vssd1 vssd1 vccd1 vccd1 _0343_ sky130_fd_sc_hd__and2_1
XFILLER_20_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6479_ _2838_ _2841_ vssd1 vssd1 vccd1 vccd1 _2842_ sky130_fd_sc_hd__nand2_1
XFILLER_58_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5850_ _2346_ _2347_ _2348_ _2349_ vssd1 vssd1 vccd1 vccd1 _2350_ sky130_fd_sc_hd__and4_1
X_4801_ _0543_ _0523_ _0907_ _0534_ _1309_ vssd1 vssd1 vccd1 vccd1 _1310_ sky130_fd_sc_hd__o221a_1
XFILLER_61_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5781_ _3276_ _3233_ _3236_ _0837_ _2281_ vssd1 vssd1 vccd1 vccd1 _2282_ sky130_fd_sc_hd__a221oi_2
X_4732_ _3185_ egd_top.BitStream_buffer.BS_buffer\[4\] vssd1 vssd1 vccd1 vccd1 _1241_
+ sky130_fd_sc_hd__nand2_1
X_4663_ _1161_ _1165_ _1168_ _1172_ vssd1 vssd1 vccd1 vccd1 _1173_ sky130_fd_sc_hd__and4_1
X_3614_ _3147_ vssd1 vssd1 vccd1 vccd1 _3148_ sky130_fd_sc_hd__buf_6
X_6402_ _2729_ _2725_ vssd1 vssd1 vccd1 vccd1 _2771_ sky130_fd_sc_hd__nor2_1
X_4594_ _0462_ _0438_ _1101_ _1102_ _1103_ vssd1 vssd1 vccd1 vccd1 _1104_ sky130_fd_sc_hd__o2111a_1
X_3545_ _2931_ vssd1 vssd1 vccd1 vccd1 _3079_ sky130_fd_sc_hd__inv_2
X_6333_ egd_top.BitStream_buffer.BitStream_buffer_output\[8\] egd_top.BitStream_buffer.BitStream_buffer_output\[7\]
+ vssd1 vssd1 vccd1 vccd1 _2704_ sky130_fd_sc_hd__nand2_1
XFILLER_88_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3476_ net10 vssd1 vssd1 vccd1 vccd1 _3014_ sky130_fd_sc_hd__buf_4
X_6264_ egd_top.BitStream_buffer.BitStream_buffer_output\[9\] vssd1 vssd1 vccd1 vccd1
+ _2635_ sky130_fd_sc_hd__clkinv_2
XFILLER_88_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5215_ _2977_ _3089_ _1717_ _1718_ _1719_ vssd1 vssd1 vccd1 vccd1 _1720_ sky130_fd_sc_hd__o2111a_1
X_6195_ egd_top.BitStream_buffer.pc_previous\[4\] _2585_ vssd1 vssd1 vccd1 vccd1 _2591_
+ sky130_fd_sc_hd__or2_1
XFILLER_84_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5146_ _0371_ _0375_ vssd1 vssd1 vccd1 vccd1 _1652_ sky130_fd_sc_hd__nand2_1
XFILLER_56_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5077_ _0622_ _0553_ vssd1 vssd1 vccd1 vccd1 _1584_ sky130_fd_sc_hd__nand2_1
XFILLER_84_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4028_ _0541_ vssd1 vssd1 vccd1 vccd1 _0542_ sky130_fd_sc_hd__buf_2
XFILLER_37_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5979_ _2441_ _0688_ vssd1 vssd1 vccd1 vccd1 _2461_ sky130_fd_sc_hd__nand2_1
XFILLER_40_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_411 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_116 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5000_ _0565_ egd_top.BitStream_buffer.BS_buffer\[11\] vssd1 vssd1 vccd1 vccd1 _1507_
+ sky130_fd_sc_hd__nand2_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5902_ _0995_ _0495_ _2401_ vssd1 vssd1 vccd1 vccd1 _2402_ sky130_fd_sc_hd__o21ai_1
XFILLER_81_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5833_ _3116_ _3149_ vssd1 vssd1 vccd1 vccd1 _2333_ sky130_fd_sc_hd__nand2_1
XFILLER_22_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5764_ _0553_ _3137_ _0579_ _3141_ _2264_ vssd1 vssd1 vccd1 vccd1 _2265_ sky130_fd_sc_hd__a221oi_1
X_4715_ _3060_ egd_top.BitStream_buffer.BS_buffer\[104\] vssd1 vssd1 vccd1 vccd1 _1224_
+ sky130_fd_sc_hd__nand2_1
X_5695_ _0642_ _0359_ _0362_ _0874_ _2195_ vssd1 vssd1 vccd1 vccd1 _2196_ sky130_fd_sc_hd__a221oi_1
X_4646_ _3288_ _3282_ _3293_ _1153_ _1155_ vssd1 vssd1 vccd1 vccd1 _1156_ sky130_fd_sc_hd__a221oi_1
X_4577_ _0362_ _0347_ vssd1 vssd1 vccd1 vccd1 _1087_ sky130_fd_sc_hd__nand2_1
XFILLER_89_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6316_ _2686_ vssd1 vssd1 vccd1 vccd1 _2687_ sky130_fd_sc_hd__inv_2
XFILLER_89_536 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3528_ egd_top.BitStream_buffer.BS_buffer\[99\] vssd1 vssd1 vccd1 vccd1 _3062_ sky130_fd_sc_hd__clkbuf_4
X_3459_ net14 vssd1 vssd1 vccd1 vccd1 _3001_ sky130_fd_sc_hd__clkbuf_4
X_6247_ _2601_ _0784_ vssd1 vssd1 vccd1 vccd1 _2620_ sky130_fd_sc_hd__nand2_1
XFILLER_39_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6178_ _2576_ _2577_ vssd1 vssd1 vccd1 vccd1 _2578_ sky130_fd_sc_hd__nand2_2
XFILLER_29_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5129_ _0324_ _3319_ vssd1 vssd1 vccd1 vccd1 _1635_ sky130_fd_sc_hd__or2_1
XFILLER_84_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6644__20 clknet_1_0__leaf__2894_ vssd1 vssd1 vccd1 vccd1 net54 sky130_fd_sc_hd__inv_2
XFILLER_75_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_80 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5480_ _3235_ _3283_ vssd1 vssd1 vccd1 vccd1 _1983_ sky130_fd_sc_hd__nand2_1
X_4500_ _1007_ _3298_ _1008_ _1009_ _1010_ vssd1 vssd1 vccd1 vccd1 _1011_ sky130_fd_sc_hd__o2111a_1
X_4431_ _0940_ _0367_ _0941_ vssd1 vssd1 vccd1 vccd1 _0942_ sky130_fd_sc_hd__o21ai_1
XFILLER_6_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_1 _0256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4362_ egd_top.BitStream_buffer.BS_buffer\[48\] vssd1 vssd1 vccd1 vccd1 _0874_ sky130_fd_sc_hd__clkbuf_4
X_4293_ _3127_ _3109_ vssd1 vssd1 vccd1 vccd1 _0805_ sky130_fd_sc_hd__nand2_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6101_ _2531_ vssd1 vssd1 vccd1 vccd1 _2533_ sky130_fd_sc_hd__clkbuf_4
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6032_ _2489_ _0865_ vssd1 vssd1 vccd1 vccd1 _2493_ sky130_fd_sc_hd__nand2_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5816_ _0330_ _3281_ _1153_ _0785_ vssd1 vssd1 vccd1 vccd1 _2316_ sky130_fd_sc_hd__a22o_1
XFILLER_10_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6796_ net40 _0255_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_5747_ _2203_ _2218_ _2233_ _2247_ vssd1 vssd1 vccd1 vccd1 _2248_ sky130_fd_sc_hd__and4_1
XFILLER_10_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5678_ _3191_ _3113_ _3117_ _3198_ _2179_ vssd1 vssd1 vccd1 vccd1 _2180_ sky130_fd_sc_hd__a221oi_1
X_4629_ egd_top.BitStream_buffer.BS_buffer\[34\] _0538_ _0364_ _0541_ _1138_ vssd1
+ vssd1 vccd1 vccd1 _1139_ sky130_fd_sc_hd__a221oi_1
XFILLER_1_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__2888_ clknet_0__2888_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__2888_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_91_531 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4980_ _0458_ _0751_ vssd1 vssd1 vccd1 vccd1 _1487_ sky130_fd_sc_hd__nand2_1
X_3931_ _0437_ _0439_ _0444_ vssd1 vssd1 vccd1 vccd1 _0445_ sky130_fd_sc_hd__o21ai_1
X_3862_ _3124_ _0338_ vssd1 vssd1 vccd1 vccd1 _0376_ sky130_fd_sc_hd__and2_1
XFILLER_31_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5601_ _0922_ _0570_ vssd1 vssd1 vccd1 vccd1 _2103_ sky130_fd_sc_hd__or2_1
X_5532_ _0469_ _3227_ vssd1 vssd1 vccd1 vccd1 _2035_ sky130_fd_sc_hd__nand2_1
X_3793_ egd_top.BitStream_buffer.BS_buffer\[91\] vssd1 vssd1 vccd1 vccd1 _3327_ sky130_fd_sc_hd__clkbuf_4
X_5463_ _3038_ _3118_ vssd1 vssd1 vccd1 vccd1 _1966_ sky130_fd_sc_hd__nand2_1
X_4414_ _0922_ _0604_ _0923_ _0924_ _0925_ vssd1 vssd1 vccd1 vccd1 _0926_ sky130_fd_sc_hd__o2111a_1
X_5394_ _3128_ _3340_ _0722_ _0323_ _1897_ vssd1 vssd1 vccd1 vccd1 _1898_ sky130_fd_sc_hd__a221oi_1
X_4345_ _3028_ _3340_ _3040_ _0323_ _0856_ vssd1 vssd1 vccd1 vccd1 _0857_ sky130_fd_sc_hd__a221oi_1
X_4276_ _0770_ _0778_ _0783_ _0788_ vssd1 vssd1 vccd1 vccd1 _0789_ sky130_fd_sc_hd__and4_1
XFILLER_86_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6015_ _2471_ _0543_ vssd1 vssd1 vccd1 vccd1 _2482_ sky130_fd_sc_hd__nand2_1
XTAP_196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_439 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6848_ net92 _0307_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[118\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_10_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6779_ net183 _0238_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[41\]
+ sky130_fd_sc_hd__dfxtp_1
X_6570__112 clknet_1_0__leaf__2888_ vssd1 vssd1 vccd1 vccd1 net146 sky130_fd_sc_hd__inv_2
XFILLER_89_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4130_ _0405_ _0642_ vssd1 vssd1 vccd1 vccd1 _0643_ sky130_fd_sc_hd__nand2_1
XFILLER_3_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4061_ _3114_ _0556_ vssd1 vssd1 vccd1 vccd1 _0575_ sky130_fd_sc_hd__nand2_1
XFILLER_76_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4963_ _0371_ _0347_ vssd1 vssd1 vccd1 vccd1 _1470_ sky130_fd_sc_hd__nand2_1
XFILLER_51_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3914_ _0412_ _0415_ _0416_ _0419_ _0427_ vssd1 vssd1 vccd1 vccd1 _0428_ sky130_fd_sc_hd__a221oi_1
X_6702_ net106 _0161_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[95\]
+ sky130_fd_sc_hd__dfxtp_1
X_4894_ _3313_ _3322_ vssd1 vssd1 vccd1 vccd1 _1402_ sky130_fd_sc_hd__nand2_1
X_3845_ _0358_ vssd1 vssd1 vccd1 vccd1 _0359_ sky130_fd_sc_hd__clkbuf_2
XFILLER_22_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3776_ _3309_ vssd1 vssd1 vccd1 vccd1 _3310_ sky130_fd_sc_hd__buf_4
X_6495_ _2854_ _2635_ _2856_ vssd1 vssd1 vccd1 vccd1 _2857_ sky130_fd_sc_hd__nand3_1
X_5515_ _0377_ _0416_ vssd1 vssd1 vccd1 vccd1 _2018_ sky130_fd_sc_hd__nand2_1
X_5446_ _0796_ _3330_ _1948_ vssd1 vssd1 vccd1 vccd1 _1949_ sky130_fd_sc_hd__o21ai_1
X_6687__59 clknet_1_1__leaf__2898_ vssd1 vssd1 vccd1 vccd1 net93 sky130_fd_sc_hd__inv_2
X_5377_ _0510_ _0613_ vssd1 vssd1 vccd1 vccd1 _1881_ sky130_fd_sc_hd__or2_1
X_4328_ _3283_ _3271_ _3276_ _3275_ _0839_ vssd1 vssd1 vccd1 vccd1 _0840_ sky130_fd_sc_hd__a221oi_1
XFILLER_74_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4259_ egd_top.BitStream_buffer.BS_buffer\[87\] vssd1 vssd1 vccd1 vccd1 _0772_ sky130_fd_sc_hd__clkbuf_4
XFILLER_27_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_391 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_80 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3630_ egd_top.BitStream_buffer.BS_buffer\[113\] vssd1 vssd1 vccd1 vccd1 _3164_ sky130_fd_sc_hd__clkbuf_4
X_3561_ _3093_ _3094_ vssd1 vssd1 vccd1 vccd1 _3095_ sky130_fd_sc_hd__nand2_1
X_5300_ _0366_ _0523_ _0940_ _0526_ _1804_ vssd1 vssd1 vccd1 vccd1 _1805_ sky130_fd_sc_hd__o221a_1
XFILLER_52_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6280_ _2650_ _1705_ vssd1 vssd1 vccd1 vccd1 _2651_ sky130_fd_sc_hd__nand2_1
X_3492_ egd_top.BitStream_buffer.BitStream_buffer_valid_n vssd1 vssd1 vccd1 vccd1
+ _3026_ sky130_fd_sc_hd__buf_2
X_5231_ _0714_ _3339_ _3128_ _0322_ _1735_ vssd1 vssd1 vccd1 vccd1 _1736_ sky130_fd_sc_hd__a221oi_1
X_5162_ _0829_ _0450_ _1665_ _1666_ _1667_ vssd1 vssd1 vccd1 vccd1 _1668_ sky130_fd_sc_hd__o2111a_1
X_5093_ _2990_ _0729_ _1598_ vssd1 vssd1 vccd1 vccd1 _1599_ sky130_fd_sc_hd__o21ai_1
XFILLER_29_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4113_ _3027_ _0625_ _0626_ vssd1 vssd1 vccd1 vccd1 _0297_ sky130_fd_sc_hd__o21a_1
XFILLER_56_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4044_ _0557_ vssd1 vssd1 vccd1 vccd1 _0558_ sky130_fd_sc_hd__buf_2
XFILLER_83_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6601__141 clknet_1_1__leaf__2890_ vssd1 vssd1 vccd1 vccd1 net175 sky130_fd_sc_hd__inv_2
X_5995_ _2464_ vssd1 vssd1 vccd1 vccd1 _2471_ sky130_fd_sc_hd__buf_2
X_4946_ _3140_ egd_top.BitStream_buffer.BS_buffer\[1\] vssd1 vssd1 vccd1 vccd1 _1454_
+ sky130_fd_sc_hd__nand2_1
X_4877_ _0513_ egd_top.BitStream_buffer.BS_buffer\[28\] vssd1 vssd1 vccd1 vccd1 _1385_
+ sky130_fd_sc_hd__nand2_1
X_3828_ _0341_ vssd1 vssd1 vccd1 vccd1 _0342_ sky130_fd_sc_hd__buf_2
X_6547_ clknet_1_1__leaf__2883_ vssd1 vssd1 vccd1 vccd1 _2886_ sky130_fd_sc_hd__buf_1
X_3759_ egd_top.BitStream_buffer.BS_buffer\[83\] vssd1 vssd1 vccd1 vccd1 _3293_ sky130_fd_sc_hd__clkbuf_4
X_6478_ _2840_ vssd1 vssd1 vccd1 vccd1 _2841_ sky130_fd_sc_hd__inv_2
X_5429_ _1931_ _1932_ vssd1 vssd1 vccd1 vccd1 _1933_ sky130_fd_sc_hd__nand2_1
XFILLER_87_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4800_ _0702_ _0530_ _0995_ _0526_ vssd1 vssd1 vccd1 vccd1 _1309_ sky130_fd_sc_hd__o22a_1
XFILLER_34_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5780_ _1574_ _3240_ _2280_ vssd1 vssd1 vccd1 vccd1 _2281_ sky130_fd_sc_hd__o21ai_1
X_4731_ _3179_ _0930_ vssd1 vssd1 vccd1 vccd1 _1240_ sky130_fd_sc_hd__nand2_1
XFILLER_61_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4662_ _0708_ _3340_ _3062_ _0323_ _1171_ vssd1 vssd1 vccd1 vccd1 _1172_ sky130_fd_sc_hd__a221oi_1
X_3613_ _3146_ vssd1 vssd1 vccd1 vccd1 _3147_ sky130_fd_sc_hd__buf_6
X_6401_ _2769_ _2765_ vssd1 vssd1 vccd1 vccd1 _2770_ sky130_fd_sc_hd__nand2_1
X_4593_ _0434_ _0447_ vssd1 vssd1 vccd1 vccd1 _1103_ sky130_fd_sc_hd__nand2_1
X_3544_ _3041_ _3077_ vssd1 vssd1 vccd1 vccd1 _3078_ sky130_fd_sc_hd__nor2_2
X_6332_ _2702_ vssd1 vssd1 vccd1 vccd1 _2703_ sky130_fd_sc_hd__inv_2
X_6263_ _2633_ vssd1 vssd1 vccd1 vccd1 _2634_ sky130_fd_sc_hd__inv_2
X_3475_ _3011_ _2976_ _3002_ _3013_ vssd1 vssd1 vccd1 vccd1 _0302_ sky130_fd_sc_hd__o211a_1
XFILLER_88_217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5214_ _0808_ _3105_ vssd1 vssd1 vccd1 vccd1 _1719_ sky130_fd_sc_hd__or2_1
X_6194_ _2590_ vssd1 vssd1 vccd1 vccd1 _0182_ sky130_fd_sc_hd__inv_2
X_5145_ _0874_ _0378_ _0948_ _0382_ _1650_ vssd1 vssd1 vccd1 vccd1 _1651_ sky130_fd_sc_hd__a221oi_1
X_5076_ _1551_ _1582_ vssd1 vssd1 vccd1 vccd1 _1583_ sky130_fd_sc_hd__nor2_1
X_4027_ _0488_ _3079_ vssd1 vssd1 vccd1 vccd1 _0541_ sky130_fd_sc_hd__nor2_2
XFILLER_44_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_331 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5978_ _3017_ _2443_ _2458_ _2460_ vssd1 vssd1 vccd1 vccd1 _0266_ sky130_fd_sc_hd__o211a_1
X_4929_ _3259_ egd_top.BitStream_buffer.BS_buffer\[78\] vssd1 vssd1 vccd1 vccd1 _1437_
+ sky130_fd_sc_hd__nand2_1
XFILLER_60_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6608__147 clknet_1_1__leaf__2891_ vssd1 vssd1 vccd1 vccd1 net181 sky130_fd_sc_hd__inv_2
XFILLER_75_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5901_ _0497_ _0365_ vssd1 vssd1 vccd1 vccd1 _2401_ sky130_fd_sc_hd__nand2_1
XFILLER_19_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5832_ _3112_ _0744_ vssd1 vssd1 vccd1 vccd1 _2332_ sky130_fd_sc_hd__nand2_1
XFILLER_22_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5763_ _0569_ _3145_ _2263_ vssd1 vssd1 vccd1 vccd1 _2264_ sky130_fd_sc_hd__o21ai_1
X_4714_ _3039_ _0716_ vssd1 vssd1 vccd1 vccd1 _1223_ sky130_fd_sc_hd__nand2_1
X_5694_ _1466_ _0367_ _2194_ vssd1 vssd1 vccd1 vccd1 _2195_ sky130_fd_sc_hd__o21ai_1
X_4645_ _0767_ _3273_ _1154_ vssd1 vssd1 vccd1 vccd1 _1155_ sky130_fd_sc_hd__o21ai_1
XFILLER_30_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4576_ _0359_ _0354_ vssd1 vssd1 vccd1 vccd1 _1086_ sky130_fd_sc_hd__nand2_1
X_3527_ _3060_ vssd1 vssd1 vccd1 vccd1 _3061_ sky130_fd_sc_hd__buf_6
X_6315_ egd_top.BitStream_buffer.BitStream_buffer_output\[6\] egd_top.BitStream_buffer.BitStream_buffer_output\[5\]
+ vssd1 vssd1 vccd1 vccd1 _2686_ sky130_fd_sc_hd__nor2_1
XFILLER_89_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6246_ _3017_ _2603_ _2611_ _2619_ vssd1 vssd1 vccd1 vccd1 _0163_ sky130_fd_sc_hd__o211a_1
X_3458_ _2998_ _2975_ _2913_ _3000_ vssd1 vssd1 vccd1 vccd1 _0306_ sky130_fd_sc_hd__o211a_1
XFILLER_76_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6177_ egd_top.BitStream_buffer.pc_previous\[1\] egd_top.BitStream_buffer.exp_golomb_len\[1\]
+ vssd1 vssd1 vccd1 vccd1 _2577_ sky130_fd_sc_hd__nand2_1
X_3389_ egd_top.BitStream_buffer.pc\[6\] _2936_ _2942_ vssd1 vssd1 vccd1 vccd1 _2943_
+ sky130_fd_sc_hd__or3b_1
XFILLER_84_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5128_ _3310_ _3338_ vssd1 vssd1 vccd1 vccd1 _1634_ sky130_fd_sc_hd__nand2_1
XFILLER_84_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5059_ _3028_ _1564_ _3341_ _3333_ _1565_ vssd1 vssd1 vccd1 vccd1 _1566_ sky130_fd_sc_hd__a221o_1
XFILLER_52_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4430_ _0370_ _0364_ vssd1 vssd1 vccd1 vccd1 _0941_ sky130_fd_sc_hd__nand2_1
XANTENNA_2 _0295_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4361_ _0389_ _0378_ _0869_ _0382_ _0872_ vssd1 vssd1 vccd1 vccd1 _0873_ sky130_fd_sc_hd__a221oi_1
X_6100_ _2531_ vssd1 vssd1 vccd1 vccd1 _2532_ sky130_fd_sc_hd__buf_2
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4292_ egd_top.BitStream_buffer.BS_buffer\[107\] vssd1 vssd1 vccd1 vccd1 _0804_ sky130_fd_sc_hd__clkinv_2
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6031_ _2982_ _2487_ _2488_ _2492_ vssd1 vssd1 vccd1 vccd1 _0245_ sky130_fd_sc_hd__o211a_1
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5815_ _3288_ _3216_ _3293_ _3220_ _2314_ vssd1 vssd1 vccd1 vccd1 _2315_ sky130_fd_sc_hd__a221oi_1
XFILLER_34_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6795_ net39 _0254_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_5746_ _2237_ _2241_ _2244_ _2246_ vssd1 vssd1 vccd1 vccd1 _2247_ sky130_fd_sc_hd__and4_1
XFILLER_41_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5677_ _2993_ _3123_ _2178_ vssd1 vssd1 vccd1 vccd1 _2179_ sky130_fd_sc_hd__o21ai_1
X_4628_ _0366_ _0545_ _1137_ vssd1 vssd1 vccd1 vccd1 _1138_ sky130_fd_sc_hd__o21ai_1
XFILLER_89_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4559_ _1066_ _1067_ _1068_ _1069_ vssd1 vssd1 vccd1 vccd1 _1070_ sky130_fd_sc_hd__and4_1
X_6229_ _2992_ _2602_ _2570_ _2610_ vssd1 vssd1 vccd1 vccd1 _0171_ sky130_fd_sc_hd__o211a_1
XFILLER_49_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__2887_ clknet_0__2887_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__2887_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_48_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3930_ _0442_ _0443_ vssd1 vssd1 vccd1 vccd1 _0444_ sky130_fd_sc_hd__nand2_1
X_6632__9 clknet_1_1__leaf__2893_ vssd1 vssd1 vccd1 vccd1 net43 sky130_fd_sc_hd__inv_2
X_3861_ egd_top.BitStream_buffer.BS_buffer\[40\] vssd1 vssd1 vccd1 vccd1 _0375_ sky130_fd_sc_hd__clkbuf_4
XFILLER_16_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5600_ _0564_ egd_top.BitStream_buffer.BS_buffer\[16\] vssd1 vssd1 vccd1 vccd1 _2102_
+ sky130_fd_sc_hd__nand2_1
X_3792_ _3325_ vssd1 vssd1 vccd1 vccd1 _3326_ sky130_fd_sc_hd__buf_2
X_6580_ clknet_1_1__leaf__2883_ vssd1 vssd1 vccd1 vccd1 _2889_ sky130_fd_sc_hd__buf_1
XFILLER_31_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5531_ _1043_ _0464_ _2031_ _2032_ _2033_ vssd1 vssd1 vccd1 vccd1 _2034_ sky130_fd_sc_hd__o2111a_1
X_6538__83 clknet_1_1__leaf__2885_ vssd1 vssd1 vccd1 vccd1 net117 sky130_fd_sc_hd__inv_2
X_5462_ _0746_ _3113_ _3117_ _3191_ _1964_ vssd1 vssd1 vccd1 vccd1 _1965_ sky130_fd_sc_hd__a221oi_1
X_6553__97 clknet_1_0__leaf__2886_ vssd1 vssd1 vccd1 vccd1 net131 sky130_fd_sc_hd__inv_2
X_4413_ _0602_ _0613_ vssd1 vssd1 vccd1 vccd1 _0925_ sky130_fd_sc_hd__or2_1
X_5393_ _3085_ _0327_ _1896_ vssd1 vssd1 vccd1 vccd1 _1897_ sky130_fd_sc_hd__o21ai_1
X_4344_ _0854_ _0327_ _0855_ vssd1 vssd1 vccd1 vccd1 _0856_ sky130_fd_sc_hd__o21ai_1
XFILLER_86_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6014_ _3014_ _2466_ _2474_ _2481_ vssd1 vssd1 vccd1 vccd1 _0251_ sky130_fd_sc_hd__o211a_1
X_4275_ _3028_ _0323_ _3341_ _3340_ _0787_ vssd1 vssd1 vccd1 vccd1 _0788_ sky130_fd_sc_hd__a221oi_2
XTAP_186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6847_ net91 _0306_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[119\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_50_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6778_ net182 _0237_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[42\]
+ sky130_fd_sc_hd__dfxtp_1
X_5729_ _0605_ _0527_ vssd1 vssd1 vccd1 vccd1 _2230_ sky130_fd_sc_hd__nand2_1
XFILLER_22_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4060_ egd_top.BitStream_buffer.BS_buffer\[11\] vssd1 vssd1 vccd1 vccd1 _0574_ sky130_fd_sc_hd__inv_2
XFILLER_49_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4962_ _0869_ _0342_ _0345_ _0393_ _1468_ vssd1 vssd1 vccd1 vccd1 _1469_ sky130_fd_sc_hd__a221oi_1
X_3913_ _0420_ _0422_ _0426_ vssd1 vssd1 vccd1 vccd1 _0427_ sky130_fd_sc_hd__o21ai_1
X_4893_ _0771_ _3298_ _1398_ _1399_ _1400_ vssd1 vssd1 vccd1 vccd1 _1401_ sky130_fd_sc_hd__o2111a_1
XFILLER_51_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3844_ _3052_ _0338_ vssd1 vssd1 vccd1 vccd1 _0358_ sky130_fd_sc_hd__and2_1
X_3775_ _3290_ _3097_ vssd1 vssd1 vccd1 vccd1 _3309_ sky130_fd_sc_hd__nor2_2
X_5514_ _0400_ _0360_ _0363_ _0407_ _2016_ vssd1 vssd1 vccd1 vccd1 _2017_ sky130_fd_sc_hd__a221oi_2
X_6494_ _2855_ egd_top.BitStream_buffer.BitStream_buffer_output\[7\] vssd1 vssd1 vccd1
+ vccd1 _2856_ sky130_fd_sc_hd__nand2_1
X_5445_ _3333_ _3062_ vssd1 vssd1 vccd1 vccd1 _1948_ sky130_fd_sc_hd__nand2_1
X_5376_ _0606_ _0515_ vssd1 vssd1 vccd1 vccd1 _1880_ sky130_fd_sc_hd__nand2_1
X_4327_ _0767_ _3279_ _0838_ vssd1 vssd1 vccd1 vccd1 _0839_ sky130_fd_sc_hd__o21ai_1
XFILLER_59_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4258_ egd_top.BitStream_buffer.BS_buffer\[86\] vssd1 vssd1 vccd1 vccd1 _0771_ sky130_fd_sc_hd__clkinv_2
XFILLER_47_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4189_ _0537_ vssd1 vssd1 vccd1 vccd1 _0702_ sky130_fd_sc_hd__inv_2
XFILLER_42_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_0__2889_ _2889_ vssd1 vssd1 vccd1 vccd1 clknet_0__2889_ sky130_fd_sc_hd__clkbuf_16
XFILLER_12_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6532__78 clknet_1_1__leaf__2884_ vssd1 vssd1 vccd1 vccd1 net112 sky130_fd_sc_hd__inv_2
XFILLER_88_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6577__119 clknet_1_0__leaf__2888_ vssd1 vssd1 vccd1 vccd1 net153 sky130_fd_sc_hd__inv_2
XFILLER_33_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3560_ egd_top.BitStream_buffer.BS_buffer\[100\] vssd1 vssd1 vccd1 vccd1 _3094_ sky130_fd_sc_hd__clkbuf_4
X_5230_ _0713_ _0326_ _1734_ vssd1 vssd1 vccd1 vccd1 _1735_ sky130_fd_sc_hd__o21ai_1
X_3491_ _3023_ _2976_ _3002_ _3025_ vssd1 vssd1 vccd1 vccd1 _0298_ sky130_fd_sc_hd__o211a_1
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5161_ _3238_ _0464_ vssd1 vssd1 vccd1 vccd1 _1667_ sky130_fd_sc_hd__or2_1
X_5092_ _3074_ _0746_ vssd1 vssd1 vccd1 vccd1 _1598_ sky130_fd_sc_hd__nand2_1
XFILLER_68_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4112_ egd_top.BitStream_buffer.BitStream_buffer_output\[15\] _2964_ _2901_ vssd1
+ vssd1 vccd1 vccd1 _0626_ sky130_fd_sc_hd__o21a_1
X_4043_ _3087_ _0556_ vssd1 vssd1 vccd1 vccd1 _0557_ sky130_fd_sc_hd__nand2_2
XFILLER_68_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6692__63 clknet_1_0__leaf__2899_ vssd1 vssd1 vccd1 vccd1 net97 sky130_fd_sc_hd__inv_2
XFILLER_83_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5994_ _2985_ _2465_ _2458_ _2470_ vssd1 vssd1 vccd1 vccd1 _0260_ sky130_fd_sc_hd__o211a_1
X_4945_ _3147_ egd_top.BitStream_buffer.BS_buffer\[127\] vssd1 vssd1 vccd1 vccd1 _1453_
+ sky130_fd_sc_hd__nand2_1
XFILLER_33_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4876_ _0503_ _0531_ vssd1 vssd1 vccd1 vccd1 _1384_ sky130_fd_sc_hd__nand2_1
XFILLER_20_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3827_ _0340_ vssd1 vssd1 vccd1 vccd1 _0341_ sky130_fd_sc_hd__clkbuf_2
X_3758_ _3291_ vssd1 vssd1 vccd1 vccd1 _3292_ sky130_fd_sc_hd__buf_4
X_3689_ _3222_ vssd1 vssd1 vccd1 vccd1 _3223_ sky130_fd_sc_hd__clkbuf_2
X_6477_ _1586_ _2839_ vssd1 vssd1 vccd1 vccd1 _2840_ sky130_fd_sc_hd__nor2_1
X_5428_ _3168_ _3133_ vssd1 vssd1 vccd1 vccd1 _1932_ sky130_fd_sc_hd__nand2_1
X_5359_ _0699_ _0495_ _1862_ vssd1 vssd1 vccd1 vccd1 _1863_ sky130_fd_sc_hd__o21ai_1
XFILLER_59_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4730_ _3175_ egd_top.BitStream_buffer.BS_buffer\[1\] vssd1 vssd1 vccd1 vccd1 _1239_
+ sky130_fd_sc_hd__nand2_1
XFILLER_14_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4661_ _1169_ _0327_ _1170_ vssd1 vssd1 vccd1 vccd1 _1171_ sky130_fd_sc_hd__o21ai_1
X_3612_ _3121_ _3134_ vssd1 vssd1 vccd1 vccd1 _3146_ sky130_fd_sc_hd__and2_1
X_6400_ _2767_ _2685_ vssd1 vssd1 vccd1 vccd1 _2769_ sky130_fd_sc_hd__nand2_1
X_4592_ _0441_ _0454_ vssd1 vssd1 vccd1 vccd1 _1102_ sky130_fd_sc_hd__nand2_1
X_6331_ egd_top.BitStream_buffer.BitStream_buffer_output\[8\] egd_top.BitStream_buffer.BitStream_buffer_output\[7\]
+ vssd1 vssd1 vccd1 vccd1 _2702_ sky130_fd_sc_hd__nor2_1
X_3543_ _3076_ vssd1 vssd1 vccd1 vccd1 _3077_ sky130_fd_sc_hd__inv_2
X_6262_ egd_top.BitStream_buffer.BitStream_buffer_output\[10\] _2632_ vssd1 vssd1
+ vccd1 vccd1 _2633_ sky130_fd_sc_hd__or2_1
X_3474_ _2989_ _3012_ vssd1 vssd1 vccd1 vccd1 _3013_ sky130_fd_sc_hd__nand2_1
XFILLER_88_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5213_ _3092_ _3070_ vssd1 vssd1 vccd1 vccd1 _1718_ sky130_fd_sc_hd__nand2_1
X_6193_ _2902_ egd_top.BitStream_buffer.pc\[5\] vssd1 vssd1 vccd1 vccd1 _2590_ sky130_fd_sc_hd__nand2_1
X_5144_ _0879_ _0385_ _1649_ vssd1 vssd1 vccd1 vccd1 _1650_ sky130_fd_sc_hd__o21ai_1
XFILLER_84_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5075_ _1567_ _1581_ vssd1 vssd1 vccd1 vccd1 _1582_ sky130_fd_sc_hd__nand2_1
XFILLER_84_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4026_ egd_top.BitStream_buffer.BS_buffer\[31\] vssd1 vssd1 vccd1 vccd1 _0540_ sky130_fd_sc_hd__clkbuf_4
XFILLER_71_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5977_ _2449_ _0611_ vssd1 vssd1 vccd1 vccd1 _2460_ sky130_fd_sc_hd__nand2_1
X_4928_ _3254_ _3302_ vssd1 vssd1 vccd1 vccd1 _1436_ sky130_fd_sc_hd__nand2_1
XFILLER_40_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4859_ _0574_ _0570_ vssd1 vssd1 vccd1 vccd1 _1367_ sky130_fd_sc_hd__or2_1
XFILLER_20_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6671__44 clknet_1_1__leaf__2897_ vssd1 vssd1 vccd1 vccd1 net78 sky130_fd_sc_hd__inv_2
XFILLER_47_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_80 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5900_ _2385_ _2399_ vssd1 vssd1 vccd1 vccd1 _2400_ sky130_fd_sc_hd__nand2_1
XFILLER_81_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5831_ _3126_ _3191_ vssd1 vssd1 vccd1 vccd1 _2331_ sky130_fd_sc_hd__nand2_1
XFILLER_61_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5762_ _3148_ _0562_ vssd1 vssd1 vccd1 vccd1 _2263_ sky130_fd_sc_hd__nand2_1
XFILLER_61_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4713_ _1210_ _1214_ _1218_ _1221_ vssd1 vssd1 vccd1 vccd1 _1222_ sky130_fd_sc_hd__and4_1
X_5693_ _0370_ _0400_ vssd1 vssd1 vccd1 vccd1 _2194_ sky130_fd_sc_hd__nand2_1
X_4644_ _3271_ _0837_ vssd1 vssd1 vccd1 vccd1 _1154_ sky130_fd_sc_hd__nand2_1
X_4575_ _0370_ _0337_ vssd1 vssd1 vccd1 vccd1 _1085_ sky130_fd_sc_hd__nand2_1
XFILLER_89_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3526_ _3041_ _3059_ vssd1 vssd1 vccd1 vccd1 _3060_ sky130_fd_sc_hd__nor2_2
X_6314_ _2683_ _2684_ vssd1 vssd1 vccd1 vccd1 _2685_ sky130_fd_sc_hd__nand2_2
X_6245_ _2608_ _0324_ vssd1 vssd1 vccd1 vccd1 _2619_ sky130_fd_sc_hd__nand2_1
X_3457_ _2989_ _2999_ vssd1 vssd1 vccd1 vccd1 _3000_ sky130_fd_sc_hd__nand2_1
XFILLER_39_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6176_ egd_top.BitStream_buffer.pc_previous\[1\] egd_top.BitStream_buffer.exp_golomb_len\[1\]
+ vssd1 vssd1 vccd1 vccd1 _2576_ sky130_fd_sc_hd__or2_1
X_3388_ _2941_ egd_top.BitStream_buffer.pc_previous\[4\] egd_top.BitStream_buffer.pc_previous\[5\]
+ egd_top.BitStream_buffer.pc_previous\[6\] vssd1 vssd1 vccd1 vccd1 _2942_ sky130_fd_sc_hd__a31o_1
XFILLER_69_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_424 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5127_ _3314_ _0330_ vssd1 vssd1 vccd1 vccd1 _1633_ sky130_fd_sc_hd__nand2_1
XFILLER_55_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5058_ _3040_ _3323_ _3325_ _0708_ vssd1 vssd1 vccd1 vccd1 _1565_ sky130_fd_sc_hd__a22o_1
X_4009_ _0522_ vssd1 vssd1 vccd1 vccd1 _0523_ sky130_fd_sc_hd__buf_2
XFILLER_55_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6614__152 clknet_1_1__leaf__2892_ vssd1 vssd1 vccd1 vccd1 net186 sky130_fd_sc_hd__inv_2
XFILLER_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_3 _0569_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4360_ _0870_ _0385_ _0871_ vssd1 vssd1 vccd1 vccd1 _0872_ sky130_fd_sc_hd__o21ai_1
XFILLER_6_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4291_ _3119_ _3089_ _0800_ _0801_ _0802_ vssd1 vssd1 vccd1 vccd1 _0803_ sky130_fd_sc_hd__o2111a_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6030_ _2489_ _0633_ vssd1 vssd1 vccd1 vccd1 _2492_ sky130_fd_sc_hd__nand2_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6650__25 clknet_1_0__leaf__2895_ vssd1 vssd1 vccd1 vccd1 net59 sky130_fd_sc_hd__inv_2
XFILLER_54_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5814_ _3317_ _1145_ _2313_ vssd1 vssd1 vccd1 vccd1 _2314_ sky130_fd_sc_hd__o21ai_1
XFILLER_34_173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6794_ net38 _0253_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_5745_ _1084_ _0522_ _0629_ _0525_ _2245_ vssd1 vssd1 vccd1 vccd1 _2246_ sky130_fd_sc_hd__o221a_1
X_5676_ _3127_ _3204_ vssd1 vssd1 vccd1 vccd1 _2178_ sky130_fd_sc_hd__nand2_1
XFILLER_30_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4627_ _0547_ egd_top.BitStream_buffer.BS_buffer\[32\] vssd1 vssd1 vccd1 vccd1 _1137_
+ sky130_fd_sc_hd__nand2_1
X_4558_ _3136_ egd_top.BitStream_buffer.BS_buffer\[125\] vssd1 vssd1 vccd1 vccd1 _1069_
+ sky130_fd_sc_hd__nand2_1
X_4489_ _0524_ _0522_ _0702_ _0525_ _0999_ vssd1 vssd1 vccd1 vccd1 _1000_ sky130_fd_sc_hd__o221a_1
X_3509_ _3042_ vssd1 vssd1 vccd1 vccd1 _3043_ sky130_fd_sc_hd__inv_2
X_6228_ _2608_ _3317_ vssd1 vssd1 vccd1 vccd1 _2610_ sky130_fd_sc_hd__nand2_1
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6159_ _3001_ _2554_ _2558_ _2566_ vssd1 vssd1 vccd1 vccd1 _0191_ sky130_fd_sc_hd__o211a_1
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_427 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_110 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1__f__2886_ clknet_0__2886_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__2886_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_63_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3860_ egd_top.BitStream_buffer.BS_buffer\[34\] _0360_ _0363_ _0364_ _0373_ vssd1
+ vssd1 vccd1 vccd1 _0374_ sky130_fd_sc_hd__a221oi_1
XFILLER_72_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3791_ _3290_ _3115_ vssd1 vssd1 vccd1 vccd1 _3325_ sky130_fd_sc_hd__nor2_2
XFILLER_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5530_ _0755_ _0449_ vssd1 vssd1 vccd1 vccd1 _2033_ sky130_fd_sc_hd__or2_1
X_5461_ _2990_ _3122_ _1963_ vssd1 vssd1 vccd1 vccd1 _1964_ sky130_fd_sc_hd__o21ai_1
X_4412_ _0609_ egd_top.BitStream_buffer.BS_buffer\[16\] vssd1 vssd1 vccd1 vccd1 _0924_
+ sky130_fd_sc_hd__nand2_1
XFILLER_8_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5392_ _0329_ _3100_ vssd1 vssd1 vccd1 vccd1 _1896_ sky130_fd_sc_hd__nand2_1
X_4343_ _0329_ _3338_ vssd1 vssd1 vccd1 vccd1 _0855_ sky130_fd_sc_hd__nand2_1
X_4274_ _0784_ _0327_ _0786_ vssd1 vssd1 vccd1 vccd1 _0787_ sky130_fd_sc_hd__o21ai_1
X_6013_ _2471_ _0699_ vssd1 vssd1 vccd1 vccd1 _2481_ sky130_fd_sc_hd__nand2_1
XTAP_187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6846_ net90 _0305_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[120\]
+ sky130_fd_sc_hd__dfxtp_2
X_6777_ net181 _0236_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[43\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_50_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3989_ _0488_ _3091_ vssd1 vssd1 vccd1 vccd1 _0503_ sky130_fd_sc_hd__nor2_2
X_5728_ _0608_ egd_top.BitStream_buffer.BS_buffer\[27\] vssd1 vssd1 vccd1 vccd1 _2229_
+ sky130_fd_sc_hd__nand2_1
XFILLER_50_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5659_ _3168_ _3173_ vssd1 vssd1 vccd1 vccd1 _2161_ sky130_fd_sc_hd__nand2_1
XFILLER_89_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4961_ _1466_ _0350_ _1467_ vssd1 vssd1 vccd1 vccd1 _1468_ sky130_fd_sc_hd__o21ai_1
XFILLER_17_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3912_ _0423_ _0425_ vssd1 vssd1 vccd1 vccd1 _0426_ sky130_fd_sc_hd__or2_1
X_4892_ _3294_ _0780_ vssd1 vssd1 vccd1 vccd1 _1400_ sky130_fd_sc_hd__nand2_1
X_3843_ _0337_ _0342_ _0345_ _0346_ _0356_ vssd1 vssd1 vccd1 vccd1 _0357_ sky130_fd_sc_hd__a221oi_1
XFILLER_32_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3774_ _3307_ vssd1 vssd1 vccd1 vccd1 _3308_ sky130_fd_sc_hd__clkbuf_4
X_5513_ _0637_ _0368_ _2015_ vssd1 vssd1 vccd1 vccd1 _2016_ sky130_fd_sc_hd__o21ai_1
X_6493_ _2723_ vssd1 vssd1 vccd1 vccd1 _2855_ sky130_fd_sc_hd__inv_2
XFILLER_8_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5444_ egd_top.BitStream_buffer.BitStream_buffer_output\[4\] _2965_ _0627_ vssd1
+ vssd1 vccd1 vccd1 _1947_ sky130_fd_sc_hd__o21ai_1
X_5375_ _0609_ _0519_ vssd1 vssd1 vccd1 vccd1 _1879_ sky130_fd_sc_hd__nand2_1
X_4326_ _3282_ _0837_ vssd1 vssd1 vccd1 vccd1 _0838_ sky130_fd_sc_hd__nand2_1
XFILLER_59_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4257_ _3293_ _3292_ _3315_ _3295_ _0769_ vssd1 vssd1 vccd1 vccd1 _0770_ sky130_fd_sc_hd__a221oi_1
X_4188_ _0528_ _0523_ _0699_ _0526_ _0700_ vssd1 vssd1 vccd1 vccd1 _0701_ sky130_fd_sc_hd__o221a_1
XFILLER_67_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6829_ net73 _0288_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BitStream_buffer_output\[6\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_23_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_0__2888_ _2888_ vssd1 vssd1 vccd1 vccd1 clknet_0__2888_ sky130_fd_sc_hd__clkbuf_16
XFILLER_23_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3490_ _2974_ _3024_ vssd1 vssd1 vccd1 vccd1 _3025_ sky130_fd_sc_hd__nand2_1
X_6677__50 clknet_1_1__leaf__2897_ vssd1 vssd1 vccd1 vccd1 net84 sky130_fd_sc_hd__inv_2
X_5160_ _0453_ _3244_ vssd1 vssd1 vccd1 vccd1 _1666_ sky130_fd_sc_hd__nand2_1
XFILLER_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5091_ _3153_ _3113_ _3117_ _3157_ _1596_ vssd1 vssd1 vccd1 vccd1 _1597_ sky130_fd_sc_hd__a221oi_1
X_4111_ _0336_ _0618_ _0624_ vssd1 vssd1 vccd1 vccd1 _0625_ sky130_fd_sc_hd__nand3_1
XFILLER_68_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4042_ _0555_ vssd1 vssd1 vccd1 vccd1 _0556_ sky130_fd_sc_hd__clkbuf_4
XFILLER_37_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5993_ _2466_ _0692_ vssd1 vssd1 vccd1 vccd1 _2470_ sky130_fd_sc_hd__nand2_1
XFILLER_91_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4944_ _1448_ _1449_ _1450_ _1451_ vssd1 vssd1 vccd1 vccd1 _1452_ sky130_fd_sc_hd__and4_1
XFILLER_64_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4875_ _0520_ _0494_ _1380_ _1381_ _1382_ vssd1 vssd1 vccd1 vccd1 _1383_ sky130_fd_sc_hd__o2111a_1
X_3826_ _3090_ _0339_ vssd1 vssd1 vccd1 vccd1 _0340_ sky130_fd_sc_hd__and2_1
X_3757_ _3290_ _3053_ vssd1 vssd1 vccd1 vccd1 _3291_ sky130_fd_sc_hd__nor2_2
XFILLER_20_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3688_ _3096_ _3213_ vssd1 vssd1 vccd1 vccd1 _3222_ sky130_fd_sc_hd__and2_1
X_6476_ egd_top.BitStream_buffer.BitStream_buffer_output\[6\] _2723_ vssd1 vssd1 vccd1
+ vccd1 _2839_ sky130_fd_sc_hd__nor2_1
X_5427_ _3163_ _3138_ vssd1 vssd1 vccd1 vccd1 _1931_ sky130_fd_sc_hd__nand2_1
X_5358_ _0497_ egd_top.BitStream_buffer.BS_buffer\[29\] vssd1 vssd1 vccd1 vccd1 _1862_
+ sky130_fd_sc_hd__nand2_1
XFILLER_58_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4309_ _3187_ _3180_ _0792_ _3186_ _0820_ vssd1 vssd1 vccd1 vccd1 _0821_ sky130_fd_sc_hd__a221oi_2
XFILLER_59_135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5289_ _0965_ _0403_ _1793_ vssd1 vssd1 vccd1 vccd1 _1794_ sky130_fd_sc_hd__o21ai_1
XFILLER_28_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6583__124 clknet_1_0__leaf__2889_ vssd1 vssd1 vccd1 vccd1 net158 sky130_fd_sc_hd__inv_2
XFILLER_48_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4660_ _0329_ egd_top.BitStream_buffer.BS_buffer\[96\] vssd1 vssd1 vccd1 vccd1 _1170_
+ sky130_fd_sc_hd__nand2_1
X_3611_ _3144_ vssd1 vssd1 vccd1 vccd1 _3145_ sky130_fd_sc_hd__inv_2
X_6330_ _2676_ _2682_ _2926_ vssd1 vssd1 vccd1 vccd1 _2701_ sky130_fd_sc_hd__a21oi_4
X_4591_ _0431_ egd_top.BitStream_buffer.BS_buffer\[58\] vssd1 vssd1 vccd1 vccd1 _1101_
+ sky130_fd_sc_hd__nand2_1
X_3542_ _2920_ _3050_ vssd1 vssd1 vccd1 vccd1 _3076_ sky130_fd_sc_hd__nor2_2
X_6261_ _2622_ _2631_ vssd1 vssd1 vccd1 vccd1 _2632_ sky130_fd_sc_hd__nand2_1
X_3473_ egd_top.BitStream_buffer.BS_buffer\[123\] vssd1 vssd1 vccd1 vccd1 _3012_ sky130_fd_sc_hd__inv_2
X_5212_ _3098_ _3082_ vssd1 vssd1 vccd1 vccd1 _1717_ sky130_fd_sc_hd__nand2_1
X_6192_ _2587_ _2589_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.pc\[5\] sky130_fd_sc_hd__nor2_4
XFILLER_69_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5143_ _0388_ _0412_ vssd1 vssd1 vccd1 vccd1 _1649_ sky130_fd_sc_hd__nand2_1
XFILLER_69_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5074_ _1570_ _1573_ _1577_ _1580_ vssd1 vssd1 vccd1 vccd1 _1581_ sky130_fd_sc_hd__and4_1
X_4025_ _0538_ vssd1 vssd1 vccd1 vccd1 _0539_ sky130_fd_sc_hd__buf_2
XFILLER_56_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5976_ _3014_ _2443_ _2458_ _2459_ vssd1 vssd1 vccd1 vccd1 _0267_ sky130_fd_sc_hd__o211a_1
XFILLER_12_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4927_ _3262_ egd_top.BitStream_buffer.BS_buffer\[79\] vssd1 vssd1 vccd1 vccd1 _1435_
+ sky130_fd_sc_hd__nand2_1
X_4858_ _0560_ egd_top.BitStream_buffer.BS_buffer\[12\] vssd1 vssd1 vccd1 vccd1 _1366_
+ sky130_fd_sc_hd__nand2_1
X_3809_ _0322_ vssd1 vssd1 vccd1 vccd1 _0323_ sky130_fd_sc_hd__clkbuf_4
X_4789_ _0469_ _0751_ vssd1 vssd1 vccd1 vccd1 _1298_ sky130_fd_sc_hd__nand2_1
X_6459_ _2816_ _2684_ vssd1 vssd1 vccd1 vccd1 _2823_ sky130_fd_sc_hd__nand2_1
X_6656__31 clknet_1_1__leaf__2895_ vssd1 vssd1 vccd1 vccd1 net65 sky130_fd_sc_hd__inv_2
XFILLER_75_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5830_ _2993_ _3089_ _2327_ _2328_ _2329_ vssd1 vssd1 vccd1 vccd1 _2330_ sky130_fd_sc_hd__o2111a_1
X_5761_ _2251_ _2255_ _2258_ _2261_ vssd1 vssd1 vccd1 vccd1 _2262_ sky130_fd_sc_hd__and4_1
X_4712_ _3062_ _3340_ _3094_ _0323_ _1220_ vssd1 vssd1 vccd1 vccd1 _1221_ sky130_fd_sc_hd__a221oi_1
X_5692_ _0948_ _0341_ _0344_ _0412_ _2192_ vssd1 vssd1 vccd1 vccd1 _2193_ sky130_fd_sc_hd__a221oi_1
X_4643_ _3278_ vssd1 vssd1 vccd1 vccd1 _1153_ sky130_fd_sc_hd__inv_2
X_4574_ _0346_ vssd1 vssd1 vccd1 vccd1 _1084_ sky130_fd_sc_hd__inv_2
X_3525_ _3058_ vssd1 vssd1 vccd1 vccd1 _3059_ sky130_fd_sc_hd__clkinv_2
X_6313_ _2924_ vssd1 vssd1 vccd1 vccd1 _2684_ sky130_fd_sc_hd__clkbuf_4
XFILLER_89_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6244_ _3014_ _2603_ _2611_ _2618_ vssd1 vssd1 vccd1 vccd1 _0164_ sky130_fd_sc_hd__o211a_1
X_3456_ egd_top.BitStream_buffer.BS_buffer\[119\] vssd1 vssd1 vccd1 vccd1 _2999_ sky130_fd_sc_hd__clkinv_2
X_3387_ egd_top.BitStream_buffer.pc_previous\[0\] egd_top.BitStream_buffer.pc_previous\[1\]
+ egd_top.BitStream_buffer.pc_previous\[2\] egd_top.BitStream_buffer.pc_previous\[3\]
+ vssd1 vssd1 vccd1 vccd1 _2941_ sky130_fd_sc_hd__and4_1
X_6175_ egd_top.BitStream_buffer.pc_previous\[5\] vssd1 vssd1 vccd1 vccd1 _2575_ sky130_fd_sc_hd__inv_2
X_5126_ _3322_ _3292_ _3327_ _3295_ _1631_ vssd1 vssd1 vccd1 vccd1 _1632_ sky130_fd_sc_hd__a221oi_1
XFILLER_57_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5057_ _3329_ vssd1 vssd1 vccd1 vccd1 _1564_ sky130_fd_sc_hd__inv_2
XFILLER_84_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4008_ _0521_ _3030_ vssd1 vssd1 vccd1 vccd1 _0522_ sky130_fd_sc_hd__nand2_2
XFILLER_52_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5959_ _2988_ _2442_ _2446_ _2450_ vssd1 vssd1 vccd1 vccd1 _0275_ sky130_fd_sc_hd__o211a_1
XFILLER_0_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6701__1 clknet_1_0__leaf__2883_ vssd1 vssd1 vccd1 vccd1 net35 sky130_fd_sc_hd__inv_2
XANTENNA_4 _0691_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6589__130 clknet_1_1__leaf__2889_ vssd1 vssd1 vccd1 vccd1 net164 sky130_fd_sc_hd__inv_2
X_4290_ _3085_ _3106_ vssd1 vssd1 vccd1 vccd1 _0802_ sky130_fd_sc_hd__or2_1
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6862_ net35 _0321_ vssd1 vssd1 vccd1 vccd1 net34 sky130_fd_sc_hd__dfxtp_2
XFILLER_34_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5813_ _3223_ _3315_ vssd1 vssd1 vccd1 vccd1 _2313_ sky130_fd_sc_hd__nand2_1
XFILLER_34_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6793_ net37 _0252_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[27\]
+ sky130_fd_sc_hd__dfxtp_4
X_5744_ _1276_ _0529_ _0348_ _0533_ vssd1 vssd1 vccd1 vccd1 _2245_ sky130_fd_sc_hd__o22a_1
X_5675_ _2980_ _3106_ _2174_ _2175_ _2176_ vssd1 vssd1 vccd1 vccd1 _2177_ sky130_fd_sc_hd__o2111a_1
X_4626_ _0699_ _0522_ _0702_ _0534_ _1135_ vssd1 vssd1 vccd1 vccd1 _1136_ sky130_fd_sc_hd__o221a_1
X_4557_ _3144_ egd_top.BitStream_buffer.BS_buffer\[123\] vssd1 vssd1 vccd1 vccd1 _1068_
+ sky130_fd_sc_hd__nand2_1
XFILLER_89_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4488_ _0699_ _0529_ _0543_ _0533_ vssd1 vssd1 vccd1 vccd1 _0999_ sky130_fd_sc_hd__o22a_1
X_3508_ egd_top.BitStream_buffer.pc\[1\] _2929_ vssd1 vssd1 vccd1 vccd1 _3042_ sky130_fd_sc_hd__or2_1
XFILLER_89_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6227_ _2988_ _2602_ _2570_ _2609_ vssd1 vssd1 vccd1 vccd1 _0172_ sky130_fd_sc_hd__o211a_1
X_3439_ egd_top.BitStream_buffer.BS_buffer\[115\] vssd1 vssd1 vccd1 vccd1 _2986_ sky130_fd_sc_hd__clkinv_2
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6158_ _2561_ _0718_ vssd1 vssd1 vccd1 vccd1 _2566_ sky130_fd_sc_hd__nand2_1
X_5109_ _0566_ _3176_ _0568_ _3180_ _1614_ vssd1 vssd1 vccd1 vccd1 _1615_ sky130_fd_sc_hd__a221oi_1
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6089_ _3011_ _2511_ _2516_ _2525_ vssd1 vssd1 vccd1 vccd1 _0220_ sky130_fd_sc_hd__o211a_1
XFILLER_45_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput30 net30 vssd1 vssd1 vccd1 vccd1 la_data_out_26_24[2] sky130_fd_sc_hd__buf_12
XFILLER_68_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__2885_ clknet_0__2885_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__2885_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_88_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3790_ _3323_ vssd1 vssd1 vccd1 vccd1 _3324_ sky130_fd_sc_hd__buf_2
XFILLER_31_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5460_ _3126_ _3157_ vssd1 vssd1 vccd1 vccd1 _1963_ sky130_fd_sc_hd__nand2_1
X_4411_ _0606_ egd_top.BitStream_buffer.BS_buffer\[14\] vssd1 vssd1 vccd1 vccd1 _0923_
+ sky130_fd_sc_hd__nand2_1
XFILLER_68_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5391_ _1169_ _3308_ _1892_ _1893_ _1894_ vssd1 vssd1 vccd1 vccd1 _1895_ sky130_fd_sc_hd__o2111a_1
X_4342_ egd_top.BitStream_buffer.BS_buffer\[95\] vssd1 vssd1 vccd1 vccd1 _0854_ sky130_fd_sc_hd__clkinv_2
X_4273_ _0329_ _0785_ vssd1 vssd1 vccd1 vccd1 _0786_ sky130_fd_sc_hd__nand2_1
XFILLER_86_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6012_ _3011_ _2466_ _2474_ _2480_ vssd1 vssd1 vccd1 vccd1 _0252_ sky130_fd_sc_hd__o211a_1
.ends

